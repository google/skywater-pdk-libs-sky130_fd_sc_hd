* File: sky130_fd_sc_hd__mux2_2.pxi.spice
* Created: Thu Aug 27 14:27:35 2020
* 
x_PM_SKY130_FD_SC_HD__MUX2_2%A_79_21# N_A_79_21#_M1008_d N_A_79_21#_M1005_d
+ N_A_79_21#_c_74_n N_A_79_21#_M1007_g N_A_79_21#_M1006_g N_A_79_21#_c_75_n
+ N_A_79_21#_M1011_g N_A_79_21#_M1009_g N_A_79_21#_c_82_n N_A_79_21#_c_76_n
+ N_A_79_21#_c_170_p N_A_79_21#_c_83_n N_A_79_21#_c_128_p N_A_79_21#_c_88_p
+ N_A_79_21#_c_94_p N_A_79_21#_c_89_p N_A_79_21#_c_113_p N_A_79_21#_c_95_p
+ N_A_79_21#_c_104_p N_A_79_21#_c_77_n N_A_79_21#_c_78_n N_A_79_21#_c_79_n
+ PM_SKY130_FD_SC_HD__MUX2_2%A_79_21#
x_PM_SKY130_FD_SC_HD__MUX2_2%A_257_199# N_A_257_199#_M1013_d
+ N_A_257_199#_M1000_d N_A_257_199#_M1004_g N_A_257_199#_M1012_g
+ N_A_257_199#_c_196_n N_A_257_199#_c_197_n N_A_257_199#_c_202_n
+ N_A_257_199#_c_203_n N_A_257_199#_c_204_n N_A_257_199#_c_205_n
+ N_A_257_199#_c_232_n N_A_257_199#_c_198_n N_A_257_199#_c_207_n
+ PM_SKY130_FD_SC_HD__MUX2_2%A_257_199#
x_PM_SKY130_FD_SC_HD__MUX2_2%A0 N_A0_M1008_g N_A0_M1001_g A0 A0 A0 A0
+ N_A0_c_287_n N_A0_c_288_n N_A0_c_289_n PM_SKY130_FD_SC_HD__MUX2_2%A0
x_PM_SKY130_FD_SC_HD__MUX2_2%A1 N_A1_M1005_g N_A1_c_338_n N_A1_c_339_n
+ N_A1_M1002_g A1 A1 N_A1_c_343_n PM_SKY130_FD_SC_HD__MUX2_2%A1
x_PM_SKY130_FD_SC_HD__MUX2_2%S N_S_M1010_g N_S_M1003_g N_S_M1013_g N_S_M1000_g S
+ S S N_S_c_393_n PM_SKY130_FD_SC_HD__MUX2_2%S
x_PM_SKY130_FD_SC_HD__MUX2_2%VPWR N_VPWR_M1006_d N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n VPWR
+ N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_435_n N_VPWR_c_444_n
+ N_VPWR_c_445_n PM_SKY130_FD_SC_HD__MUX2_2%VPWR
x_PM_SKY130_FD_SC_HD__MUX2_2%X N_X_M1007_s N_X_M1006_s N_X_c_498_n N_X_c_499_n
+ N_X_c_501_n N_X_c_496_n X X PM_SKY130_FD_SC_HD__MUX2_2%X
x_PM_SKY130_FD_SC_HD__MUX2_2%VGND N_VGND_M1007_d N_VGND_M1011_d N_VGND_M1010_d
+ N_VGND_c_532_n N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n VGND
+ N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n N_VGND_c_540_n
+ N_VGND_c_541_n PM_SKY130_FD_SC_HD__MUX2_2%VGND
cc_1 VNB N_A_79_21#_c_74_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_75_n 0.0164012f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_76_n 0.00688196f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.72
cc_4 VNB N_A_79_21#_c_77_n 0.00229788f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_5 VNB N_A_79_21#_c_78_n 0.0480844f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_6 VNB N_A_79_21#_c_79_n 0.00180654f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB N_A_257_199#_M1004_g 0.0288566f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB N_A_257_199#_c_196_n 6.23272e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_9 VNB N_A_257_199#_c_197_n 0.0253246f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_10 VNB N_A_257_199#_c_198_n 0.0433249f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=0.635
cc_11 VNB A0 0.0225985f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_12 VNB N_A0_c_287_n 0.0325495f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_13 VNB N_A0_c_288_n 0.0226851f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_14 VNB N_A0_c_289_n 0.00690845f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.72
cc_15 VNB N_A1_M1005_g 0.0152081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A1_c_338_n 0.0155208f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A1_c_339_n 0.00819149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_M1002_g 0.0236688f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB A1 0.00195435f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB A1 0.00780429f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_21 VNB N_A1_c_343_n 0.0258665f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_22 VNB N_S_M1010_g 0.0275685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_S_M1013_g 0.0340185f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_24 VNB S 0.00504577f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_25 VNB N_S_c_393_n 0.0432042f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.92
cc_26 VNB N_VPWR_c_435_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_27 VNB N_X_c_496_n 7.9516e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_28 VNB N_VGND_c_532_n 0.00997339f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_29 VNB N_VGND_c_533_n 0.0330373f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_30 VNB N_VGND_c_534_n 0.00268492f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_31 VNB N_VGND_c_535_n 0.0048408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_536_n 0.0152056f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.835
cc_33 VNB N_VGND_c_537_n 0.0523715f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=0.465
cc_34 VNB N_VGND_c_538_n 0.0177117f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=2.34
cc_35 VNB N_VGND_c_539_n 0.218849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_540_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_37 VNB N_VGND_c_541_n 0.00381743f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_38 VPB N_A_79_21#_M1006_g 0.0253019f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_39 VPB N_A_79_21#_M1009_g 0.0201564f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_40 VPB N_A_79_21#_c_82_n 0.00209021f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.835
cc_41 VPB N_A_79_21#_c_83_n 0.00455708f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.92
cc_42 VPB N_A_79_21#_c_77_n 0.00123788f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_43 VPB N_A_79_21#_c_78_n 0.00829412f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_44 VPB N_A_257_199#_M1012_g 0.0462187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_257_199#_c_196_n 0.00113049f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_46 VPB N_A_257_199#_c_197_n 0.00508966f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_47 VPB N_A_257_199#_c_202_n 0.0164186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_257_199#_c_203_n 0.00157448f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=0.805
cc_49 VPB N_A_257_199#_c_204_n 0.00453643f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.325
cc_50 VPB N_A_257_199#_c_205_n 0.0157254f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.835
cc_51 VPB N_A_257_199#_c_198_n 0.0223369f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=0.635
cc_52 VPB N_A_257_199#_c_207_n 0.0254451f $X=-0.19 $Y=1.305 $X2=1.605 $Y2=0.38
cc_53 VPB N_A0_M1001_g 0.0261971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB A0 6.02903e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_55 VPB A0 0.0105489f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_56 VPB N_A0_c_289_n 0.019355f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=0.72
cc_57 VPB N_A1_M1005_g 0.0471733f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_S_M1003_g 0.0355658f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_59 VPB N_S_M1000_g 0.0450009f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_60 VPB S 0.00644757f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_61 VPB N_S_c_393_n 0.00469193f $X=-0.19 $Y=1.305 $X2=1.165 $Y2=1.92
cc_62 VPB N_VPWR_c_436_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_63 VPB N_VPWR_c_437_n 0.0431346f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_64 VPB N_VPWR_c_438_n 0.00537922f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_65 VPB N_VPWR_c_439_n 0.00495318f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=0.995
cc_66 VPB N_VPWR_c_440_n 0.0183487f $X=-0.19 $Y=1.305 $X2=1.165 $Y2=0.72
cc_67 VPB N_VPWR_c_441_n 0.0498767f $X=-0.19 $Y=1.305 $X2=1.57 $Y2=2.005
cc_68 VPB N_VPWR_c_442_n 0.0171691f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.16
cc_69 VPB N_VPWR_c_435_n 0.0439198f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_70 VPB N_VPWR_c_444_n 0.00554993f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_71 VPB N_VPWR_c_445_n 0.00420071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_496_n 0.0011566f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_73 N_A_79_21#_c_75_n N_A_257_199#_M1004_g 0.0181578f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_74 N_A_79_21#_c_76_n N_A_257_199#_M1004_g 0.0124727f $X=1.435 $Y=0.72 $X2=0
+ $Y2=0
cc_75 N_A_79_21#_c_88_p N_A_257_199#_M1004_g 0.00459008f $X=1.52 $Y=0.635 $X2=0
+ $Y2=0
cc_76 N_A_79_21#_c_89_p N_A_257_199#_M1004_g 0.00380967f $X=1.605 $Y=0.38 $X2=0
+ $Y2=0
cc_77 N_A_79_21#_c_79_n N_A_257_199#_M1004_g 0.002206f $X=1.01 $Y=0.995 $X2=0
+ $Y2=0
cc_78 N_A_79_21#_M1009_g N_A_257_199#_M1012_g 0.0260928f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_79 N_A_79_21#_c_82_n N_A_257_199#_M1012_g 0.00290526f $X=1.08 $Y=1.835 $X2=0
+ $Y2=0
cc_80 N_A_79_21#_c_83_n N_A_257_199#_M1012_g 0.0117505f $X=1.485 $Y=1.92 $X2=0
+ $Y2=0
cc_81 N_A_79_21#_c_94_p N_A_257_199#_M1012_g 0.00794397f $X=1.57 $Y=2.255 $X2=0
+ $Y2=0
cc_82 N_A_79_21#_c_95_p N_A_257_199#_M1012_g 0.00601411f $X=1.655 $Y=2.34 $X2=0
+ $Y2=0
cc_83 N_A_79_21#_c_76_n N_A_257_199#_c_196_n 0.0123545f $X=1.435 $Y=0.72 $X2=0
+ $Y2=0
cc_84 N_A_79_21#_c_77_n N_A_257_199#_c_196_n 0.0374964f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_85 N_A_79_21#_c_78_n N_A_257_199#_c_196_n 3.17464e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_86 N_A_79_21#_c_76_n N_A_257_199#_c_197_n 0.00288902f $X=1.435 $Y=0.72 $X2=0
+ $Y2=0
cc_87 N_A_79_21#_c_83_n N_A_257_199#_c_197_n 0.00160571f $X=1.485 $Y=1.92 $X2=0
+ $Y2=0
cc_88 N_A_79_21#_c_77_n N_A_257_199#_c_197_n 0.00199269f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_79_21#_c_78_n N_A_257_199#_c_197_n 0.0202785f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_90 N_A_79_21#_c_83_n N_A_257_199#_c_202_n 0.0122822f $X=1.485 $Y=1.92 $X2=0
+ $Y2=0
cc_91 N_A_79_21#_c_104_p N_A_257_199#_c_202_n 0.00510386f $X=2.63 $Y=2.34 $X2=0
+ $Y2=0
cc_92 N_A_79_21#_c_82_n N_A_257_199#_c_203_n 0.0140957f $X=1.08 $Y=1.835 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_83_n N_A_257_199#_c_203_n 0.0133813f $X=1.485 $Y=1.92 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_82_n N_A_257_199#_c_204_n 0.00462643f $X=1.08 $Y=1.835 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_M1005_d N_A_257_199#_c_205_n 0.00406618f $X=2.395 $Y=1.845
+ $X2=0 $Y2=0
cc_96 N_A_79_21#_c_104_p N_A_257_199#_c_205_n 0.0311958f $X=2.63 $Y=2.34 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_83_n N_A_257_199#_c_232_n 0.0153287f $X=1.485 $Y=1.92 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_104_p N_A_257_199#_c_232_n 0.00920022f $X=2.63 $Y=2.34 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_76_n A0 0.00299654f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_113_p A0 0.0278634f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_79_n A0 0.00519686f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_113_p N_A0_c_287_n 5.87272e-19 $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_76_n N_A0_c_288_n 0.00388645f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_88_p N_A0_c_288_n 0.00360534f $X=1.52 $Y=0.635 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_113_p N_A0_c_288_n 0.0100917f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_83_n N_A1_M1005_g 3.43672e-19 $X=1.485 $Y=1.92 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_94_p N_A1_M1005_g 0.00367717f $X=1.57 $Y=2.255 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_104_p N_A1_M1005_g 0.0123885f $X=2.63 $Y=2.34 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_113_p N_A1_c_338_n 0.00452893f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_113_p N_A1_c_339_n 9.12852e-19 $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_113_p A1 0.00401739f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_113_p N_A1_c_343_n 4.68028e-19 $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_82_n N_VPWR_M1009_d 0.00664553f $X=1.08 $Y=1.835 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_83_n N_VPWR_M1009_d 0.00387091f $X=1.485 $Y=1.92 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_128_p N_VPWR_M1009_d 0.00283359f $X=1.165 $Y=1.92 $X2=0
+ $Y2=0
cc_116 N_A_79_21#_M1006_g N_VPWR_c_437_n 0.00450113f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_79_21#_M1009_g N_VPWR_c_438_n 0.00441646f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_79_21#_c_83_n N_VPWR_c_438_n 0.0115988f $X=1.485 $Y=1.92 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_128_p N_VPWR_c_438_n 0.0119477f $X=1.165 $Y=1.92 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_94_p N_VPWR_c_438_n 0.00582421f $X=1.57 $Y=2.255 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_95_p N_VPWR_c_438_n 0.0138777f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_122 N_A_79_21#_M1006_g N_VPWR_c_440_n 0.00541359f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_M1009_g N_VPWR_c_440_n 0.00571722f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_c_128_p N_VPWR_c_440_n 2.56506e-19 $X=1.165 $Y=1.92 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_83_n N_VPWR_c_441_n 0.00199439f $X=1.485 $Y=1.92 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_95_p N_VPWR_c_441_n 0.00780487f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_104_p N_VPWR_c_441_n 0.0538314f $X=2.63 $Y=2.34 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1005_d N_VPWR_c_435_n 0.00337207f $X=2.395 $Y=1.845 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_M1006_g N_VPWR_c_435_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_79_21#_M1009_g N_VPWR_c_435_n 0.0106088f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_83_n N_VPWR_c_435_n 0.00461221f $X=1.485 $Y=1.92 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_128_p N_VPWR_c_435_n 0.00149576f $X=1.165 $Y=1.92 $X2=0
+ $Y2=0
cc_133 N_A_79_21#_c_95_p N_VPWR_c_435_n 0.00617983f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_104_p N_VPWR_c_435_n 0.0407251f $X=2.63 $Y=2.34 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_74_n N_X_c_498_n 0.00437631f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_74_n N_X_c_499_n 0.00247572f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_78_n N_X_c_499_n 0.00156696f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_79_21#_M1006_g N_X_c_501_n 0.00351251f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_79_21#_M1009_g N_X_c_501_n 0.00371318f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_78_n N_X_c_501_n 0.00159703f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_74_n N_X_c_496_n 0.0076095f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_79_21#_M1006_g N_X_c_496_n 0.00984046f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_75_n N_X_c_496_n 0.00184881f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_79_21#_M1009_g N_X_c_496_n 0.00203892f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_82_n N_X_c_496_n 0.0104184f $X=1.08 $Y=1.835 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_77_n N_X_c_496_n 0.0234482f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_78_n N_X_c_496_n 0.0245558f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_79_n N_X_c_496_n 0.00726529f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_79_21#_M1006_g X 0.00825361f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_79_21#_M1009_g X 0.0087236f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_94_p X 0.00388105f $X=1.57 $Y=2.255 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_83_n A_306_369# 0.0016033f $X=1.485 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_79_21#_c_94_p A_306_369# 0.00412407f $X=1.57 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_79_21#_c_95_p A_306_369# 7.2174e-19 $X=1.655 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_79_21#_c_104_p A_306_369# 0.0166683f $X=2.63 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_79_21#_c_76_n N_VGND_M1011_d 0.00255482f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_170_p N_VGND_M1011_d 0.00230163f $X=1.165 $Y=0.72 $X2=0
+ $Y2=0
cc_158 N_A_79_21#_c_79_n N_VGND_M1011_d 0.00117765f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_74_n N_VGND_c_533_n 0.00312028f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_79_21#_c_74_n N_VGND_c_534_n 4.79856e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_75_n N_VGND_c_534_n 0.0071592f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_76_n N_VGND_c_534_n 0.00515539f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_170_p N_VGND_c_534_n 0.0120512f $X=1.165 $Y=0.72 $X2=0 $Y2=0
cc_164 N_A_79_21#_c_77_n N_VGND_c_534_n 0.00132593f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_78_n N_VGND_c_534_n 2.49234e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_74_n N_VGND_c_536_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_75_n N_VGND_c_536_n 0.0046653f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_76_n N_VGND_c_537_n 0.00260098f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_89_p N_VGND_c_537_n 0.00781925f $X=1.605 $Y=0.38 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_113_p N_VGND_c_537_n 0.0530528f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_171 N_A_79_21#_M1008_d N_VGND_c_539_n 0.00680618f $X=1.915 $Y=0.235 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_c_74_n N_VGND_c_539_n 0.0104557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_79_21#_c_75_n N_VGND_c_539_n 0.00789179f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_76_n N_VGND_c_539_n 0.00447974f $X=1.435 $Y=0.72 $X2=0 $Y2=0
cc_175 N_A_79_21#_c_170_p N_VGND_c_539_n 8.57032e-19 $X=1.165 $Y=0.72 $X2=0
+ $Y2=0
cc_176 N_A_79_21#_c_89_p N_VGND_c_539_n 0.00634027f $X=1.605 $Y=0.38 $X2=0 $Y2=0
cc_177 N_A_79_21#_c_113_p N_VGND_c_539_n 0.040112f $X=2.565 $Y=0.38 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_76_n A_288_47# 2.68783e-19 $X=1.435 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_79_21#_c_88_p A_288_47# 0.00193592f $X=1.52 $Y=0.635 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_79_21#_c_89_p A_288_47# 0.00114114f $X=1.605 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_79_21#_c_113_p A_288_47# 0.00493536f $X=2.565 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_257_199#_c_205_n N_A0_M1001_g 0.0125485f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_183 N_A_257_199#_M1004_g A0 7.18533e-19 $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_257_199#_c_196_n A0 0.0141669f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_257_199#_c_197_n A0 0.00239318f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_257_199#_c_202_n A0 0.0215416f $X=1.825 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A_257_199#_c_205_n A0 0.0212354f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_188 N_A_257_199#_c_205_n A0 0.042641f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_189 N_A_257_199#_c_196_n N_A0_c_287_n 3.23688e-19 $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_257_199#_c_197_n N_A0_c_287_n 0.00601779f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_257_199#_c_202_n N_A0_c_287_n 0.00251637f $X=1.825 $Y=1.58 $X2=0
+ $Y2=0
cc_192 N_A_257_199#_M1004_g N_A0_c_288_n 0.0323878f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A_257_199#_c_205_n N_A0_c_289_n 0.00103148f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_194 N_A_257_199#_M1012_g N_A1_M1005_g 0.0154518f $X=1.455 $Y=2.165 $X2=0
+ $Y2=0
cc_195 N_A_257_199#_c_197_n N_A1_M1005_g 0.00289638f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_257_199#_c_202_n N_A1_M1005_g 0.00246702f $X=1.825 $Y=1.58 $X2=0
+ $Y2=0
cc_197 N_A_257_199#_c_204_n N_A1_M1005_g 0.00374475f $X=1.91 $Y=1.835 $X2=0
+ $Y2=0
cc_198 N_A_257_199#_c_205_n N_A1_M1005_g 0.0132249f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_199 N_A_257_199#_c_198_n A1 0.00405973f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_200 N_A_257_199#_c_198_n A1 5.69346e-19 $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_201 N_A_257_199#_c_198_n N_S_M1010_g 6.08856e-19 $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_257_199#_c_205_n N_S_M1003_g 0.0162198f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_203 N_A_257_199#_c_198_n N_S_M1003_g 0.00109105f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_204 N_A_257_199#_c_207_n N_S_M1003_g 8.41605e-19 $X=3.88 $Y=2 $X2=0 $Y2=0
cc_205 N_A_257_199#_c_198_n N_S_M1013_g 0.0162888f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_206 N_A_257_199#_c_205_n N_S_M1000_g 0.012927f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_207 N_A_257_199#_c_198_n N_S_M1000_g 0.0168146f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_208 N_A_257_199#_c_207_n N_S_M1000_g 0.00673256f $X=3.88 $Y=2 $X2=0 $Y2=0
cc_209 N_A_257_199#_c_205_n S 0.0136816f $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_210 N_A_257_199#_c_198_n S 0.0646093f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_211 N_A_257_199#_c_205_n N_S_c_393_n 3.29564e-19 $X=3.715 $Y=1.92 $X2=0 $Y2=0
cc_212 N_A_257_199#_c_198_n N_S_c_393_n 0.0117966f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_213 N_A_257_199#_c_205_n N_VPWR_M1003_d 0.00161592f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_214 N_A_257_199#_M1012_g N_VPWR_c_438_n 0.00677196f $X=1.455 $Y=2.165 $X2=0
+ $Y2=0
cc_215 N_A_257_199#_c_205_n N_VPWR_c_439_n 0.012179f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_216 N_A_257_199#_M1012_g N_VPWR_c_441_n 0.00415313f $X=1.455 $Y=2.165 $X2=0
+ $Y2=0
cc_217 N_A_257_199#_c_205_n N_VPWR_c_441_n 0.00658059f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_218 N_A_257_199#_c_205_n N_VPWR_c_442_n 0.00208295f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_219 N_A_257_199#_c_207_n N_VPWR_c_442_n 0.021418f $X=3.88 $Y=2 $X2=0 $Y2=0
cc_220 N_A_257_199#_M1000_d N_VPWR_c_435_n 0.00217517f $X=3.735 $Y=1.845 $X2=0
+ $Y2=0
cc_221 N_A_257_199#_M1012_g N_VPWR_c_435_n 0.00691693f $X=1.455 $Y=2.165 $X2=0
+ $Y2=0
cc_222 N_A_257_199#_c_205_n N_VPWR_c_435_n 0.0190896f $X=3.715 $Y=1.92 $X2=0
+ $Y2=0
cc_223 N_A_257_199#_c_207_n N_VPWR_c_435_n 0.0126651f $X=3.88 $Y=2 $X2=0 $Y2=0
cc_224 N_A_257_199#_M1012_g X 6.93109e-19 $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_225 N_A_257_199#_c_205_n A_306_369# 0.00295934f $X=3.715 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_226 N_A_257_199#_c_232_n A_306_369# 0.00511624f $X=1.995 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_227 N_A_257_199#_c_205_n A_591_369# 0.0018249f $X=3.715 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_228 N_A_257_199#_M1004_g N_VGND_c_534_n 0.00310635f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_257_199#_M1004_g N_VGND_c_537_n 0.00423121f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_230 N_A_257_199#_c_198_n N_VGND_c_538_n 0.0210771f $X=3.88 $Y=0.42 $X2=0
+ $Y2=0
cc_231 N_A_257_199#_M1013_d N_VGND_c_539_n 0.00217517f $X=3.735 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_257_199#_M1004_g N_VGND_c_539_n 0.00594789f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_233 N_A_257_199#_c_198_n N_VGND_c_539_n 0.0124954f $X=3.88 $Y=0.42 $X2=0
+ $Y2=0
cc_234 N_A0_M1001_g N_A1_M1005_g 0.0285362f $X=2.88 $Y=2.165 $X2=0 $Y2=0
cc_235 A0 N_A1_M1005_g 0.0300135f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A0_c_289_n N_A1_M1005_g 0.0155275f $X=2.88 $Y=1.42 $X2=0 $Y2=0
cc_237 A0 N_A1_c_338_n 0.00661777f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_238 A0 N_A1_c_338_n 0.00611141f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_239 A0 N_A1_c_339_n 0.00613143f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_240 N_A0_c_287_n N_A1_c_339_n 0.0110204f $X=1.9 $Y=0.93 $X2=0 $Y2=0
cc_241 N_A0_c_287_n N_A1_M1002_g 3.75339e-19 $X=1.9 $Y=0.93 $X2=0 $Y2=0
cc_242 A0 A1 0.0211163f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_243 A0 A1 0.0235718f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_244 N_A0_c_287_n A1 2.08447e-19 $X=1.9 $Y=0.93 $X2=0 $Y2=0
cc_245 N_A0_c_289_n A1 0.00114405f $X=2.88 $Y=1.42 $X2=0 $Y2=0
cc_246 A0 N_A1_c_343_n 5.73679e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_247 A0 N_A1_c_343_n 0.00119563f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_248 N_A0_c_287_n N_A1_c_343_n 0.00169542f $X=1.9 $Y=0.93 $X2=0 $Y2=0
cc_249 N_A0_c_289_n N_A1_c_343_n 0.0212283f $X=2.88 $Y=1.42 $X2=0 $Y2=0
cc_250 N_A0_M1001_g N_S_M1003_g 0.0418775f $X=2.88 $Y=2.165 $X2=0 $Y2=0
cc_251 A0 S 0.0188995f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_252 A0 N_S_c_393_n 0.00270151f $X=2.91 $Y=1.445 $X2=0 $Y2=0
cc_253 N_A0_c_289_n N_S_c_393_n 0.0418775f $X=2.88 $Y=1.42 $X2=0 $Y2=0
cc_254 N_A0_M1001_g N_VPWR_c_441_n 0.00436487f $X=2.88 $Y=2.165 $X2=0 $Y2=0
cc_255 N_A0_M1001_g N_VPWR_c_435_n 0.00622759f $X=2.88 $Y=2.165 $X2=0 $Y2=0
cc_256 N_A0_c_288_n N_VGND_c_537_n 0.00366111f $X=1.9 $Y=0.765 $X2=0 $Y2=0
cc_257 N_A0_c_288_n N_VGND_c_539_n 0.00672884f $X=1.9 $Y=0.765 $X2=0 $Y2=0
cc_258 N_A1_M1002_g N_S_M1010_g 0.0289474f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_259 A1 N_S_M1010_g 0.00316198f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_260 A1 N_S_M1010_g 0.00255209f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_261 N_A1_c_343_n N_S_M1010_g 0.0169127f $X=2.79 $Y=0.94 $X2=0 $Y2=0
cc_262 A1 S 0.0159208f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_263 N_A1_c_343_n S 2.83278e-19 $X=2.79 $Y=0.94 $X2=0 $Y2=0
cc_264 N_A1_M1005_g N_VPWR_c_441_n 0.00366111f $X=2.32 $Y=2.165 $X2=0 $Y2=0
cc_265 N_A1_M1005_g N_VPWR_c_435_n 0.00643646f $X=2.32 $Y=2.165 $X2=0 $Y2=0
cc_266 N_A1_M1002_g N_VGND_c_537_n 0.00439206f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_267 A1 N_VGND_c_537_n 0.00538049f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_268 A1 N_VGND_c_537_n 0.00237968f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_269 N_A1_M1002_g N_VGND_c_539_n 0.00744578f $X=2.815 $Y=0.445 $X2=0 $Y2=0
cc_270 A1 N_VGND_c_539_n 0.00640177f $X=2.91 $Y=0.425 $X2=0 $Y2=0
cc_271 A1 N_VGND_c_539_n 0.00411784f $X=2.91 $Y=0.765 $X2=0 $Y2=0
cc_272 A1 A_578_47# 0.00558936f $X=2.91 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_273 N_S_M1003_g N_VPWR_c_439_n 0.00298136f $X=3.24 $Y=2.165 $X2=0 $Y2=0
cc_274 N_S_M1000_g N_VPWR_c_439_n 0.00281335f $X=3.66 $Y=2.165 $X2=0 $Y2=0
cc_275 N_S_M1003_g N_VPWR_c_441_n 0.00436487f $X=3.24 $Y=2.165 $X2=0 $Y2=0
cc_276 N_S_M1000_g N_VPWR_c_442_n 0.00427495f $X=3.66 $Y=2.165 $X2=0 $Y2=0
cc_277 N_S_M1003_g N_VPWR_c_435_n 0.00567152f $X=3.24 $Y=2.165 $X2=0 $Y2=0
cc_278 N_S_M1000_g N_VPWR_c_435_n 0.00668913f $X=3.66 $Y=2.165 $X2=0 $Y2=0
cc_279 N_S_M1010_g N_VGND_c_535_n 0.00281288f $X=3.24 $Y=0.445 $X2=0 $Y2=0
cc_280 N_S_M1013_g N_VGND_c_535_n 0.00281288f $X=3.66 $Y=0.445 $X2=0 $Y2=0
cc_281 S N_VGND_c_535_n 0.0152508f $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_282 N_S_c_393_n N_VGND_c_535_n 4.13159e-19 $X=3.66 $Y=1.16 $X2=0 $Y2=0
cc_283 N_S_M1010_g N_VGND_c_537_n 0.00585385f $X=3.24 $Y=0.445 $X2=0 $Y2=0
cc_284 N_S_M1013_g N_VGND_c_538_n 0.00564131f $X=3.66 $Y=0.445 $X2=0 $Y2=0
cc_285 N_S_M1010_g N_VGND_c_539_n 0.0106164f $X=3.24 $Y=0.445 $X2=0 $Y2=0
cc_286 N_S_M1013_g N_VGND_c_539_n 0.0109824f $X=3.66 $Y=0.445 $X2=0 $Y2=0
cc_287 S N_VGND_c_539_n 7.73929e-19 $X=3.37 $Y=0.765 $X2=0 $Y2=0
cc_288 N_VPWR_c_435_n N_X_M1006_s 0.00215201f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_438_n X 0.0195756f $X=1.15 $Y=2.34 $X2=0 $Y2=0
cc_290 N_VPWR_c_440_n X 0.0175403f $X=1.025 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_435_n X 0.0115429f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_435_n A_306_369# 0.00586504f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_293 N_VPWR_c_435_n A_591_369# 0.00269901f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_294 N_VPWR_c_437_n N_VGND_c_533_n 0.0086775f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_295 N_X_c_498_n N_VGND_c_536_n 0.0150329f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_296 N_X_M1007_s N_VGND_c_539_n 0.0038878f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_297 N_X_c_498_n N_VGND_c_539_n 0.00932112f $X=0.68 $Y=0.42 $X2=0 $Y2=0
cc_298 N_VGND_c_539_n A_288_47# 0.00263843f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_299 N_VGND_c_539_n A_578_47# 0.00503489f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

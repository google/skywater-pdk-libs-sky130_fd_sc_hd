* File: sky130_fd_sc_hd__nand4_1.spice.SKY130_FD_SC_HD__NAND4_1.pxi
* Created: Thu Aug 27 14:30:06 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4_1%D N_D_c_44_n N_D_M1007_g N_D_M1005_g D N_D_c_46_n
+ PM_SKY130_FD_SC_HD__NAND4_1%D
x_PM_SKY130_FD_SC_HD__NAND4_1%C N_C_c_69_n N_C_M1002_g N_C_M1001_g C C C
+ N_C_c_71_n N_C_c_72_n PM_SKY130_FD_SC_HD__NAND4_1%C
x_PM_SKY130_FD_SC_HD__NAND4_1%B N_B_M1004_g N_B_M1000_g N_B_c_108_n N_B_c_109_n
+ N_B_c_110_n B N_B_c_111_n PM_SKY130_FD_SC_HD__NAND4_1%B
x_PM_SKY130_FD_SC_HD__NAND4_1%A N_A_c_151_n N_A_M1006_g N_A_M1003_g A A
+ N_A_c_153_n PM_SKY130_FD_SC_HD__NAND4_1%A
x_PM_SKY130_FD_SC_HD__NAND4_1%VPWR N_VPWR_M1005_s N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n N_VPWR_c_183_n N_VPWR_c_184_n
+ N_VPWR_c_185_n N_VPWR_c_186_n VPWR N_VPWR_c_187_n N_VPWR_c_179_n
+ PM_SKY130_FD_SC_HD__NAND4_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND4_1%Y N_Y_M1006_d N_Y_M1005_d N_Y_M1000_d N_Y_c_218_n
+ N_Y_c_219_n N_Y_c_224_n N_Y_c_255_n N_Y_c_215_n N_Y_c_236_n Y N_Y_c_216_n
+ PM_SKY130_FD_SC_HD__NAND4_1%Y
x_PM_SKY130_FD_SC_HD__NAND4_1%VGND N_VGND_M1007_s N_VGND_c_261_n N_VGND_c_262_n
+ VGND N_VGND_c_263_n N_VGND_c_264_n PM_SKY130_FD_SC_HD__NAND4_1%VGND
cc_1 VNB N_D_c_44_n 0.0212957f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB D 0.0139673f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_D_c_46_n 0.0355062f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_C_c_69_n 0.0164311f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB C 0.00226512f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_C_c_71_n 0.0213808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_C_c_72_n 0.00235574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_108_n 0.00109375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_109_n 0.00208581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_c_110_n 0.0232548f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_11 VNB N_B_c_111_n 0.016344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_c_151_n 0.0221199f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB A 0.0133408f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_A_c_153_n 0.0367295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_179_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_215_n 0.00261864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_216_n 0.0249997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_261_n 0.0102727f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_19 VNB N_VGND_c_262_n 0.0262359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB N_VGND_c_263_n 0.0492405f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_264_n 0.141941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_D_M1005_g 0.0263149f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_23 VPB D 0.00475375f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_24 VPB N_D_c_46_n 0.0094694f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_25 VPB N_C_M1001_g 0.0191664f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_26 VPB N_C_c_71_n 0.00397839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_C_c_72_n 0.0016008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_B_M1000_g 0.0197878f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_29 VPB N_B_c_109_n 9.48942e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_B_c_110_n 0.00399403f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_31 VPB N_A_M1003_g 0.0219896f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB A 0.0152386f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_c_153_n 0.0124663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_180_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_35 VPB N_VPWR_c_181_n 0.0429032f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_36 VPB N_VPWR_c_182_n 0.00415222f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_183_n 0.0109102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_184_n 0.0298835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_185_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_186_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_187_n 0.0200551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_179_n 0.0428917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_215_n 0.00132625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 N_D_c_44_n N_C_c_69_n 0.0353923f $X=0.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_45 N_D_M1005_g N_C_M1001_g 0.0151563f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_46 N_D_c_44_n C 0.00513227f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_47 D N_C_c_71_n 2.49652e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_48 N_D_c_46_n N_C_c_71_n 0.0207259f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_49 D N_C_c_72_n 0.023096f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_50 N_D_c_46_n N_C_c_72_n 0.00264953f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_51 N_D_M1005_g N_VPWR_c_181_n 0.00321781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_52 D N_VPWR_c_181_n 0.0191671f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_53 N_D_c_46_n N_VPWR_c_181_n 0.00171514f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_54 N_D_M1005_g N_VPWR_c_185_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_55 N_D_M1005_g N_VPWR_c_179_n 0.0104829f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_56 N_D_M1005_g N_Y_c_218_n 0.00338192f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_57 N_D_M1005_g N_Y_c_219_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_58 N_D_c_44_n N_VGND_c_262_n 0.0141323f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_59 D N_VGND_c_262_n 0.0210629f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_60 N_D_c_46_n N_VGND_c_262_n 0.00195936f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_61 N_D_c_44_n N_VGND_c_263_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 N_D_c_44_n N_VGND_c_264_n 0.00799591f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 N_C_M1001_g N_B_M1000_g 0.0292916f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_64 N_C_c_69_n N_B_c_108_n 0.00123452f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_65 C N_B_c_108_n 0.006646f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_66 N_C_c_71_n N_B_c_109_n 0.00197607f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_67 N_C_c_72_n N_B_c_109_n 0.0263533f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_68 N_C_c_71_n N_B_c_110_n 0.020191f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_69 N_C_c_72_n N_B_c_110_n 3.16067e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_70 N_C_c_71_n B 5.13678e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C_c_69_n N_B_c_111_n 0.0392711f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_72 N_C_M1001_g N_VPWR_c_182_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_73 N_C_M1001_g N_VPWR_c_185_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_74 N_C_M1001_g N_VPWR_c_179_n 0.00955595f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_75 N_C_M1001_g N_Y_c_218_n 8.84614e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_76 N_C_c_71_n N_Y_c_218_n 0.00122405f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_c_72_n N_Y_c_218_n 0.0183056f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_M1001_g N_Y_c_219_n 0.00983512f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_79 N_C_M1001_g N_Y_c_224_n 0.0106747f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_80 N_C_c_71_n N_Y_c_224_n 0.00123493f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_81 N_C_c_72_n N_Y_c_224_n 0.00891084f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C_c_69_n N_VGND_c_262_n 0.00151754f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_83 N_C_c_69_n N_VGND_c_263_n 0.00585385f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_84 C N_VGND_c_263_n 0.0101172f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_85 N_C_c_69_n N_VGND_c_264_n 0.0108681f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_86 C N_VGND_c_264_n 0.00802479f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_87 C A_109_47# 0.00607973f $X=0.61 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_88 B N_A_c_151_n 7.81004e-19 $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_89 N_B_c_111_n N_A_c_151_n 0.030612f $X=1.37 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_90 N_B_M1000_g N_A_M1003_g 0.010807f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B_c_109_n N_A_c_153_n 3.15088e-19 $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B_c_110_n N_A_c_153_n 0.02024f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_M1000_g N_VPWR_c_182_n 0.00268723f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B_M1000_g N_VPWR_c_187_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_VPWR_c_179_n 0.0107321f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B_M1000_g N_Y_c_219_n 6.26017e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B_M1000_g N_Y_c_224_n 0.0128868f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B_c_109_n N_Y_c_224_n 0.0156236f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_99 B N_Y_c_224_n 0.00347602f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_100 N_B_M1000_g N_Y_c_215_n 0.00233229f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B_c_108_n N_Y_c_215_n 0.0060434f $X=1.247 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B_c_109_n N_Y_c_215_n 0.0246541f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_110_n N_Y_c_215_n 0.00190138f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_c_111_n N_Y_c_215_n 7.5826e-19 $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_109_n N_Y_c_236_n 0.00322248f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_106 N_B_c_110_n N_Y_c_236_n 0.00367907f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_107 B N_Y_c_216_n 0.0434018f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_108 N_B_c_111_n N_Y_c_216_n 0.00518446f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_109 B N_VGND_c_263_n 0.016572f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_110 N_B_c_111_n N_VGND_c_263_n 0.0041935f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_111 B N_VGND_c_264_n 0.0125298f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_112 N_B_c_111_n N_VGND_c_264_n 0.00681121f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_108_n A_193_47# 6.5878e-19 $X=1.247 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_114 B A_193_47# 0.00523732f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_115 A N_VPWR_M1003_d 0.0052728f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A_M1003_g N_VPWR_c_184_n 0.00452839f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_117 A N_VPWR_c_184_n 0.0197361f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_c_153_n N_VPWR_c_184_n 0.00260772f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_M1003_g N_VPWR_c_187_n 0.00585385f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1003_g N_VPWR_c_179_n 0.0116954f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_c_151_n N_Y_c_215_n 0.00933112f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_M1003_g N_Y_c_215_n 0.00380538f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_123 A N_Y_c_215_n 0.0342212f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_153_n N_Y_c_215_n 0.00842855f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_Y_c_236_n 0.00653595f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_126 A N_Y_c_236_n 0.0130944f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_c_151_n N_Y_c_216_n 0.0182263f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_128 A N_Y_c_216_n 0.0206713f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A_c_153_n N_Y_c_216_n 0.00518508f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_c_151_n N_VGND_c_263_n 0.00357668f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_151_n N_VGND_c_264_n 0.00638972f $X=1.79 $Y=0.995 $X2=0 $Y2=0
cc_132 N_VPWR_c_179_n N_Y_M1005_d 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_179_n N_Y_M1000_d 0.0026338f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_185_n N_Y_c_219_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_c_179_n N_Y_c_219_n 0.0122217f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_136 N_VPWR_M1001_d N_Y_c_224_n 0.00452985f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_137 N_VPWR_c_182_n N_Y_c_224_n 0.0126919f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_138 N_VPWR_c_187_n N_Y_c_255_n 0.0191632f $X=1.915 $Y=2.72 $X2=0 $Y2=0
cc_139 N_VPWR_c_179_n N_Y_c_255_n 0.0126319f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_140 N_VPWR_c_181_n N_VGND_c_262_n 7.14544e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_141 N_Y_c_216_n N_VGND_c_263_n 0.0440555f $X=2 $Y=0.38 $X2=0 $Y2=0
cc_142 N_Y_M1006_d N_VGND_c_264_n 0.00242111f $X=1.865 $Y=0.235 $X2=0 $Y2=0
cc_143 N_Y_c_216_n N_VGND_c_264_n 0.0258385f $X=2 $Y=0.38 $X2=0 $Y2=0
cc_144 N_Y_c_216_n A_277_47# 0.0087441f $X=2 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_145 N_VGND_c_264_n A_109_47# 0.00416909f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
cc_146 N_VGND_c_264_n A_193_47# 0.00344225f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
cc_147 N_VGND_c_264_n A_277_47# 0.0073712f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdfxbp_1.pex.spice
* Created: Thu Aug 27 14:47:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%CLK 1 2 3 5 6 8 11 13
c42 1 0 2.71124e-20 $X=0.31 $Y=1.325
r43 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r44 9 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.31 $Y=1.665
+ $X2=0.47 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r47 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r50 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_27_47# 1 2 9 13 17 19 20 25 29 31 35 39
+ 43 44 45 49 50 52 55 56 57 58 59 60 69 74 77 78 79 81 85
c246 85 0 1.77381e-19 $X=6.65 $Y=1.41
c247 52 0 8.70797e-20 $X=0.76 $Y=1.235
c248 50 0 1.8506e-19 $X=0.73 $Y=1.795
c249 45 0 5.65522e-20 $X=0.615 $Y=1.88
c250 29 0 4.21632e-20 $X=6.655 $Y=2.275
c251 19 0 1.57835e-19 $X=4.965 $Y=1.32
r252 84 86 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.41
+ $X2=6.65 $Y2=1.575
r253 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.65
+ $Y=1.41 $X2=6.65 $Y2=1.41
r254 81 84 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.65 $Y=1.32 $X2=6.65
+ $Y2=1.41
r255 77 80 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.74
+ $X2=5.1 $Y2=1.905
r256 77 79 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.74
+ $X2=5.1 $Y2=1.575
r257 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.74 $X2=5.1 $Y2=1.74
r258 70 85 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=6.66 $Y=1.87
+ $X2=6.66 $Y2=1.41
r259 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.66 $Y=1.87
+ $X2=6.66 $Y2=1.87
r260 66 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.25 $Y=1.87
+ $X2=5.25 $Y2=1.87
r261 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r262 60 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.395 $Y=1.87
+ $X2=5.25 $Y2=1.87
r263 59 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.515 $Y=1.87
+ $X2=6.66 $Y2=1.87
r264 59 60 1.38614 $w=1.4e-07 $l=1.12e-06 $layer=MET1_cond $X=6.515 $Y=1.87
+ $X2=5.395 $Y2=1.87
r265 58 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r266 57 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.105 $Y=1.87
+ $X2=5.25 $Y2=1.87
r267 57 58 5.23514 $w=1.4e-07 $l=4.23e-06 $layer=MET1_cond $X=5.105 $Y=1.87
+ $X2=0.875 $Y2=1.87
r268 53 74 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.76 $Y=1.235
+ $X2=0.89 $Y2=1.235
r269 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.235 $X2=0.76 $Y2=1.235
r270 50 63 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.88
r271 50 52 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.795
+ $X2=0.73 $Y2=1.235
r272 49 56 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=0.97
r273 49 52 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.73 $Y=1.085
+ $X2=0.73 $Y2=1.235
r274 47 56 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.712 $Y=0.805
+ $X2=0.712 $Y2=0.97
r275 46 55 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r276 45 63 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.73 $Y2=1.88
r277 45 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=1.88
+ $X2=0.345 $Y2=1.88
r278 43 47 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.712 $Y2=0.805
r279 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=0.72
+ $X2=0.345 $Y2=0.72
r280 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r281 37 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r282 33 35 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.3 $Y=1.245
+ $X2=7.3 $Y2=0.415
r283 32 81 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.785 $Y=1.32
+ $X2=6.65 $Y2=1.32
r284 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=1.32
+ $X2=7.3 $Y2=1.245
r285 31 32 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=7.225 $Y=1.32
+ $X2=6.785 $Y2=1.32
r286 29 86 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.655 $Y=2.275
+ $X2=6.655 $Y2=1.575
r287 25 80 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.04 $Y=2.275
+ $X2=5.04 $Y2=1.905
r288 21 79 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.04 $Y=1.395
+ $X2=5.04 $Y2=1.575
r289 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.965 $Y=1.32
+ $X2=5.04 $Y2=1.395
r290 19 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.965 $Y=1.32
+ $X2=4.655 $Y2=1.32
r291 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=1.245
+ $X2=4.655 $Y2=1.32
r292 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.58 $Y=1.245
+ $X2=4.58 $Y2=0.415
r293 11 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r294 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r295 7 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r296 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r297 2 55 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r298 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%SCE 3 7 9 13 17 19 21 22 24 26 30 31 35 36
c117 26 0 1.66295e-19 $X=3.065 $Y=0.7
c118 24 0 1.76484e-19 $X=2.455 $Y=0.7
r119 40 41 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.58
+ $X2=1.845 $Y2=1.655
r120 34 36 6.65455 $w=1.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.542 $Y=0.615
+ $X2=2.542 $Y2=0.51
r121 34 35 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.542 $Y=0.615
+ $X2=2.542 $Y2=0.7
r122 31 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.95
+ $X2=3.15 $Y2=0.785
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=0.95 $X2=3.15 $Y2=0.95
r124 28 30 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0.785
+ $X2=3.15 $Y2=0.95
r125 27 35 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.63 $Y=0.7
+ $X2=2.542 $Y2=0.7
r126 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.065 $Y=0.7
+ $X2=3.15 $Y2=0.785
r127 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.065 $Y=0.7
+ $X2=2.63 $Y2=0.7
r128 25 33 1.50975 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.01 $Y=0.7
+ $X2=1.885 $Y2=0.7
r129 24 35 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=2.455 $Y=0.7
+ $X2=2.542 $Y2=0.7
r130 24 25 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.455 $Y=0.7
+ $X2=2.01 $Y2=0.7
r131 22 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.845 $Y=1.52
+ $X2=1.845 $Y2=1.58
r132 22 39 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.845 $Y=1.52
+ $X2=1.845 $Y2=1.385
r133 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.52 $X2=1.845 $Y2=1.52
r134 19 33 11.5378 $w=1.94e-07 $l=1.98997e-07 $layer=LI1_cond $X=1.845 $Y=0.88
+ $X2=1.885 $Y2=0.7
r135 19 21 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.845 $Y=0.88
+ $X2=1.845 $Y2=1.52
r136 17 43 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.21 $Y=0.445
+ $X2=3.21 $Y2=0.785
r137 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.25 $Y=1.655
+ $X2=2.25 $Y2=2.165
r138 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.58
+ $X2=1.845 $Y2=1.58
r139 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.175 $Y=1.58
+ $X2=2.25 $Y2=1.655
r140 9 10 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.175 $Y=1.58
+ $X2=2.01 $Y2=1.58
r141 7 41 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.83 $Y=2.165
+ $X2=1.83 $Y2=1.655
r142 3 39 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.83 $Y=0.445 $X2=1.83
+ $Y2=1.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_299_47# 1 2 9 13 16 19 21 24 25 28 32 34
+ 38 39 41 43 44
c126 43 0 1.84493e-19 $X=3.17 $Y=1.52
c127 41 0 1.81307e-19 $X=2.185 $Y=1.967
c128 39 0 1.12087e-19 $X=2.28 $Y=1.04
c129 24 0 1.59836e-19 $X=2.185 $Y=1.86
c130 9 0 1.20015e-19 $X=2.34 $Y=0.445
r131 44 52 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.52
+ $X2=3.17 $Y2=1.685
r132 43 46 9.59627 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.157 $Y=1.52
+ $X2=3.157 $Y2=1.685
r133 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.52 $X2=3.17 $Y2=1.52
r134 39 48 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.28 $Y=1.04
+ $X2=2.28 $Y2=0.905
r135 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.04 $X2=2.28 $Y2=1.04
r136 35 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.185 $Y=1.04
+ $X2=2.28 $Y2=1.04
r137 29 32 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.505 $Y=0.42
+ $X2=1.62 $Y2=0.42
r138 28 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.145 $Y=1.86
+ $X2=3.145 $Y2=1.685
r139 26 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=1.967
+ $X2=2.185 $Y2=1.967
r140 25 28 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.06 $Y=1.967
+ $X2=3.145 $Y2=1.86
r141 25 26 42.3456 $w=2.13e-07 $l=7.9e-07 $layer=LI1_cond $X=3.06 $Y=1.967
+ $X2=2.27 $Y2=1.967
r142 24 41 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.185 $Y=1.86
+ $X2=2.185 $Y2=1.967
r143 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=1.125
+ $X2=2.185 $Y2=1.04
r144 23 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.185 $Y=1.125
+ $X2=2.185 $Y2=1.86
r145 22 34 1.54683 $w=2.15e-07 $l=1.43e-07 $layer=LI1_cond $X=1.705 $Y=1.967
+ $X2=1.562 $Y2=1.967
r146 21 41 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=1.967
+ $X2=2.185 $Y2=1.967
r147 21 22 21.1728 $w=2.13e-07 $l=3.95e-07 $layer=LI1_cond $X=2.1 $Y=1.967
+ $X2=1.705 $Y2=1.967
r148 17 34 4.92743 $w=2.27e-07 $l=1.08e-07 $layer=LI1_cond $X=1.562 $Y=2.075
+ $X2=1.562 $Y2=1.967
r149 17 19 4.04366 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=1.562 $Y=2.075
+ $X2=1.562 $Y2=2.175
r150 16 34 4.92743 $w=2.27e-07 $l=1.32469e-07 $layer=LI1_cond $X=1.505 $Y=1.86
+ $X2=1.562 $Y2=1.967
r151 15 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.585
+ $X2=1.505 $Y2=0.42
r152 15 16 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=1.505 $Y=0.585
+ $X2=1.505 $Y2=1.86
r153 13 52 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.125 $Y=2.165
+ $X2=3.125 $Y2=1.685
r154 9 48 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.34 $Y=0.445
+ $X2=2.34 $Y2=0.905
r155 2 19 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=2.175
r156 1 32 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%D 3 7 9 12 13
c50 13 0 2.8857e-19 $X=2.69 $Y=1.52
r51 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.52
+ $X2=2.69 $Y2=1.685
r52 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.52
+ $X2=2.69 $Y2=1.355
r53 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.52 $X2=2.69 $Y2=1.52
r54 9 13 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=1.52 $X2=2.69
+ $Y2=1.52
r55 7 14 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.73 $Y=0.445
+ $X2=2.73 $Y2=1.355
r56 3 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.705 $Y=2.165
+ $X2=2.705 $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%SCD 3 7 9 12
c49 7 0 1.84493e-19 $X=3.59 $Y=2.165
c50 3 0 1.66295e-19 $X=3.59 $Y=0.445
r51 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.355
+ $X2=3.65 $Y2=1.52
r52 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.355
+ $X2=3.65 $Y2=1.19
r53 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.355 $X2=3.65 $Y2=1.355
r54 9 13 4.98366 $w=5.98e-07 $l=2.5e-07 $layer=LI1_cond $X=3.9 $Y=1.355 $X2=3.65
+ $Y2=1.355
r55 7 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.59 $Y=2.165
+ $X2=3.59 $Y2=1.52
r56 3 14 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.59 $Y=0.445
+ $X2=3.59 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_193_47# 1 2 9 13 14 16 19 23 24 27 28 32
+ 33 35 36 37 38 45 47 54 56 61 69
c212 61 0 1.77381e-19 $X=6.88 $Y=0.87
c213 37 0 1.57835e-19 $X=6.525 $Y=0.85
r214 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=0.87 $X2=6.88 $Y2=0.87
r215 58 61 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.785 $Y=0.87
+ $X2=6.88 $Y2=0.87
r216 54 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=0.87 $X2=5
+ $Y2=0.705
r217 48 62 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.67 $Y=0.87
+ $X2=6.88 $Y2=0.87
r218 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0.85
+ $X2=6.67 $Y2=0.85
r219 45 78 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.83 $Y=0.87
+ $X2=4.625 $Y2=0.87
r220 45 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5 $Y=0.87
+ $X2=5 $Y2=0.87
r221 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0.85
+ $X2=4.83 $Y2=0.85
r222 41 73 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=1.1 $Y=0.85
+ $X2=1.1 $Y2=1.96
r223 41 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.1 $Y=0.85 $X2=1.1
+ $Y2=0.51
r224 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=0.85 $X2=1.1
+ $Y2=0.85
r225 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=0.85
+ $X2=4.83 $Y2=0.85
r226 37 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.525 $Y=0.85
+ $X2=6.67 $Y2=0.85
r227 37 38 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=6.525 $Y=0.85
+ $X2=4.975 $Y2=0.85
r228 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=0.85
+ $X2=1.1 $Y2=0.85
r229 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=4.83 $Y2=0.85
r230 35 36 4.25742 $w=1.4e-07 $l=3.44e-06 $layer=MET1_cond $X=4.685 $Y=0.85
+ $X2=1.245 $Y2=0.85
r231 33 64 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=7.16 $Y=1.74
+ $X2=7.075 $Y2=1.74
r232 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.16
+ $Y=1.74 $X2=7.16 $Y2=1.74
r233 29 32 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.02 $Y=1.74
+ $X2=7.16 $Y2=1.74
r234 28 62 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.925 $Y=0.87
+ $X2=6.88 $Y2=0.87
r235 27 29 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.02 $Y=1.575
+ $X2=7.02 $Y2=1.74
r236 26 28 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.02 $Y=1.035
+ $X2=6.925 $Y2=0.87
r237 26 27 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.02 $Y=1.035
+ $X2=7.02 $Y2=1.575
r238 24 52 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.59 $Y=1.74
+ $X2=4.59 $Y2=1.875
r239 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.59
+ $Y=1.74 $X2=4.59 $Y2=1.74
r240 21 78 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=1.035
+ $X2=4.625 $Y2=0.87
r241 21 23 33.853 $w=2.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.625 $Y=1.035
+ $X2=4.625 $Y2=1.74
r242 17 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.075 $Y=1.875
+ $X2=7.075 $Y2=1.74
r243 17 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.075 $Y=1.875
+ $X2=7.075 $Y2=2.275
r244 14 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.785 $Y=0.705
+ $X2=6.785 $Y2=0.87
r245 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.785 $Y=0.705
+ $X2=6.785 $Y2=0.415
r246 13 56 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.06 $Y=0.415
+ $X2=5.06 $Y2=0.705
r247 9 52 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.575 $Y=2.275
+ $X2=4.575 $Y2=1.875
r248 2 73 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r249 1 69 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_1089_183# 1 2 9 13 15 18 21 23 29 30 32
+ 33 36
r95 35 36 5.54023 $w=2.61e-07 $l=3e-08 $layer=POLY_cond $X=5.52 $Y=0.93 $X2=5.55
+ $Y2=0.93
r96 32 33 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=2.3
+ $X2=6.35 $Y2=2.135
r97 27 36 24.0077 $w=2.61e-07 $l=1.3e-07 $layer=POLY_cond $X=5.68 $Y=0.93
+ $X2=5.55 $Y2=0.93
r98 26 29 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=0.93
+ $X2=5.765 $Y2=0.93
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=0.93 $X2=5.68 $Y2=0.93
r100 21 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.395 $Y=0.45
+ $X2=6.52 $Y2=0.45
r101 19 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.31 $Y=1.065
+ $X2=6.31 $Y2=0.915
r102 19 33 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.31 $Y=1.065
+ $X2=6.31 $Y2=2.135
r103 18 30 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.31 $Y=0.765
+ $X2=6.31 $Y2=0.915
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.31 $Y=0.535
+ $X2=6.395 $Y2=0.45
r105 17 18 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.31 $Y=0.535
+ $X2=6.31 $Y2=0.765
r106 15 30 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=0.915
+ $X2=6.31 $Y2=0.915
r107 15 29 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.225 $Y=0.915
+ $X2=5.765 $Y2=0.915
r108 11 36 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.55 $Y=0.795
+ $X2=5.55 $Y2=0.93
r109 11 13 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=5.55 $Y=0.795
+ $X2=5.55 $Y2=0.445
r110 7 35 15.717 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.52 $Y=1.065
+ $X2=5.52 $Y2=0.93
r111 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=5.52 $Y=1.065
+ $X2=5.52 $Y2=2.275
r112 2 32 600 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.735 $X2=6.39 $Y2=2.3
r113 1 23 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.235 $X2=6.52 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_930_413# 1 2 8 11 13 15 18 20 21 22 26 31
+ 33 35
c108 31 0 1.42307e-19 $X=5.34 $Y=1.315
r109 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=1.41 $X2=5.97 $Y2=1.41
r110 35 37 17.1405 $w=2.42e-07 $l=3.4e-07 $layer=LI1_cond $X=5.63 $Y=1.41
+ $X2=5.97 $Y2=1.41
r111 32 35 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=1.575
+ $X2=5.63 $Y2=1.41
r112 32 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.63 $Y=1.575
+ $X2=5.63 $Y2=2.19
r113 31 35 14.6198 $w=2.42e-07 $l=2.9e-07 $layer=LI1_cond $X=5.34 $Y=1.41
+ $X2=5.63 $Y2=1.41
r114 30 31 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.34 $Y=0.535
+ $X2=5.34 $Y2=1.315
r115 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.255 $Y=0.45
+ $X2=5.34 $Y2=0.535
r116 26 28 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.255 $Y=0.45
+ $X2=4.85 $Y2=0.45
r117 22 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.545 $Y=2.275
+ $X2=5.63 $Y2=2.19
r118 22 24 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.545 $Y=2.275
+ $X2=4.81 $Y2=2.275
r119 20 38 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.105 $Y=1.41
+ $X2=5.97 $Y2=1.41
r120 20 21 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=6.105 $Y=1.41
+ $X2=6.18 $Y2=1.41
r121 16 18 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.18 $Y=1.025
+ $X2=6.28 $Y2=1.025
r122 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.28 $Y=0.95
+ $X2=6.28 $Y2=1.025
r123 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.28 $Y=0.95
+ $X2=6.28 $Y2=0.555
r124 9 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.18 $Y=1.545
+ $X2=6.18 $Y2=1.41
r125 9 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=6.18 $Y=1.545
+ $X2=6.18 $Y2=2.11
r126 8 21 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.18 $Y=1.275
+ $X2=6.18 $Y2=1.41
r127 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.18 $Y=1.1 $X2=6.18
+ $Y2=1.025
r128 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.18 $Y=1.1 $X2=6.18
+ $Y2=1.275
r129 2 24 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=4.65
+ $Y=2.065 $X2=4.81 $Y2=2.275
r130 1 28 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.235 $X2=4.85 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_1517_315# 1 2 9 13 15 17 20 22 24 26 28
+ 31 34 35 36 39 43 47 50 52 55 56 58 59 60
c125 56 0 4.4412e-19 $X=9.135 $Y=1.16
c126 34 0 1.53472e-19 $X=10.047 $Y=1.515
r127 61 63 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.66 $Y=1.74
+ $X2=7.775 $Y2=1.74
r128 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.135
+ $Y=1.16 $X2=9.135 $Y2=1.16
r129 53 60 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=8.67 $Y=1.16
+ $X2=8.577 $Y2=1.16
r130 53 55 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.67 $Y=1.16
+ $X2=9.135 $Y2=1.16
r131 52 59 6.72893 $w=2.37e-07 $l=1.89222e-07 $layer=LI1_cond $X=8.577 $Y=1.575
+ $X2=8.525 $Y2=1.74
r132 51 60 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=8.577 $Y=1.325
+ $X2=8.577 $Y2=1.16
r133 51 52 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=8.577 $Y=1.325
+ $X2=8.577 $Y2=1.575
r134 50 60 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=8.577 $Y=0.995
+ $X2=8.577 $Y2=1.16
r135 50 58 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=8.577 $Y=0.995
+ $X2=8.577 $Y2=0.825
r136 45 59 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=8.525 $Y=1.905
+ $X2=8.525 $Y2=1.74
r137 45 47 1.78827 $w=2.88e-07 $l=4.5e-08 $layer=LI1_cond $X=8.525 $Y=1.905
+ $X2=8.525 $Y2=1.95
r138 41 58 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=0.66
+ $X2=8.505 $Y2=0.825
r139 41 43 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.505 $Y=0.66
+ $X2=8.505 $Y2=0.385
r140 39 63 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.84 $Y=1.74
+ $X2=7.775 $Y2=1.74
r141 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.84
+ $Y=1.74 $X2=7.84 $Y2=1.74
r142 36 59 0.189605 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=8.38 $Y=1.74
+ $X2=8.525 $Y2=1.74
r143 36 38 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.38 $Y=1.74
+ $X2=7.84 $Y2=1.74
r144 34 35 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=10.047 $Y=1.515
+ $X2=10.047 $Y2=1.665
r145 31 35 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=10.075 $Y=2.165
+ $X2=10.075 $Y2=1.665
r146 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.075 $Y=0.73
+ $X2=10.075 $Y2=0.445
r147 24 34 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.02 $Y=1.325
+ $X2=10.02 $Y2=1.515
r148 23 56 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=9.21 $Y=1.16
+ $X2=9.105 $Y2=1.16
r149 22 24 49.1818 $w=1.63e-07 $l=1.77989e-07 $layer=POLY_cond $X=10.047 $Y=1.16
+ $X2=10.02 $Y2=1.325
r150 22 26 127.544 $w=1.63e-07 $l=4.43779e-07 $layer=POLY_cond $X=10.047 $Y=1.16
+ $X2=10.075 $Y2=0.73
r151 22 23 128.523 $w=3.3e-07 $l=7.35e-07 $layer=POLY_cond $X=9.945 $Y=1.16
+ $X2=9.21 $Y2=1.16
r152 18 56 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=9.135 $Y=1.325
+ $X2=9.105 $Y2=1.16
r153 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.135 $Y=1.325
+ $X2=9.135 $Y2=1.985
r154 15 56 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=9.135 $Y=0.995
+ $X2=9.105 $Y2=1.16
r155 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.135 $Y=0.995
+ $X2=9.135 $Y2=0.56
r156 11 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.775 $Y=1.575
+ $X2=7.775 $Y2=1.74
r157 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=7.775 $Y=1.575
+ $X2=7.775 $Y2=0.445
r158 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.905
+ $X2=7.66 $Y2=1.74
r159 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.66 $Y=1.905
+ $X2=7.66 $Y2=2.275
r160 2 47 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=8.38
+ $Y=1.485 $X2=8.505 $Y2=1.95
r161 1 43 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=8.38
+ $Y=0.235 $X2=8.505 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_1346_413# 1 2 7 9 12 14 15 16 20 27 30 33
+ 34
c88 30 0 1.02967e-19 $X=8.23 $Y=1.16
c89 27 0 4.21632e-20 $X=7.5 $Y=2.165
c90 15 0 1.25869e-19 $X=8.715 $Y=1.16
c91 12 0 9.95676e-20 $X=8.715 $Y=1.985
r92 33 35 11.5578 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=7.435 $Y=1.16
+ $X2=7.435 $Y2=1.405
r93 33 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=1.16
+ $X2=7.435 $Y2=0.995
r94 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.16 $X2=8.23 $Y2=1.16
r95 28 33 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.585 $Y=1.16
+ $X2=7.435 $Y2=1.16
r96 28 30 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=7.585 $Y=1.16
+ $X2=8.23 $Y2=1.16
r97 27 35 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.5 $Y=2.165 $X2=7.5
+ $Y2=1.405
r98 24 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.37 $Y=0.535
+ $X2=7.37 $Y2=0.995
r99 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.285 $Y=0.45
+ $X2=7.37 $Y2=0.535
r100 20 22 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.285 $Y=0.45
+ $X2=7.08 $Y2=0.45
r101 16 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.415 $Y=2.25
+ $X2=7.5 $Y2=2.165
r102 16 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.415 $Y=2.25
+ $X2=6.865 $Y2=2.25
r103 14 31 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=8.64 $Y=1.16
+ $X2=8.23 $Y2=1.16
r104 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.64 $Y=1.16
+ $X2=8.715 $Y2=1.16
r105 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.715 $Y=1.325
+ $X2=8.715 $Y2=1.16
r106 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.715 $Y=1.325
+ $X2=8.715 $Y2=1.985
r107 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.715 $Y=0.995
+ $X2=8.715 $Y2=1.16
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.715 $Y=0.995
+ $X2=8.715 $Y2=0.56
r109 2 18 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=2.065 $X2=6.865 $Y2=2.25
r110 1 22 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=6.86
+ $Y=0.235 $X2=7.08 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_1948_47# 1 2 9 12 14 16 19 24 25 28 31 32
+ 34
r60 28 30 6.2579 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=9.825 $Y=0.51
+ $X2=9.825 $Y2=0.62
r61 25 35 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=10.487 $Y=1.16
+ $X2=10.487 $Y2=1.325
r62 25 34 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=10.487 $Y=1.16
+ $X2=10.487 $Y2=0.995
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.475
+ $Y=1.16 $X2=10.475 $Y2=1.16
r64 22 32 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=10.03 $Y=1.16
+ $X2=9.905 $Y2=1.16
r65 22 24 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=10.03 $Y=1.16
+ $X2=10.475 $Y2=1.16
r66 20 32 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=9.905 $Y=1.325
+ $X2=9.905 $Y2=1.16
r67 20 31 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=9.905 $Y=1.325
+ $X2=9.905 $Y2=1.685
r68 19 32 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=9.865 $Y=0.995
+ $X2=9.905 $Y2=1.16
r69 19 30 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.865 $Y=0.995
+ $X2=9.865 $Y2=0.62
r70 14 31 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.85
+ $X2=9.865 $Y2=1.685
r71 14 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=9.865 $Y=1.85
+ $X2=9.865 $Y2=2
r72 12 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.56 $Y=1.985
+ $X2=10.56 $Y2=1.325
r73 9 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.56 $Y=0.56
+ $X2=10.56 $Y2=0.995
r74 2 16 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=9.74
+ $Y=1.845 $X2=9.865 $Y2=2
r75 1 28 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=9.74
+ $Y=0.235 $X2=9.865 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 53
+ 54 56 57 59 60 61 63 68 92 96 103 104 107 110 113 116
c169 104 0 1.8506e-19 $X=10.81 $Y=2.72
c170 48 0 1.53472e-19 $X=10.35 $Y=1.66
c171 44 0 1.70577e-19 $X=8.925 $Y=1.79
c172 2 0 3.41142e-19 $X=1.905 $Y=1.845
c173 1 0 5.65522e-20 $X=0.545 $Y=1.815
r174 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r175 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r176 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r177 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r178 104 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r179 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r180 101 116 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=10.515 $Y=2.72
+ $X2=10.362 $Y2=2.72
r181 101 103 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.515 $Y=2.72
+ $X2=10.81 $Y2=2.72
r182 100 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r183 100 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=8.97 $Y2=2.72
r184 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r185 97 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=2.72
+ $X2=8.925 $Y2=2.72
r186 97 99 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.01 $Y=2.72
+ $X2=9.89 $Y2=2.72
r187 96 116 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=10.21 $Y=2.72
+ $X2=10.362 $Y2=2.72
r188 96 99 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.21 $Y=2.72
+ $X2=9.89 $Y2=2.72
r189 95 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r190 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r191 92 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.84 $Y=2.72
+ $X2=8.925 $Y2=2.72
r192 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.84 $Y=2.72
+ $X2=8.51 $Y2=2.72
r193 91 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r194 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r195 88 91 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r196 87 90 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=7.59 $Y2=2.72
r197 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r198 85 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r199 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r200 82 85 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r201 81 84 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.75 $Y2=2.72
r202 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r203 79 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r204 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r205 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 76 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r207 75 78 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r208 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r209 73 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.04 $Y2=2.72
r210 73 75 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.53 $Y2=2.72
r211 72 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r212 72 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r213 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r214 69 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r215 69 71 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r216 68 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=2.04 $Y2=2.72
r217 68 71 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=1.61 $Y2=2.72
r218 63 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r219 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r220 61 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r221 61 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r222 59 90 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.765 $Y=2.72
+ $X2=7.59 $Y2=2.72
r223 59 60 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=7.765 $Y=2.72
+ $X2=7.917 $Y2=2.72
r224 58 94 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.07 $Y=2.72
+ $X2=8.51 $Y2=2.72
r225 58 60 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.07 $Y=2.72
+ $X2=7.917 $Y2=2.72
r226 56 84 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=2.72
+ $X2=5.75 $Y2=2.72
r227 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=2.72
+ $X2=5.97 $Y2=2.72
r228 55 87 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=6.21 $Y2=2.72
r229 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.72
+ $X2=5.97 $Y2=2.72
r230 54 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.91 $Y2=2.72
r231 53 78 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=2.72
+ $X2=3.45 $Y2=2.72
r232 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=2.72
+ $X2=3.825 $Y2=2.72
r233 48 51 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=10.362 $Y=1.66
+ $X2=10.362 $Y2=2
r234 46 116 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=10.362 $Y=2.635
+ $X2=10.362 $Y2=2.72
r235 46 51 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=10.362 $Y=2.635
+ $X2=10.362 $Y2=2
r236 42 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.925 $Y=2.635
+ $X2=8.925 $Y2=2.72
r237 42 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.925 $Y=2.635
+ $X2=8.925 $Y2=1.79
r238 38 60 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.917 $Y=2.635
+ $X2=7.917 $Y2=2.72
r239 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=7.917 $Y=2.635
+ $X2=7.917 $Y2=2.3
r240 34 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=2.635
+ $X2=5.97 $Y2=2.72
r241 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.97 $Y=2.635
+ $X2=5.97 $Y2=2
r242 30 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=2.635
+ $X2=3.825 $Y2=2.72
r243 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.825 $Y=2.635
+ $X2=3.825 $Y2=2.33
r244 26 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r245 26 28 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.33
r246 22 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r247 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r248 7 51 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=10.15
+ $Y=1.845 $X2=10.35 $Y2=2
r249 7 48 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=10.15
+ $Y=1.845 $X2=10.35 $Y2=1.66
r250 6 44 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=8.79
+ $Y=1.485 $X2=8.925 $Y2=1.79
r251 5 40 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=2.065 $X2=7.98 $Y2=2.3
r252 4 36 300 $w=1.7e-07 $l=4.06202e-07 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=2.065 $X2=5.97 $Y2=2
r253 3 32 600 $w=1.7e-07 $l=5.59308e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.845 $X2=3.825 $Y2=2.33
r254 2 28 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2.33
r255 1 24 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%A_556_369# 1 2 3 4 13 17 22 24 25 26 27 28
+ 30 32 36 38 39
c113 17 0 1.20015e-19 $X=3.405 $Y=0.36
r114 39 41 18.6318 $w=2.39e-07 $l=3.65e-07 $layer=LI1_cond $X=4.307 $Y=1.91
+ $X2=4.307 $Y2=2.275
r115 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.25 $Y=0.45 $X2=4.35
+ $Y2=0.45
r116 32 39 5.37298 $w=2.39e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.25 $Y=1.825
+ $X2=4.307 $Y2=1.91
r117 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.885
+ $X2=4.25 $Y2=0.8
r118 31 32 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.25 $Y=0.885
+ $X2=4.25 $Y2=1.825
r119 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.715
+ $X2=4.25 $Y2=0.8
r120 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.25 $Y=0.535
+ $X2=4.25 $Y2=0.45
r121 29 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.25 $Y=0.535
+ $X2=4.25 $Y2=0.715
r122 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=0.8
+ $X2=4.25 $Y2=0.8
r123 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.165 $Y=0.8
+ $X2=3.575 $Y2=0.8
r124 25 39 2.73298 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.165 $Y=1.91
+ $X2=4.307 $Y2=1.91
r125 25 26 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.165 $Y=1.91
+ $X2=3.57 $Y2=1.91
r126 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.49 $Y=0.715
+ $X2=3.575 $Y2=0.8
r127 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.49 $Y=0.445
+ $X2=3.49 $Y2=0.715
r128 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.485 $Y=1.995
+ $X2=3.57 $Y2=1.91
r129 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.485 $Y=1.995
+ $X2=3.485 $Y2=2.245
r130 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.405 $Y=0.36
+ $X2=3.49 $Y2=0.445
r131 17 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.405 $Y=0.36
+ $X2=2.995 $Y2=0.36
r132 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.4 $Y=2.33
+ $X2=3.485 $Y2=2.245
r133 13 15 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.4 $Y=2.33
+ $X2=2.915 $Y2=2.33
r134 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=2.065 $X2=4.365 $Y2=2.275
r135 3 15 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.845 $X2=2.915 $Y2=2.33
r136 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.235 $X2=4.35 $Y2=0.45
r137 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.995 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%Q 1 2 9 12 13 14 17
c43 12 0 2.25437e-19 $X=9.5 $Y=1.43
r44 14 17 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=9.355 $Y=0.51
+ $X2=9.355 $Y2=0.395
r45 13 14 7.07929 $w=3.48e-07 $l=2.15e-07 $layer=LI1_cond $X=9.355 $Y=0.725
+ $X2=9.355 $Y2=0.51
r46 11 13 3.07305 $w=3.97e-07 $l=1.88481e-07 $layer=LI1_cond $X=9.5 $Y=0.825
+ $X2=9.355 $Y2=0.725
r47 11 12 31.6922 $w=2.18e-07 $l=6.05e-07 $layer=LI1_cond $X=9.5 $Y=0.825
+ $X2=9.5 $Y2=1.43
r48 7 12 4.41447 $w=3.04e-07 $l=1.81865e-07 $layer=LI1_cond $X=9.365 $Y=1.54
+ $X2=9.5 $Y2=1.43
r49 7 9 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.365 $Y=1.54
+ $X2=9.365 $Y2=1.67
r50 2 9 300 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=2 $X=9.21
+ $Y=1.485 $X2=9.345 $Y2=1.67
r51 1 17 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=9.21
+ $Y=0.235 $X2=9.345 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%Q_N 1 2 7 11 12 26
r15 16 26 1.89814 $w=2.53e-07 $l=4.2e-08 $layer=LI1_cond $X=10.812 $Y=1.572
+ $X2=10.812 $Y2=1.53
r16 12 26 0.994265 $w=2.53e-07 $l=2.2e-08 $layer=LI1_cond $X=10.812 $Y=1.508
+ $X2=10.812 $Y2=1.53
r17 12 19 10.259 $w=2.53e-07 $l=2.27e-07 $layer=LI1_cond $X=10.812 $Y=1.593
+ $X2=10.812 $Y2=1.82
r18 12 16 0.949071 $w=2.53e-07 $l=2.1e-08 $layer=LI1_cond $X=10.812 $Y=1.593
+ $X2=10.812 $Y2=1.572
r19 11 12 21.7855 $w=3.63e-07 $l=6.5e-07 $layer=LI1_cond $X=10.835 $Y=0.795
+ $X2=10.835 $Y2=1.445
r20 7 11 6.13261 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=10.812 $Y=0.668
+ $X2=10.812 $Y2=0.795
r21 7 9 1.81804 $w=2.55e-07 $l=3.8e-08 $layer=LI1_cond $X=10.812 $Y=0.668
+ $X2=10.812 $Y2=0.63
r22 2 19 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=10.635
+ $Y=1.485 $X2=10.77 $Y2=1.82
r23 1 9 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=10.635
+ $Y=0.235 $X2=10.77 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__SDFXBP_1%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 46 50
+ 53 54 55 57 62 67 82 86 93 94 97 100 103 106 109 112
c179 94 0 2.71124e-20 $X=10.81 $Y=0
c180 46 0 1.70577e-19 $X=8.925 $Y=0.53
r181 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r182 109 110 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r183 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r184 104 107 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.75 $Y2=0
r185 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r186 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r187 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r188 94 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=10.35 $Y2=0
r189 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r190 91 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.35 $Y2=0
r191 91 93 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.81 $Y2=0
r192 90 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r193 90 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=8.97 $Y2=0
r194 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r195 87 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0 $X2=8.925
+ $Y2=0
r196 87 89 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.01 $Y=0 $X2=9.89
+ $Y2=0
r197 86 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=10.35 $Y2=0
r198 86 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=9.89 $Y2=0
r199 85 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r200 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r201 82 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.84 $Y=0 $X2=8.925
+ $Y2=0
r202 82 84 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=8.51
+ $Y2=0
r203 81 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r204 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r205 78 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.59 $Y2=0
r206 78 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r207 77 80 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=7.59
+ $Y2=0
r208 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r209 75 106 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.045 $Y=0
+ $X2=5.86 $Y2=0
r210 75 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=0
+ $X2=6.21 $Y2=0
r211 74 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r212 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r213 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r214 71 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r215 70 73 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r216 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r217 68 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0
+ $X2=2.12 $Y2=0
r218 68 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.53
+ $Y2=0
r219 67 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.845
+ $Y2=0
r220 67 73 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.45
+ $Y2=0
r221 66 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r222 66 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r223 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r224 63 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r225 63 65 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r226 62 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0
+ $X2=2.12 $Y2=0
r227 62 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.61
+ $Y2=0
r228 57 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r229 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r230 55 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r231 55 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r232 53 80 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.7 $Y=0 $X2=7.59
+ $Y2=0
r233 53 54 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.7 $Y=0 $X2=7.885
+ $Y2=0
r234 52 84 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=8.51
+ $Y2=0
r235 52 54 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.07 $Y=0 $X2=7.885
+ $Y2=0
r236 48 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.35 $Y=0.085
+ $X2=10.35 $Y2=0
r237 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.35 $Y=0.085
+ $X2=10.35 $Y2=0.38
r238 44 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.925 $Y=0.085
+ $X2=8.925 $Y2=0
r239 44 46 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.925 $Y=0.085
+ $X2=8.925 $Y2=0.53
r240 40 54 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=0.085
+ $X2=7.885 $Y2=0
r241 40 42 11.3687 $w=3.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.885 $Y=0.085
+ $X2=7.885 $Y2=0.45
r242 36 106 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=0.085
+ $X2=5.86 $Y2=0
r243 36 38 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.86 $Y=0.085
+ $X2=5.86 $Y2=0.42
r244 35 103 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.845
+ $Y2=0
r245 34 106 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.675 $Y=0
+ $X2=5.86 $Y2=0
r246 34 35 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=5.675 $Y=0
+ $X2=3.945 $Y2=0
r247 30 103 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0
r248 30 32 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.845 $Y=0.085
+ $X2=3.845 $Y2=0.38
r249 26 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0
r250 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.36
r251 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r252 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r253 7 50 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=10.15
+ $Y=0.235 $X2=10.35 $Y2=0.38
r254 6 46 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=8.79
+ $Y=0.235 $X2=8.925 $Y2=0.53
r255 5 42 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=7.85
+ $Y=0.235 $X2=7.985 $Y2=0.45
r256 4 38 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.93 $Y2=0.42
r257 3 32 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.235 $X2=3.83 $Y2=0.38
r258 2 28 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.12 $Y2=0.36
r259 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


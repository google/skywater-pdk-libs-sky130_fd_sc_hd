* File: sky130_fd_sc_hd__a2bb2oi_2.spice
* Created: Thu Aug 27 14:03:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2bb2oi_2.pex.spice"
.subckt sky130_fd_sc_hd__a2bb2oi_2  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1002 N_A_136_47#_M1002_d N_B1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1011_d N_B2_M1011_g N_A_136_47#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1016 N_Y_M1011_d N_B2_M1016_g N_A_136_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_136_47#_M1016_s N_B1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_A_442_21#_M1001_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1001_d N_A_442_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1006_s N_A1_N_M1014_g N_A_442_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A1_N_M1017_g N_A_442_21#_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75003.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_A_442_21#_M1012_d N_A2_N_M1012_g N_VGND_M1017_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_A_442_21#_M1012_d N_A2_N_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75004.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_54_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1004_d N_B2_M1007_g N_A_54_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_B2_M1008_g N_A_54_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1008_d N_B1_M1005_g N_A_54_297#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_442_21#_M1000_g N_A_54_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1000_d N_A_442_21#_M1015_g N_A_54_297#_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_N_M1009_g N_A_662_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1009_d N_A1_N_M1019_g N_A_662_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1010 N_A_662_297#_M1019_s N_A2_N_M1010_g N_A_442_21#_M1010_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1013 N_A_662_297#_M1013_d N_A2_N_M1013_g N_A_442_21#_M1010_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__a2bb2oi_2.pxi.spice"
*
.ends
*
*

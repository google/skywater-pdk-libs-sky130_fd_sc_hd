* File: sky130_fd_sc_hd__o32a_4.spice
* Created: Thu Aug 27 14:41:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o32a_4.pex.spice"
.subckt sky130_fd_sc_hd__o32a_4  VNB VPB A1 A2 A3 B1 B2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B2	B2
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1012 N_A_27_47#_M1012_d N_A1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1027 N_A_27_47#_M1027_d N_A1_M1027_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1016 N_A_27_47#_M1027_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1018 N_A_27_47#_M1018_d N_A2_M1018_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1018_d N_A3_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.08775 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_27_47#_M1017_d N_A3_M1017_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_549_297#_M1001_d N_B1_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1023 N_A_549_297#_M1023_d N_B1_M1023_g N_A_27_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_A_549_297#_M1023_d N_B2_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.0975 PD=0.92 PS=0.95 NRD=0 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_549_297#_M1006_d N_B2_M1006_g N_A_27_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.0975 PD=1.82 PS=0.95 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_A_549_297#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1000_d N_A_549_297#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1024 N_X_M1024_d N_A_549_297#_M1024_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1025 N_X_M1024_d N_A_549_297#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_297#_M1007_d N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1019 N_A_27_297#_M1019_d N_A1_M1019_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1003 N_A_277_297#_M1003_d N_A2_M1003_g N_A_27_297#_M1019_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1026 N_A_277_297#_M1003_d N_A2_M1026_g N_A_27_297#_M1026_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_277_297#_M1009_d N_A3_M1009_g N_A_549_297#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_A_277_297#_M1015_d N_A3_M1015_g N_A_549_297#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1011 N_A_739_297#_M1011_d N_B1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1013 N_A_739_297#_M1013_d N_B1_M1013_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1008 N_A_549_297#_M1008_d N_B2_M1008_g N_A_739_297#_M1013_d VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_549_297#_M1008_d N_B2_M1010_g N_A_739_297#_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.15 AS=0.26 PD=1.3 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_549_297#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1002_d N_A_549_297#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1020 N_X_M1020_d N_A_549_297#_M1020_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1022 N_X_M1020_d N_A_549_297#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX28_noxref VNB VPB NWDIODE A=13.8993 P=20.53
c_77 VNB 0 1.81415e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__o32a_4.pxi.spice"
*
.ends
*
*

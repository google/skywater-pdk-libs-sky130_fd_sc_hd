* File: sky130_fd_sc_hd__or2_4.pxi.spice
* Created: Thu Aug 27 14:42:48 2020
* 
x_PM_SKY130_FD_SC_HD__OR2_4%B N_B_c_58_n N_B_M1011_g N_B_M1006_g B B N_B_c_60_n
+ PM_SKY130_FD_SC_HD__OR2_4%B
x_PM_SKY130_FD_SC_HD__OR2_4%A N_A_M1009_g N_A_M1002_g A N_A_c_89_n N_A_c_90_n
+ PM_SKY130_FD_SC_HD__OR2_4%A
x_PM_SKY130_FD_SC_HD__OR2_4%A_35_297# N_A_35_297#_M1011_d N_A_35_297#_M1006_s
+ N_A_35_297#_c_122_n N_A_35_297#_M1001_g N_A_35_297#_M1000_g
+ N_A_35_297#_c_123_n N_A_35_297#_M1004_g N_A_35_297#_M1003_g
+ N_A_35_297#_c_124_n N_A_35_297#_M1005_g N_A_35_297#_M1007_g
+ N_A_35_297#_c_125_n N_A_35_297#_M1008_g N_A_35_297#_M1010_g
+ N_A_35_297#_c_132_n N_A_35_297#_c_138_n N_A_35_297#_c_126_n
+ N_A_35_297#_c_153_n N_A_35_297#_c_156_n N_A_35_297#_c_134_n
+ N_A_35_297#_c_188_p N_A_35_297#_c_135_n N_A_35_297#_c_145_n
+ N_A_35_297#_c_127_n PM_SKY130_FD_SC_HD__OR2_4%A_35_297#
x_PM_SKY130_FD_SC_HD__OR2_4%VPWR N_VPWR_M1002_d N_VPWR_M1003_s N_VPWR_M1010_s
+ N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n
+ N_VPWR_c_258_n N_VPWR_c_259_n VPWR N_VPWR_c_260_n N_VPWR_c_261_n
+ N_VPWR_c_252_n PM_SKY130_FD_SC_HD__OR2_4%VPWR
x_PM_SKY130_FD_SC_HD__OR2_4%X N_X_M1001_d N_X_M1005_d N_X_M1000_d N_X_M1007_d
+ N_X_c_310_n N_X_c_301_n N_X_c_302_n N_X_c_322_n N_X_c_326_n N_X_c_329_n
+ N_X_c_335_n N_X_c_338_n N_X_c_303_n N_X_c_343_n N_X_c_345_n N_X_c_304_n
+ N_X_c_355_n X N_X_c_307_n PM_SKY130_FD_SC_HD__OR2_4%X
x_PM_SKY130_FD_SC_HD__OR2_4%VGND N_VGND_M1011_s N_VGND_M1009_d N_VGND_M1004_s
+ N_VGND_M1008_s N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n
+ N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n
+ VGND N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n
+ PM_SKY130_FD_SC_HD__OR2_4%VGND
cc_1 VNB N_B_c_58_n 0.0187567f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB B 0.0206831f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_B_c_60_n 0.0383638f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_4 VNB A 0.00389478f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_A_c_89_n 0.0229788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_c_90_n 0.0172147f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_7 VNB N_A_35_297#_c_122_n 0.0168999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_35_297#_c_123_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_9 VNB N_A_35_297#_c_124_n 0.0157966f $X=-0.19 $Y=-0.24 $X2=0.217 $Y2=1.16
cc_10 VNB N_A_35_297#_c_125_n 0.0191474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_35_297#_c_126_n 0.00285945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_35_297#_c_127_n 0.0659673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_252_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_X_c_301_n 0.00217862f $X=-0.19 $Y=-0.24 $X2=0.217 $Y2=0.85
cc_15 VNB N_X_c_302_n 0.00222241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_X_c_303_n 0.0108848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_304_n 0.00222466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0224311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_391_n 0.0100926f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_20 VNB N_VGND_c_392_n 0.0185095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_393_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.217 $Y2=0.85
cc_22 VNB N_VGND_c_394_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_395_n 0.00419326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_396_n 0.0198074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_397_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_398_n 0.0188761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_399_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_400_n 0.0169753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_401_n 0.0133346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_402_n 0.181386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_B_M1006_g 0.0245932f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.985
cc_32 VPB B 0.00503328f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_33 VPB N_B_c_60_n 0.0108454f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_34 VPB N_A_M1002_g 0.0193101f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.985
cc_35 VPB A 0.00155218f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_36 VPB N_A_c_89_n 0.00401838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_35_297#_M1000_g 0.0190563f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_38 VPB N_A_35_297#_M1003_g 0.0184657f $X=-0.19 $Y=1.305 $X2=0.217 $Y2=0.85
cc_39 VPB N_A_35_297#_M1007_g 0.018496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_35_297#_M1010_g 0.021884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_35_297#_c_132_n 0.0307964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_35_297#_c_126_n 0.00162205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_35_297#_c_134_n 0.00152908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_35_297#_c_135_n 0.00716461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_35_297#_c_127_n 0.0114336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_253_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_47 VPB N_VPWR_c_254_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_48 VPB N_VPWR_c_255_n 0.00419326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_256_n 0.0323675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_257_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_258_n 0.0185656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_259_n 0.00323604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_260_n 0.017296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_261_n 0.0139971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_252_n 0.0507576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB X 0.010445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_X_c_307_n 0.0127598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 N_B_M1006_g N_A_M1002_g 0.0489446f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_59 N_B_c_60_n A 3.14407e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B_c_60_n N_A_c_89_n 0.0489446f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_61 N_B_c_58_n N_A_c_90_n 0.0114141f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_62 N_B_M1006_g N_A_35_297#_c_132_n 0.016289f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_63 N_B_c_58_n N_A_35_297#_c_138_n 0.0064372f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_64 N_B_c_58_n N_A_35_297#_c_126_n 0.00263079f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_65 N_B_M1006_g N_A_35_297#_c_126_n 0.00838774f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_66 N_B_c_60_n N_A_35_297#_c_126_n 0.0100446f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_M1006_g N_A_35_297#_c_135_n 0.0115914f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_68 B N_A_35_297#_c_135_n 0.0163216f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_69 N_B_c_60_n N_A_35_297#_c_135_n 0.00528653f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_70 N_B_c_58_n N_A_35_297#_c_145_n 0.00525302f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_71 B N_A_35_297#_c_145_n 0.0355419f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_72 N_B_M1006_g N_VPWR_c_256_n 0.00495816f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_73 N_B_M1006_g N_VPWR_c_252_n 0.00946309f $X=0.53 $Y=1.985 $X2=0 $Y2=0
cc_74 B N_VGND_M1011_s 0.00274532f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_75 B N_VGND_c_391_n 2.18612e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_76 N_B_c_58_n N_VGND_c_392_n 0.00448362f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_77 B N_VGND_c_392_n 0.0200799f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B_c_60_n N_VGND_c_392_n 0.00101431f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B_c_58_n N_VGND_c_396_n 0.00542757f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_c_58_n N_VGND_c_402_n 0.0104852f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_81 B N_VGND_c_402_n 0.0013663f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_A_35_297#_c_122_n 0.0158653f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_A_35_297#_M1000_g 0.0220703f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_A_35_297#_c_132_n 0.00285278f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_c_90_n N_A_35_297#_c_138_n 0.00457432f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_86 A N_A_35_297#_c_126_n 0.0251226f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_c_90_n N_A_35_297#_c_126_n 0.00905168f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_A_35_297#_c_153_n 0.0159973f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_89 A N_A_35_297#_c_153_n 0.0260143f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_A_35_297#_c_153_n 0.00256542f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_91 A N_A_35_297#_c_156_n 0.0144732f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_A_35_297#_c_134_n 8.50012e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 A N_A_35_297#_c_134_n 0.00610147f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A_c_90_n N_A_35_297#_c_145_n 0.00271381f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_95 A N_A_35_297#_c_127_n 0.0042063f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_89_n N_A_35_297#_c_127_n 0.018698f $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_M1002_g N_VPWR_c_253_n 0.00730536f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_M1002_g N_VPWR_c_256_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_VPWR_c_252_n 0.0108133f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_c_90_n N_X_c_302_n 4.02691e-19 $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_101 A N_VGND_c_393_n 0.0144654f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_c_89_n N_VGND_c_393_n 5.59096e-19 $X=0.95 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_c_90_n N_VGND_c_393_n 0.00620502f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_90_n N_VGND_c_396_n 0.00542757f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_c_90_n N_VGND_c_402_n 0.00995006f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_35_297#_c_153_n A_121_297# 0.00360686f $X=1.41 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_35_297#_c_135_n A_121_297# 0.00144354f $X=0.32 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_35_297#_c_153_n N_VPWR_M1002_d 0.00762776f $X=1.41 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_35_297#_M1000_g N_VPWR_c_253_n 0.00490039f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_110 N_A_35_297#_c_132_n N_VPWR_c_253_n 0.0187663f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_111 N_A_35_297#_c_153_n N_VPWR_c_253_n 0.0136682f $X=1.41 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_35_297#_M1003_g N_VPWR_c_254_n 0.00268723f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_A_35_297#_M1007_g N_VPWR_c_254_n 0.00146448f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_35_297#_M1010_g N_VPWR_c_255_n 0.00316354f $X=2.655 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_35_297#_c_132_n N_VPWR_c_256_n 0.0230561f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_116 N_A_35_297#_M1000_g N_VPWR_c_258_n 0.00541359f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_117 N_A_35_297#_M1003_g N_VPWR_c_258_n 0.00422241f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_35_297#_M1007_g N_VPWR_c_260_n 0.00422241f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_35_297#_M1010_g N_VPWR_c_260_n 0.00541359f $X=2.655 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_35_297#_M1006_s N_VPWR_c_252_n 0.00225715f $X=0.175 $Y=1.485 $X2=0
+ $Y2=0
cc_121 N_A_35_297#_M1000_g N_VPWR_c_252_n 0.00982391f $X=1.395 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_35_297#_M1003_g N_VPWR_c_252_n 0.00569656f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_35_297#_M1007_g N_VPWR_c_252_n 0.00569656f $X=2.235 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_35_297#_M1010_g N_VPWR_c_252_n 0.0105352f $X=2.655 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_35_297#_c_132_n N_VPWR_c_252_n 0.0134449f $X=0.32 $Y=2.3 $X2=0 $Y2=0
cc_126 N_A_35_297#_c_153_n N_X_M1000_d 0.00354302f $X=1.41 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_35_297#_c_122_n N_X_c_310_n 0.00565046f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_35_297#_c_123_n N_X_c_310_n 0.00632248f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_35_297#_c_124_n N_X_c_310_n 5.22228e-19 $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_35_297#_c_123_n N_X_c_301_n 0.00850187f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_35_297#_c_124_n N_X_c_301_n 0.00850187f $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_35_297#_c_188_p N_X_c_301_n 0.0355133f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_35_297#_c_127_n N_X_c_301_n 0.00221825f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_35_297#_c_122_n N_X_c_302_n 0.00338648f $X=1.395 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_35_297#_c_123_n N_X_c_302_n 0.00110527f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_35_297#_c_156_n N_X_c_302_n 0.015237f $X=1.512 $Y=1.245 $X2=0 $Y2=0
cc_137 N_A_35_297#_c_188_p N_X_c_302_n 0.012274f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_35_297#_c_127_n N_X_c_302_n 0.00230123f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_35_297#_M1003_g N_X_c_322_n 0.0100318f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_35_297#_M1007_g N_X_c_322_n 0.0100318f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_35_297#_c_188_p N_X_c_322_n 0.0113082f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_35_297#_c_127_n N_X_c_322_n 0.00159731f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_35_297#_c_123_n N_X_c_326_n 5.22228e-19 $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_35_297#_c_124_n N_X_c_326_n 0.00632248f $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_35_297#_c_125_n N_X_c_326_n 0.0109442f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_35_297#_M1003_g N_X_c_329_n 5.29007e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_35_297#_M1007_g N_X_c_329_n 0.00388148f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_35_297#_M1010_g N_X_c_329_n 9.81519e-19 $X=2.655 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_35_297#_c_153_n N_X_c_329_n 0.00498257f $X=1.41 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_35_297#_c_188_p N_X_c_329_n 0.0152981f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_35_297#_c_127_n N_X_c_329_n 0.00221277f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_35_297#_M1003_g N_X_c_335_n 8.34775e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_35_297#_M1007_g N_X_c_335_n 0.00310792f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_35_297#_M1010_g N_X_c_335_n 0.00734931f $X=2.655 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_35_297#_M1003_g N_X_c_338_n 5.19281e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_35_297#_M1007_g N_X_c_338_n 0.00620543f $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_35_297#_M1010_g N_X_c_338_n 0.00528656f $X=2.655 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_35_297#_c_125_n N_X_c_303_n 0.0115817f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_35_297#_c_188_p N_X_c_303_n 6.43913e-19 $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_35_297#_M1010_g N_X_c_343_n 0.0138268f $X=2.655 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_35_297#_c_188_p N_X_c_343_n 4.73169e-19 $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_35_297#_M1000_g N_X_c_345_n 0.00789006f $X=1.395 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_35_297#_M1003_g N_X_c_345_n 0.00747389f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_35_297#_M1007_g N_X_c_345_n 5.19281e-19 $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_35_297#_c_153_n N_X_c_345_n 0.0102191f $X=1.41 $Y=1.58 $X2=0 $Y2=0
cc_166 N_A_35_297#_c_188_p N_X_c_345_n 0.00348915f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_35_297#_c_127_n N_X_c_345_n 8.87525e-19 $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_35_297#_c_124_n N_X_c_304_n 0.00110527f $X=2.235 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_35_297#_c_125_n N_X_c_304_n 0.00110527f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_35_297#_c_188_p N_X_c_304_n 0.0262212f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_35_297#_c_127_n N_X_c_304_n 0.00230227f $X=2.655 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_35_297#_M1007_g N_X_c_355_n 4.64231e-19 $X=2.235 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_35_297#_M1010_g N_X_c_355_n 0.00187637f $X=2.655 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_35_297#_c_125_n X 0.024109f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_35_297#_c_188_p X 0.0141433f $X=2.255 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_35_297#_c_122_n N_VGND_c_393_n 0.00583105f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_35_297#_c_138_n N_VGND_c_393_n 0.0329353f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_178 N_A_35_297#_c_123_n N_VGND_c_394_n 0.00268723f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_35_297#_c_124_n N_VGND_c_394_n 0.00146448f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_35_297#_c_125_n N_VGND_c_395_n 0.00316354f $X=2.655 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_35_297#_c_138_n N_VGND_c_396_n 0.0153821f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_182 N_A_35_297#_c_122_n N_VGND_c_398_n 0.00541763f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_35_297#_c_123_n N_VGND_c_398_n 0.0042482f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_35_297#_c_124_n N_VGND_c_400_n 0.0042482f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_35_297#_c_125_n N_VGND_c_400_n 0.0042482f $X=2.655 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_35_297#_M1011_d N_VGND_c_402_n 0.00217091f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_187 N_A_35_297#_c_122_n N_VGND_c_402_n 0.00990849f $X=1.395 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_35_297#_c_123_n N_VGND_c_402_n 0.00573646f $X=1.815 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_35_297#_c_124_n N_VGND_c_402_n 0.00573646f $X=2.235 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_35_297#_c_125_n N_VGND_c_402_n 0.00677017f $X=2.655 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_35_297#_c_138_n N_VGND_c_402_n 0.0119633f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_192 A_121_297# N_VPWR_c_252_n 0.00897657f $X=0.605 $Y=1.485 $X2=0.605
+ $Y2=1.495
cc_193 N_VPWR_c_252_n N_X_M1000_d 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_252_n N_X_M1007_d 0.00215201f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_M1003_s N_X_c_322_n 0.00440038f $X=1.89 $Y=1.485 $X2=0 $Y2=0
cc_196 N_VPWR_c_254_n N_X_c_322_n 0.012179f $X=2.025 $Y=2.34 $X2=0 $Y2=0
cc_197 N_VPWR_c_258_n N_X_c_322_n 0.0020257f $X=1.94 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_260_n N_X_c_322_n 0.0020257f $X=2.78 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_252_n N_X_c_322_n 0.00841425f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_260_n N_X_c_338_n 0.0189039f $X=2.78 $Y=2.72 $X2=0 $Y2=0
cc_201 N_VPWR_c_252_n N_X_c_338_n 0.0122217f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_253_n N_X_c_345_n 0.0401692f $X=1.145 $Y=2.01 $X2=0 $Y2=0
cc_203 N_VPWR_c_258_n N_X_c_345_n 0.0188215f $X=1.94 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_c_252_n N_X_c_345_n 0.0121968f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_M1010_s N_X_c_307_n 0.00544116f $X=2.73 $Y=1.485 $X2=0 $Y2=0
cc_206 N_VPWR_c_255_n N_X_c_307_n 0.0142906f $X=2.865 $Y=2 $X2=0 $Y2=0
cc_207 N_X_c_301_n N_VGND_M1004_s 0.00162006f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_208 N_X_c_303_n N_VGND_M1008_s 0.00321757f $X=2.79 $Y=0.82 $X2=0 $Y2=0
cc_209 N_X_c_310_n N_VGND_c_393_n 0.0294569f $X=1.605 $Y=0.4 $X2=0 $Y2=0
cc_210 N_X_c_302_n N_VGND_c_393_n 0.00600337f $X=1.77 $Y=0.82 $X2=0 $Y2=0
cc_211 N_X_c_301_n N_VGND_c_394_n 0.0122414f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_212 N_X_c_303_n N_VGND_c_395_n 0.0134722f $X=2.79 $Y=0.82 $X2=0 $Y2=0
cc_213 N_X_c_310_n N_VGND_c_398_n 0.017716f $X=1.605 $Y=0.4 $X2=0 $Y2=0
cc_214 N_X_c_301_n N_VGND_c_398_n 0.00193763f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_215 N_X_c_301_n N_VGND_c_400_n 0.00193763f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_216 N_X_c_326_n N_VGND_c_400_n 0.017716f $X=2.445 $Y=0.4 $X2=0 $Y2=0
cc_217 N_X_c_303_n N_VGND_c_400_n 0.00194519f $X=2.79 $Y=0.82 $X2=0 $Y2=0
cc_218 N_X_c_303_n N_VGND_c_401_n 0.00306906f $X=2.79 $Y=0.82 $X2=0 $Y2=0
cc_219 N_X_M1001_d N_VGND_c_402_n 0.00215535f $X=1.47 $Y=0.235 $X2=0 $Y2=0
cc_220 N_X_M1005_d N_VGND_c_402_n 0.00215535f $X=2.31 $Y=0.235 $X2=0 $Y2=0
cc_221 N_X_c_310_n N_VGND_c_402_n 0.0121406f $X=1.605 $Y=0.4 $X2=0 $Y2=0
cc_222 N_X_c_301_n N_VGND_c_402_n 0.00825759f $X=2.28 $Y=0.82 $X2=0 $Y2=0
cc_223 N_X_c_326_n N_VGND_c_402_n 0.0121406f $X=2.445 $Y=0.4 $X2=0 $Y2=0
cc_224 N_X_c_303_n N_VGND_c_402_n 0.0097057f $X=2.79 $Y=0.82 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__edfxtp_1.spice.SKY130_FD_SC_HD__EDFXTP_1.pxi
* Created: Thu Aug 27 14:19:54 2020
* 
x_PM_SKY130_FD_SC_HD__EDFXTP_1%CLK N_CLK_c_220_n N_CLK_c_224_n N_CLK_c_221_n
+ N_CLK_M1031_g N_CLK_c_225_n N_CLK_M1015_g N_CLK_c_226_n CLK
+ PM_SKY130_FD_SC_HD__EDFXTP_1%CLK
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_27_47# N_A_27_47#_M1031_s N_A_27_47#_M1015_s
+ N_A_27_47#_M1017_g N_A_27_47#_M1000_g N_A_27_47#_M1006_g N_A_27_47#_M1010_g
+ N_A_27_47#_M1030_g N_A_27_47#_c_262_n N_A_27_47#_M1007_g N_A_27_47#_c_498_p
+ N_A_27_47#_c_264_n N_A_27_47#_c_265_n N_A_27_47#_c_277_n N_A_27_47#_c_398_p
+ N_A_27_47#_c_266_n N_A_27_47#_c_267_n N_A_27_47#_c_268_n N_A_27_47#_c_269_n
+ N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n N_A_27_47#_c_283_n
+ N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_c_286_n N_A_27_47#_c_270_n
+ N_A_27_47#_c_288_n N_A_27_47#_c_271_n N_A_27_47#_c_272_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%D N_D_M1002_g N_D_M1021_g N_D_c_512_n N_D_c_516_n
+ D N_D_c_514_n PM_SKY130_FD_SC_HD__EDFXTP_1%D
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_423_343# N_A_423_343#_M1029_s
+ N_A_423_343#_M1013_s N_A_423_343#_c_568_n N_A_423_343#_M1025_g
+ N_A_423_343#_M1018_g N_A_423_343#_c_569_n N_A_423_343#_c_563_n
+ N_A_423_343#_c_564_n N_A_423_343#_c_565_n N_A_423_343#_c_566_n
+ N_A_423_343#_c_567_n PM_SKY130_FD_SC_HD__EDFXTP_1%A_423_343#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%DE N_DE_M1004_g N_DE_c_651_n N_DE_c_652_n
+ N_DE_M1029_g N_DE_c_654_n N_DE_M1013_g N_DE_c_659_n N_DE_M1016_g N_DE_c_655_n
+ N_DE_c_661_n DE PM_SKY130_FD_SC_HD__EDFXTP_1%DE
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_791_264# N_A_791_264#_M1012_s
+ N_A_791_264#_M1027_s N_A_791_264#_M1032_g N_A_791_264#_M1026_g
+ N_A_791_264#_M1019_g N_A_791_264#_M1020_g N_A_791_264#_c_748_n
+ N_A_791_264#_c_749_n N_A_791_264#_c_750_n N_A_791_264#_c_737_n
+ N_A_791_264#_c_751_n N_A_791_264#_c_752_n N_A_791_264#_c_753_n
+ N_A_791_264#_c_738_n N_A_791_264#_c_739_n N_A_791_264#_c_740_n
+ N_A_791_264#_c_741_n N_A_791_264#_c_742_n N_A_791_264#_c_743_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%A_791_264#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_193_47# N_A_193_47#_M1017_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1009_g N_A_193_47#_c_902_n N_A_193_47#_M1028_g
+ N_A_193_47#_c_904_n N_A_193_47#_M1003_g N_A_193_47#_M1024_g
+ N_A_193_47#_c_905_n N_A_193_47#_c_906_n N_A_193_47#_c_914_n
+ N_A_193_47#_c_915_n N_A_193_47#_c_916_n N_A_193_47#_c_917_n
+ N_A_193_47#_c_960_n N_A_193_47#_c_907_n N_A_193_47#_c_908_n
+ N_A_193_47#_c_909_n N_A_193_47#_c_921_n N_A_193_47#_c_910_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_1150_159# N_A_1150_159#_M1022_d
+ N_A_1150_159#_M1014_d N_A_1150_159#_M1001_g N_A_1150_159#_M1033_g
+ N_A_1150_159#_M1023_g N_A_1150_159#_M1011_g N_A_1150_159#_c_1101_n
+ N_A_1150_159#_c_1102_n N_A_1150_159#_c_1103_n N_A_1150_159#_c_1104_n
+ N_A_1150_159#_c_1113_n N_A_1150_159#_c_1105_n N_A_1150_159#_c_1106_n
+ N_A_1150_159#_c_1107_n N_A_1150_159#_c_1108_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%A_1150_159#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_986_413# N_A_986_413#_M1006_d
+ N_A_986_413#_M1009_d N_A_986_413#_c_1216_n N_A_986_413#_M1014_g
+ N_A_986_413#_M1022_g N_A_986_413#_c_1217_n N_A_986_413#_c_1218_n
+ N_A_986_413#_c_1219_n N_A_986_413#_c_1220_n N_A_986_413#_c_1230_n
+ N_A_986_413#_c_1236_n N_A_986_413#_c_1221_n N_A_986_413#_c_1226_n
+ N_A_986_413#_c_1222_n PM_SKY130_FD_SC_HD__EDFXTP_1%A_986_413#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_1591_413# N_A_1591_413#_M1003_d
+ N_A_1591_413#_M1030_d N_A_1591_413#_M1012_g N_A_1591_413#_M1027_g
+ N_A_1591_413#_c_1323_n N_A_1591_413#_c_1324_n N_A_1591_413#_M1008_g
+ N_A_1591_413#_M1005_g N_A_1591_413#_c_1325_n N_A_1591_413#_c_1326_n
+ N_A_1591_413#_c_1327_n N_A_1591_413#_c_1339_n N_A_1591_413#_c_1342_n
+ N_A_1591_413#_c_1328_n N_A_1591_413#_c_1337_n N_A_1591_413#_c_1329_n
+ N_A_1591_413#_c_1330_n PM_SKY130_FD_SC_HD__EDFXTP_1%A_1591_413#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%VPWR N_VPWR_M1015_d N_VPWR_M1025_d N_VPWR_M1013_d
+ N_VPWR_M1001_d N_VPWR_M1023_s N_VPWR_M1019_d N_VPWR_M1027_d N_VPWR_c_1433_n
+ N_VPWR_c_1434_n N_VPWR_c_1435_n N_VPWR_c_1436_n N_VPWR_c_1437_n
+ N_VPWR_c_1438_n N_VPWR_c_1439_n N_VPWR_c_1440_n N_VPWR_c_1441_n
+ N_VPWR_c_1442_n N_VPWR_c_1443_n N_VPWR_c_1444_n N_VPWR_c_1445_n
+ N_VPWR_c_1446_n VPWR N_VPWR_c_1447_n N_VPWR_c_1448_n N_VPWR_c_1449_n
+ N_VPWR_c_1450_n N_VPWR_c_1432_n N_VPWR_c_1452_n N_VPWR_c_1453_n
+ N_VPWR_c_1454_n N_VPWR_c_1455_n PM_SKY130_FD_SC_HD__EDFXTP_1%VPWR
x_PM_SKY130_FD_SC_HD__EDFXTP_1%A_299_47# N_A_299_47#_M1002_s N_A_299_47#_M1032_d
+ N_A_299_47#_M1021_s N_A_299_47#_M1026_d N_A_299_47#_c_1596_n
+ N_A_299_47#_c_1588_n N_A_299_47#_c_1598_n N_A_299_47#_c_1589_n
+ N_A_299_47#_c_1590_n N_A_299_47#_c_1591_n N_A_299_47#_c_1592_n
+ N_A_299_47#_c_1593_n N_A_299_47#_c_1594_n N_A_299_47#_c_1595_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%A_299_47#
x_PM_SKY130_FD_SC_HD__EDFXTP_1%Q N_Q_M1008_d N_Q_M1005_d Q N_Q_c_1718_n
+ PM_SKY130_FD_SC_HD__EDFXTP_1%Q
x_PM_SKY130_FD_SC_HD__EDFXTP_1%VGND N_VGND_M1031_d N_VGND_M1004_d N_VGND_M1029_d
+ N_VGND_M1033_d N_VGND_M1011_s N_VGND_M1020_d N_VGND_M1012_d N_VGND_c_1735_n
+ N_VGND_c_1736_n N_VGND_c_1737_n N_VGND_c_1738_n N_VGND_c_1739_n
+ N_VGND_c_1740_n N_VGND_c_1741_n N_VGND_c_1742_n N_VGND_c_1743_n
+ N_VGND_c_1744_n N_VGND_c_1745_n N_VGND_c_1746_n N_VGND_c_1747_n
+ N_VGND_c_1748_n N_VGND_c_1749_n VGND N_VGND_c_1750_n N_VGND_c_1751_n
+ N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n N_VGND_c_1755_n
+ N_VGND_c_1756_n N_VGND_c_1757_n PM_SKY130_FD_SC_HD__EDFXTP_1%VGND
cc_1 VNB N_CLK_c_220_n 0.0573151f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_221_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0185843f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1017_g 0.0373293f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1006_g 0.0222595f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_6 VNB N_A_27_47#_c_262_n 0.0139254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1007_g 0.0461694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_264_n 0.00191938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_265_n 0.00646065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_266_n 0.0024678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_267_n 0.0042825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_268_n 0.0298396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_269_n 0.00478196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_270_n 0.0236749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_271_n 0.00915868f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_272_n 0.00210612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1002_g 0.0308382f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_18 VNB N_D_c_512_n 0.0161793f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_19 VNB D 0.00399003f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_20 VNB N_D_c_514_n 0.0145063f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_21 VNB N_A_423_343#_M1018_g 0.0217809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_423_343#_c_563_n 0.00769004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_423_343#_c_564_n 0.00185686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_423_343#_c_565_n 0.00333068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_423_343#_c_566_n 0.0291606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_423_343#_c_567_n 0.00198824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_DE_M1004_g 0.0211774f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_28 VNB N_DE_c_651_n 0.0423212f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_29 VNB N_DE_c_652_n 0.032977f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_30 VNB N_DE_M1029_g 0.0242274f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_31 VNB N_DE_c_654_n 0.0180937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_DE_c_655_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB DE 0.0110099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_791_264#_M1032_g 0.0534418f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_35 VNB N_A_791_264#_M1020_g 0.0480681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_791_264#_c_737_n 0.00377528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_791_264#_c_738_n 0.00469958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_791_264#_c_739_n 0.0395002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_791_264#_c_740_n 0.00419717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_791_264#_c_741_n 0.0132319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_791_264#_c_742_n 0.0013422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_791_264#_c_743_n 0.00158979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_902_n 0.0136524f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_44 VNB N_A_193_47#_M1028_g 0.0429795f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_45 VNB N_A_193_47#_c_904_n 0.0180286f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_46 VNB N_A_193_47#_c_905_n 0.00392862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_906_n 0.0296727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_907_n 0.0032859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_193_47#_c_908_n 0.0119889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_c_909_n 0.00248621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_193_47#_c_910_n 0.0122334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1150_159#_M1001_g 0.0138674f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_53 VNB N_A_1150_159#_M1033_g 0.0197771f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_54 VNB N_A_1150_159#_M1011_g 0.0283997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1150_159#_c_1101_n 0.0223712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1150_159#_c_1102_n 0.00481399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1150_159#_c_1103_n 0.00932364f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1150_159#_c_1104_n 0.00611738f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1150_159#_c_1105_n 0.0048611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1150_159#_c_1106_n 0.0162827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1150_159#_c_1107_n 0.00249997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1150_159#_c_1108_n 0.0317753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_986_413#_c_1216_n 0.0113827f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_64 VNB N_A_986_413#_c_1217_n 0.0181892f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_65 VNB N_A_986_413#_c_1218_n 0.0133197f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_66 VNB N_A_986_413#_c_1219_n 0.00937183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_986_413#_c_1220_n 0.00117523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_986_413#_c_1221_n 0.0117046f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_986_413#_c_1222_n 0.00182328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1591_413#_M1012_g 0.0350674f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_71 VNB N_A_1591_413#_c_1323_n 0.0145702f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_72 VNB N_A_1591_413#_c_1324_n 0.0205457f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_73 VNB N_A_1591_413#_c_1325_n 0.0384709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1591_413#_c_1326_n 0.004935f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1591_413#_c_1327_n 0.0137821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1591_413#_c_1328_n 0.00719187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1591_413#_c_1329_n 0.00330077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1591_413#_c_1330_n 0.002763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VPWR_c_1432_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_299_47#_c_1588_n 0.0139151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_299_47#_c_1589_n 0.00311002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_299_47#_c_1590_n 0.00675947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_299_47#_c_1591_n 0.00419923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_299_47#_c_1592_n 4.93883e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_299_47#_c_1593_n 0.00440827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_299_47#_c_1594_n 0.00402556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_299_47#_c_1595_n 0.00400821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_Q_c_1718_n 0.0401252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1735_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1736_n 0.00461568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1737_n 4.14e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1738_n 0.00284902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1739_n 0.00256722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1740_n 0.00698438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1741_n 0.00947199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1742_n 0.0365941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1743_n 0.00507461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1744_n 0.0222458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1745_n 0.00408091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1746_n 0.042635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1747_n 0.0049096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1748_n 0.0189086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1749_n 0.00471252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1750_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1751_n 0.0165213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1752_n 0.0645626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1753_n 0.0230523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1754_n 0.525311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1755_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1756_n 0.00436942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1757_n 0.00597188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VPB N_CLK_c_220_n 0.0047794f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_113 VPB N_CLK_c_224_n 0.0162092f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_114 VPB N_CLK_c_225_n 0.01861f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_115 VPB N_CLK_c_226_n 0.0230979f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_116 VPB CLK 0.0175757f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_117 VPB N_A_27_47#_M1000_g 0.0377949f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_118 VPB N_A_27_47#_M1010_g 0.0194293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_M1030_g 0.033317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_262_n 0.0198419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_277_n 0.0018131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_266_n 0.00333071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_269_n 0.00290992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_280_n 0.00357396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_281_n 0.0245693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_282_n 0.00167507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_283_n 0.0139626f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_284_n 0.00136166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_285_n 0.00815911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_286_n 0.0048201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_270_n 0.0117983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_288_n 0.0276115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_271_n 0.0212228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_272_n 0.00662783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_D_M1021_g 0.0238916f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_136 VPB N_D_c_516_n 0.0159446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB D 0.00181411f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_138 VPB N_D_c_514_n 0.0165468f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_139 VPB N_A_423_343#_c_568_n 0.0753975f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_140 VPB N_A_423_343#_c_569_n 0.0076426f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_141 VPB N_A_423_343#_c_564_n 0.00615569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_DE_c_654_n 0.0104063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_DE_M1013_g 0.0255037f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_144 VPB N_DE_c_659_n 0.0220855f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_145 VPB N_DE_M1016_g 0.0236724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_DE_c_661_n 0.00456175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB DE 0.00246649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_791_264#_M1032_g 8.98279e-19 $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_149 VPB N_A_791_264#_M1026_g 0.0248815f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_150 VPB N_A_791_264#_M1019_g 0.0241837f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_151 VPB N_A_791_264#_M1020_g 0.0184691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_791_264#_c_748_n 0.011879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_791_264#_c_749_n 0.040689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_791_264#_c_750_n 0.00761748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_791_264#_c_751_n 0.00659101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_791_264#_c_752_n 0.0310969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_791_264#_c_753_n 0.00248001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_791_264#_c_741_n 6.77134e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_791_264#_c_743_n 0.00225466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_193_47#_M1009_g 0.0469787f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_161 VPB N_A_193_47#_c_902_n 0.0138415f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_162 VPB N_A_193_47#_M1024_g 0.0210318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_193_47#_c_914_n 0.0361515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_193_47#_c_915_n 0.00566519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_193_47#_c_916_n 0.0211513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_193_47#_c_917_n 0.0012313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_193_47#_c_907_n 0.00673154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_193_47#_c_908_n 0.0201772f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_193_47#_c_909_n 0.00152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_193_47#_c_921_n 0.0265183f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_193_47#_c_910_n 0.00945279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1150_159#_M1001_g 0.0519779f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_173 VPB N_A_1150_159#_M1023_g 0.0564064f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_174 VPB N_A_1150_159#_c_1102_n 0.00955004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1150_159#_c_1103_n 0.00154645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1150_159#_c_1113_n 0.0154933f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1150_159#_c_1105_n 0.00366659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_986_413#_M1014_g 0.0274355f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_179 VPB N_A_986_413#_c_1219_n 0.018904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_986_413#_c_1220_n 0.0102534f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_986_413#_c_1226_n 0.00394568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_986_413#_c_1222_n 0.00924579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1591_413#_M1027_g 0.0451789f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_184 VPB N_A_1591_413#_c_1323_n 0.00439136f $X=-0.19 $Y=1.305 $X2=0.33
+ $Y2=1.16
cc_185 VPB N_A_1591_413#_M1005_g 0.0237506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1591_413#_c_1325_n 0.0157863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1591_413#_c_1326_n 3.18387e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1591_413#_c_1327_n 8.89166e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1591_413#_c_1337_n 0.00704026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1591_413#_c_1329_n 0.00292829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1433_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1434_n 0.00843162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1435_n 0.00704186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1436_n 0.00505269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1437_n 0.0192928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1438_n 0.00629264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1439_n 0.00924361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1440_n 0.010598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1441_n 0.0365367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1442_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1443_n 0.0432692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1444_n 0.00497475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1445_n 0.0224066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1446_n 0.00468329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1447_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1448_n 0.0193581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1449_n 0.0730926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1450_n 0.0230248f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1432_n 0.0721263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1452_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1453_n 0.00372488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1454_n 0.00449095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1455_n 0.00442865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_299_47#_c_1596_n 0.00772563f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_A_299_47#_c_1588_n 0.00994696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_299_47#_c_1598_n 0.00581789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_299_47#_c_1589_n 0.00950245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_Q_c_1718_n 0.0436448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 N_CLK_c_220_n N_A_27_47#_M1017_g 0.00520193f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_220 N_CLK_c_221_n N_A_27_47#_M1017_g 0.0200589f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_221 CLK N_A_27_47#_M1017_g 3.12184e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_222 N_CLK_c_224_n N_A_27_47#_M1000_g 0.00541775f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_223 N_CLK_c_226_n N_A_27_47#_M1000_g 0.0276441f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_224 CLK N_A_27_47#_M1000_g 5.77812e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_225 N_CLK_c_220_n N_A_27_47#_c_264_n 0.00775742f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_226 N_CLK_c_221_n N_A_27_47#_c_264_n 0.00684762f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_227 CLK N_A_27_47#_c_264_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_228 N_CLK_c_220_n N_A_27_47#_c_265_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_229 CLK N_A_27_47#_c_265_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_230 N_CLK_c_225_n N_A_27_47#_c_277_n 0.0126874f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_231 N_CLK_c_226_n N_A_27_47#_c_277_n 0.00142281f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_232 CLK N_A_27_47#_c_277_n 0.00766156f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_233 N_CLK_c_220_n N_A_27_47#_c_266_n 0.0046428f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_234 N_CLK_c_224_n N_A_27_47#_c_266_n 7.07325e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_235 N_CLK_c_226_n N_A_27_47#_c_266_n 0.00436768f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_236 CLK N_A_27_47#_c_266_n 0.0511211f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_237 N_CLK_c_220_n N_A_27_47#_c_280_n 2.46885e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_238 N_CLK_c_225_n N_A_27_47#_c_280_n 2.17882e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_239 N_CLK_c_226_n N_A_27_47#_c_280_n 0.00343236f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_240 CLK N_A_27_47#_c_280_n 0.0153591f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_241 N_CLK_c_225_n N_A_27_47#_c_282_n 0.00101286f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_220_n N_A_27_47#_c_270_n 0.0169118f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_243 CLK N_A_27_47#_c_270_n 0.00161603f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_244 N_CLK_c_225_n N_VPWR_c_1433_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_245 N_CLK_c_225_n N_VPWR_c_1447_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_246 N_CLK_c_225_n N_VPWR_c_1432_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_247 N_CLK_c_221_n N_VGND_c_1735_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_248 N_CLK_c_220_n N_VGND_c_1750_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_249 N_CLK_c_221_n N_VGND_c_1750_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_250 N_CLK_c_221_n N_VGND_c_1754_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_281_n N_D_M1021_g 0.00440395f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1017_g N_D_c_512_n 0.00269191f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1000_g N_D_c_516_n 0.00269191f $X=0.89 $Y=2.135 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_281_n N_D_c_516_n 0.00153919f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_281_n D 0.00497736f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_270_n N_D_c_514_n 0.00269191f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_281_n N_A_423_343#_c_568_n 0.0120018f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_281_n N_A_423_343#_c_569_n 0.0221661f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_281_n N_A_423_343#_c_564_n 0.00660521f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_281_n N_DE_M1013_g 0.00347932f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_281_n N_DE_c_659_n 0.00132678f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_281_n N_DE_M1016_g 0.00575563f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_267_n N_A_791_264#_M1032_g 2.53945e-19 $X=5.15 $Y=0.845
+ $X2=0 $Y2=0
cc_264 N_A_27_47#_c_268_n N_A_791_264#_M1032_g 0.00303165f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_281_n N_A_791_264#_M1026_g 0.0043253f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1007_g N_A_791_264#_M1020_g 0.0443098f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_281_n N_A_791_264#_c_751_n 0.00923372f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_281_n N_A_791_264#_c_752_n 0.00184708f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1007_g N_A_791_264#_c_739_n 0.00644693f $X=8.51 $Y=0.415
+ $X2=0 $Y2=0
cc_270 N_A_27_47#_c_267_n N_A_791_264#_c_739_n 0.0294334f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_268_n N_A_791_264#_c_739_n 0.00161772f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_271_n N_A_791_264#_c_739_n 8.58822e-19 $X=7.875 $Y=1.32
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_272_n N_A_791_264#_c_739_n 0.00521916f $X=7.875 $Y=1.41
+ $X2=0 $Y2=0
cc_274 N_A_27_47#_c_281_n N_A_193_47#_M1000_d 0.00126326f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_269_n N_A_193_47#_M1009_g 7.3078e-19 $X=5.235 $Y=1.655 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_281_n N_A_193_47#_M1009_g 0.00666456f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_285_n N_A_193_47#_M1009_g 0.00270517f $X=5.295 $Y=1.87 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_288_n N_A_193_47#_M1009_g 0.0273982f $X=5.405 $Y=1.74 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_269_n N_A_193_47#_c_902_n 0.0120754f $X=5.235 $Y=1.655 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_285_n N_A_193_47#_c_902_n 0.00149465f $X=5.295 $Y=1.87 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_288_n N_A_193_47#_c_902_n 0.018371f $X=5.405 $Y=1.74 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_M1006_g N_A_193_47#_M1028_g 0.0124733f $X=4.99 $Y=0.415 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_267_n N_A_193_47#_M1028_g 0.00145899f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_268_n N_A_193_47#_M1028_g 0.0168195f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_269_n N_A_193_47#_M1028_g 0.00509325f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_286 N_A_27_47#_M1007_g N_A_193_47#_c_904_n 0.0144865f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_M1030_g N_A_193_47#_M1024_g 0.0175064f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1007_g N_A_193_47#_c_905_n 0.00658103f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_271_n N_A_193_47#_c_905_n 9.61914e-19 $X=7.875 $Y=1.32 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_M1007_g N_A_193_47#_c_906_n 0.0213226f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_271_n N_A_193_47#_c_906_n 0.0204217f $X=7.875 $Y=1.32 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_272_n N_A_193_47#_c_906_n 5.64291e-19 $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_281_n N_A_193_47#_c_914_n 0.279301f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1000_g N_A_193_47#_c_915_n 0.00457449f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_266_n N_A_193_47#_c_915_n 0.00673509f $X=0.76 $Y=1.235 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_281_n N_A_193_47#_c_915_n 0.0262177f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_262_n N_A_193_47#_c_916_n 0.00218822f $X=8.435 $Y=1.32 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_267_n N_A_193_47#_c_916_n 0.00220528f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_269_n N_A_193_47#_c_916_n 0.0122906f $X=5.235 $Y=1.655 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_281_n N_A_193_47#_c_916_n 0.00995021f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_283_n N_A_193_47#_c_916_n 0.185323f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_284_n N_A_193_47#_c_916_n 0.0254049f $X=5.44 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_285_n N_A_193_47#_c_916_n 0.00659382f $X=5.295 $Y=1.87 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_286_n N_A_193_47#_c_916_n 0.026031f $X=7.885 $Y=1.87 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_288_n N_A_193_47#_c_916_n 0.00183443f $X=5.405 $Y=1.74 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_271_n N_A_193_47#_c_916_n 0.00372733f $X=7.875 $Y=1.32 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_272_n N_A_193_47#_c_916_n 0.0147985f $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_267_n N_A_193_47#_c_917_n 0.00129557f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_269_n N_A_193_47#_c_917_n 0.00254764f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_281_n N_A_193_47#_c_917_n 0.0267692f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_272_n N_A_193_47#_c_960_n 6.47753e-19 $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_M1030_g N_A_193_47#_c_907_n 0.0020271f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_262_n N_A_193_47#_c_907_n 0.0169581f $X=8.435 $Y=1.32 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_M1007_g N_A_193_47#_c_907_n 0.00640774f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_286_n N_A_193_47#_c_907_n 0.00821717f $X=7.885 $Y=1.87 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_271_n N_A_193_47#_c_907_n 0.00345899f $X=7.875 $Y=1.32 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_272_n N_A_193_47#_c_907_n 0.051449f $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_267_n N_A_193_47#_c_908_n 0.00116173f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_268_n N_A_193_47#_c_908_n 0.0213517f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_269_n N_A_193_47#_c_908_n 0.00139632f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_281_n N_A_193_47#_c_908_n 5.87167e-19 $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_267_n N_A_193_47#_c_909_n 0.0115307f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_268_n N_A_193_47#_c_909_n 0.00111596f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_269_n N_A_193_47#_c_909_n 0.0369678f $X=5.235 $Y=1.655 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_281_n N_A_193_47#_c_909_n 0.00453285f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_285_n N_A_193_47#_c_909_n 0.00526954f $X=5.295 $Y=1.87 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_288_n N_A_193_47#_c_909_n 3.45729e-19 $X=5.405 $Y=1.74 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_M1030_g N_A_193_47#_c_921_n 0.0130792f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_262_n N_A_193_47#_c_921_n 0.0224153f $X=8.435 $Y=1.32 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_272_n N_A_193_47#_c_921_n 6.57469e-19 $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_M1017_g N_A_193_47#_c_910_n 0.0188272f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_264_n N_A_193_47#_c_910_n 0.0127744f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_398_p N_A_193_47#_c_910_n 0.00850019f $X=0.73 $Y=1.795 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_266_n N_A_193_47#_c_910_n 0.0695916f $X=0.76 $Y=1.235 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_c_281_n N_A_193_47#_c_910_n 0.0124318f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_282_n N_A_193_47#_c_910_n 0.00241841f $X=0.865 $Y=1.87 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_M1010_g N_A_1150_159#_M1001_g 0.0243723f $X=5.31 $Y=2.275
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_269_n N_A_1150_159#_M1001_g 0.00146118f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_283_n N_A_1150_159#_M1001_g 0.0013651f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_c_285_n N_A_1150_159#_M1001_g 0.00196903f $X=5.295 $Y=1.87
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_288_n N_A_1150_159#_M1001_g 0.0206078f $X=5.405 $Y=1.74
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_M1030_g N_A_1150_159#_M1023_g 0.0428173f $X=7.88 $Y=2.275
+ $X2=0 $Y2=0
cc_343 N_A_27_47#_c_283_n N_A_1150_159#_M1023_g 0.00780647f $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_344 N_A_27_47#_c_286_n N_A_1150_159#_M1023_g 0.00131932f $X=7.885 $Y=1.87
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_272_n N_A_1150_159#_M1023_g 0.00605027f $X=7.875 $Y=1.41
+ $X2=0 $Y2=0
cc_346 N_A_27_47#_c_271_n N_A_1150_159#_c_1102_n 0.0189308f $X=7.875 $Y=1.32
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_272_n N_A_1150_159#_c_1102_n 0.00198129f $X=7.875 $Y=1.41
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_283_n N_A_1150_159#_c_1113_n 0.0261908f $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_271_n N_A_1150_159#_c_1105_n 5.17694e-19 $X=7.875 $Y=1.32
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_272_n N_A_1150_159#_c_1105_n 0.00546887f $X=7.875 $Y=1.41
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_283_n N_A_986_413#_M1014_g 0.00324412f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_283_n N_A_986_413#_c_1219_n 2.40114e-19 $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_M1010_g N_A_986_413#_c_1230_n 0.00947181f $X=5.31 $Y=2.275
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_c_281_n N_A_986_413#_c_1230_n 0.00579806f $X=5.15 $Y=1.87
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_c_283_n N_A_986_413#_c_1230_n 0.0054742f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_284_n N_A_986_413#_c_1230_n 0.00117338f $X=5.44 $Y=1.87
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_285_n N_A_986_413#_c_1230_n 0.0279213f $X=5.295 $Y=1.87
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_288_n N_A_986_413#_c_1230_n 7.4902e-19 $X=5.405 $Y=1.74
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_M1006_g N_A_986_413#_c_1236_n 0.00838591f $X=4.99 $Y=0.415
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_267_n N_A_986_413#_c_1236_n 0.0197321f $X=5.15 $Y=0.845
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_268_n N_A_986_413#_c_1236_n 0.00160367f $X=4.98 $Y=0.87
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_267_n N_A_986_413#_c_1221_n 0.0151383f $X=5.15 $Y=0.845
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_269_n N_A_986_413#_c_1221_n 0.024597f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_M1010_g N_A_986_413#_c_1226_n 0.00104479f $X=5.31 $Y=2.275
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_269_n N_A_986_413#_c_1226_n 0.00207816f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_c_283_n N_A_986_413#_c_1226_n 0.0129147f $X=7.74 $Y=1.87 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_284_n N_A_986_413#_c_1226_n 4.13019e-19 $X=5.44 $Y=1.87
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_285_n N_A_986_413#_c_1226_n 0.0255803f $X=5.295 $Y=1.87
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_288_n N_A_986_413#_c_1226_n 6.18409e-19 $X=5.405 $Y=1.74
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_269_n N_A_986_413#_c_1222_n 0.0144717f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_283_n N_A_986_413#_c_1222_n 0.00326146f $X=7.74 $Y=1.87
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_285_n N_A_986_413#_c_1222_n 0.00725124f $X=5.295 $Y=1.87
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_288_n N_A_986_413#_c_1222_n 5.89706e-19 $X=5.405 $Y=1.74
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_M1030_g N_A_1591_413#_c_1339_n 0.00428769f $X=7.88 $Y=2.275
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_c_286_n N_A_1591_413#_c_1339_n 0.0021332f $X=7.885 $Y=1.87
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_c_272_n N_A_1591_413#_c_1339_n 0.00225822f $X=7.875 $Y=1.41
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_M1007_g N_A_1591_413#_c_1342_n 0.0121553f $X=8.51 $Y=0.415
+ $X2=0 $Y2=0
cc_378 N_A_27_47#_M1007_g N_A_1591_413#_c_1328_n 0.00499822f $X=8.51 $Y=0.415
+ $X2=0 $Y2=0
cc_379 N_A_27_47#_c_262_n N_A_1591_413#_c_1337_n 6.71564e-19 $X=8.435 $Y=1.32
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_M1007_g N_A_1591_413#_c_1330_n 0.00301916f $X=8.51 $Y=0.415
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_398_p N_VPWR_M1015_d 6.67509e-19 $X=0.73 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_382 N_A_27_47#_c_282_n N_VPWR_M1015_d 0.00178771f $X=0.865 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_383 N_A_27_47#_c_281_n N_VPWR_M1013_d 0.00132004f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_384 N_A_27_47#_c_283_n N_VPWR_M1001_d 0.00515584f $X=7.74 $Y=1.87 $X2=0 $Y2=0
cc_385 N_A_27_47#_M1000_g N_VPWR_c_1433_n 0.00944765f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_277_n N_VPWR_c_1433_n 0.00346278f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_398_p N_VPWR_c_1433_n 0.013292f $X=0.73 $Y=1.795 $X2=0 $Y2=0
cc_388 N_A_27_47#_c_280_n N_VPWR_c_1433_n 0.012721f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_389 N_A_27_47#_c_282_n N_VPWR_c_1433_n 0.003216f $X=0.865 $Y=1.87 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_281_n N_VPWR_c_1434_n 0.0177398f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_391 N_A_27_47#_c_281_n N_VPWR_c_1435_n 0.0144415f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_392 N_A_27_47#_c_283_n N_VPWR_c_1436_n 0.0124077f $X=7.74 $Y=1.87 $X2=0 $Y2=0
cc_393 N_A_27_47#_M1030_g N_VPWR_c_1438_n 0.00239883f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_283_n N_VPWR_c_1438_n 0.010979f $X=7.74 $Y=1.87 $X2=0 $Y2=0
cc_395 N_A_27_47#_M1000_g N_VPWR_c_1441_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_M1030_g N_VPWR_c_1443_n 0.00429356f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_272_n N_VPWR_c_1443_n 0.00157744f $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_277_n N_VPWR_c_1447_n 0.0018545f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_280_n N_VPWR_c_1447_n 0.0120313f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_400 N_A_27_47#_M1010_g N_VPWR_c_1449_n 0.00375986f $X=5.31 $Y=2.275 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_M1000_g N_VPWR_c_1432_n 0.00534571f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_M1010_g N_VPWR_c_1432_n 0.00556927f $X=5.31 $Y=2.275 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_M1030_g N_VPWR_c_1432_n 0.00573395f $X=7.88 $Y=2.275 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_277_n N_VPWR_c_1432_n 0.00404038f $X=0.615 $Y=1.88 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_c_280_n N_VPWR_c_1432_n 0.00646745f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_281_n N_VPWR_c_1432_n 0.206468f $X=5.15 $Y=1.87 $X2=0 $Y2=0
cc_407 N_A_27_47#_c_282_n N_VPWR_c_1432_n 0.0145601f $X=0.865 $Y=1.87 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_283_n N_VPWR_c_1432_n 0.11007f $X=7.74 $Y=1.87 $X2=0 $Y2=0
cc_409 N_A_27_47#_c_284_n N_VPWR_c_1432_n 0.0144472f $X=5.44 $Y=1.87 $X2=0 $Y2=0
cc_410 N_A_27_47#_c_286_n N_VPWR_c_1432_n 0.0159851f $X=7.885 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_272_n N_VPWR_c_1432_n 0.00101559f $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_281_n N_A_299_47#_c_1596_n 0.020151f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_413 N_A_27_47#_c_281_n N_A_299_47#_c_1588_n 0.00810658f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_281_n N_A_299_47#_c_1598_n 0.0236561f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_281_n N_A_299_47#_c_1589_n 0.00348201f $X=5.15 $Y=1.87 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_c_285_n N_A_299_47#_c_1589_n 0.00630988f $X=5.295 $Y=1.87
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_268_n N_A_299_47#_c_1590_n 3.24335e-19 $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_269_n N_A_299_47#_c_1590_n 0.00462079f $X=5.235 $Y=1.655
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_M1006_g N_A_299_47#_c_1592_n 0.00516494f $X=4.99 $Y=0.415
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_M1006_g N_A_299_47#_c_1594_n 0.00870068f $X=4.99 $Y=0.415
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_c_267_n N_A_299_47#_c_1594_n 0.00702182f $X=5.15 $Y=0.845
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_268_n N_A_299_47#_c_1594_n 0.00130091f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1017_g N_A_299_47#_c_1595_n 0.00143698f $X=0.89 $Y=0.445
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_281_n A_381_369# 0.00298073f $X=5.15 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_425 N_A_27_47#_c_281_n A_729_369# 0.00510983f $X=5.15 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_426 N_A_27_47#_c_264_n N_VGND_M1031_d 0.00164502f $X=0.615 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_427 N_A_27_47#_M1017_g N_VGND_c_1735_n 0.0090859f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_264_n N_VGND_c_1735_n 0.0172929f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_429 N_A_27_47#_c_270_n N_VGND_c_1735_n 5.70216e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_430 N_A_27_47#_M1007_g N_VGND_c_1740_n 0.00155843f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_M1017_g N_VGND_c_1742_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_M1007_g N_VGND_c_1746_n 0.00373071f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_498_p N_VGND_c_1750_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_264_n N_VGND_c_1750_n 0.00243651f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_M1006_g N_VGND_c_1752_n 0.00406674f $X=4.99 $Y=0.415 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_267_n N_VGND_c_1752_n 0.00253275f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_268_n N_VGND_c_1752_n 0.00134958f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_M1031_s N_VGND_c_1754_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_M1017_g N_VGND_c_1754_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_M1006_g N_VGND_c_1754_n 0.00693963f $X=4.99 $Y=0.415 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_M1007_g N_VGND_c_1754_n 0.00568812f $X=8.51 $Y=0.415 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_498_p N_VGND_c_1754_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_264_n N_VGND_c_1754_n 0.00580457f $X=0.615 $Y=0.72 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_c_267_n N_VGND_c_1754_n 0.00206503f $X=5.15 $Y=0.845 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_268_n N_VGND_c_1754_n 0.00141025f $X=4.98 $Y=0.87 $X2=0
+ $Y2=0
cc_446 N_D_M1021_g N_A_423_343#_c_568_n 0.059369f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_447 N_D_c_516_n N_A_423_343#_c_568_n 0.00202148f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_448 D N_A_423_343#_c_568_n 0.00175679f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_449 N_D_c_514_n N_A_423_343#_c_568_n 0.00564261f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_450 D N_A_423_343#_c_564_n 0.00775821f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_451 N_D_c_514_n N_A_423_343#_c_564_n 0.00112085f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_452 N_D_M1002_g N_DE_M1004_g 0.0501357f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_453 D N_DE_M1004_g 3.59802e-19 $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_454 N_D_M1002_g N_DE_c_652_n 0.00609422f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_455 N_D_c_512_n N_DE_c_652_n 0.0121267f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_456 D N_DE_c_652_n 5.46011e-19 $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_457 N_D_M1002_g DE 7.68806e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_458 N_D_c_512_n DE 0.00538864f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_459 D DE 0.0433254f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_460 N_D_c_516_n N_A_193_47#_c_914_n 0.00238342f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_461 D N_A_193_47#_c_914_n 0.0215563f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_462 N_D_c_514_n N_A_193_47#_c_914_n 0.00384385f $X=1.78 $Y=1.145 $X2=0 $Y2=0
cc_463 N_D_M1021_g N_VPWR_c_1434_n 0.00282543f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_464 N_D_M1021_g N_VPWR_c_1441_n 0.00541359f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_465 N_D_M1021_g N_VPWR_c_1432_n 0.00735355f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_466 N_D_M1021_g N_A_299_47#_c_1596_n 0.00949347f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_467 N_D_c_516_n N_A_299_47#_c_1596_n 0.00320688f $X=1.765 $Y=1.65 $X2=0 $Y2=0
cc_468 D N_A_299_47#_c_1596_n 0.00525464f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_469 N_D_M1002_g N_A_299_47#_c_1588_n 0.00738489f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_470 N_D_M1021_g N_A_299_47#_c_1588_n 0.00462667f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_471 N_D_c_512_n N_A_299_47#_c_1588_n 0.00752867f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_472 D N_A_299_47#_c_1588_n 0.0697065f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_473 N_D_M1002_g N_A_299_47#_c_1591_n 7.51093e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_474 N_D_M1002_g N_A_299_47#_c_1593_n 0.00320603f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_475 N_D_c_512_n N_A_299_47#_c_1593_n 0.00203556f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_476 D N_A_299_47#_c_1593_n 0.00827304f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_477 N_D_M1002_g N_A_299_47#_c_1595_n 0.00424642f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_478 N_D_c_512_n N_A_299_47#_c_1595_n 0.00228287f $X=1.765 $Y=1.13 $X2=0 $Y2=0
cc_479 D N_A_299_47#_c_1595_n 0.00347931f $X=1.72 $Y=1.105 $X2=0 $Y2=0
cc_480 N_D_M1002_g N_VGND_c_1736_n 0.00200661f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_481 N_D_M1002_g N_VGND_c_1742_n 0.00539883f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_482 N_D_M1002_g N_VGND_c_1754_n 0.00608889f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_483 N_A_423_343#_c_563_n N_DE_M1004_g 0.00526826f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_484 N_A_423_343#_c_568_n N_DE_c_651_n 0.0080968f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_485 N_A_423_343#_c_564_n N_DE_c_651_n 0.005738f $X=2.932 $Y=1.355 $X2=0 $Y2=0
cc_486 N_A_423_343#_c_567_n N_DE_c_651_n 0.0178991f $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_487 N_A_423_343#_c_568_n N_DE_c_652_n 0.00919986f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_488 N_A_423_343#_c_567_n N_DE_c_652_n 6.99116e-19 $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_489 N_A_423_343#_M1018_g N_DE_M1029_g 0.0148047f $X=3.57 $Y=0.445 $X2=0 $Y2=0
cc_490 N_A_423_343#_c_563_n N_DE_M1029_g 0.00862574f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_491 N_A_423_343#_c_565_n N_DE_M1029_g 0.00220234f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_492 N_A_423_343#_c_566_n N_DE_M1029_g 0.0213224f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_493 N_A_423_343#_c_567_n N_DE_M1029_g 5.67233e-19 $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_494 N_A_423_343#_c_568_n N_DE_c_654_n 0.0152313f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_495 N_A_423_343#_c_564_n N_DE_c_654_n 0.0179184f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_496 N_A_423_343#_c_565_n N_DE_c_654_n 0.00575309f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_497 N_A_423_343#_c_567_n N_DE_c_654_n 0.00317696f $X=2.932 $Y=1.01 $X2=0
+ $Y2=0
cc_498 N_A_423_343#_c_569_n N_DE_M1013_g 0.0105135f $X=2.92 $Y=1.99 $X2=0 $Y2=0
cc_499 N_A_423_343#_c_564_n N_DE_M1013_g 0.00362978f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_500 N_A_423_343#_c_565_n N_DE_c_659_n 0.00580736f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_501 N_A_423_343#_c_566_n N_DE_c_659_n 0.0122629f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_502 N_A_423_343#_c_569_n N_DE_M1016_g 8.04992e-19 $X=2.92 $Y=1.99 $X2=0 $Y2=0
cc_503 N_A_423_343#_c_564_n N_DE_M1016_g 5.26012e-19 $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_504 N_A_423_343#_c_565_n N_DE_c_655_n 0.00305763f $X=3.55 $Y=1.01 $X2=0 $Y2=0
cc_505 N_A_423_343#_c_567_n N_DE_c_655_n 4.2374e-19 $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_506 N_A_423_343#_c_564_n N_DE_c_661_n 0.00610053f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_507 N_A_423_343#_c_568_n DE 0.00845936f $X=2.19 $Y=1.77 $X2=0 $Y2=0
cc_508 N_A_423_343#_c_563_n DE 0.00561932f $X=2.92 $Y=0.51 $X2=0 $Y2=0
cc_509 N_A_423_343#_c_564_n DE 0.0143622f $X=2.932 $Y=1.355 $X2=0 $Y2=0
cc_510 N_A_423_343#_c_567_n DE 0.0240519f $X=2.932 $Y=1.01 $X2=0 $Y2=0
cc_511 N_A_423_343#_M1018_g N_A_791_264#_M1032_g 0.0251313f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_423_343#_c_566_n N_A_791_264#_M1032_g 0.0108934f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_513 N_A_423_343#_M1018_g N_A_791_264#_c_740_n 0.0021118f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_514 N_A_423_343#_c_565_n N_A_791_264#_c_740_n 0.00406567f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_515 N_A_423_343#_c_566_n N_A_791_264#_c_740_n 0.00242559f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_516 N_A_423_343#_M1018_g N_A_791_264#_c_741_n 0.00307938f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_517 N_A_423_343#_c_565_n N_A_791_264#_c_741_n 0.0248957f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_518 N_A_423_343#_c_566_n N_A_791_264#_c_741_n 0.00233652f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_519 N_A_423_343#_c_568_n N_A_193_47#_c_914_n 0.00463103f $X=2.19 $Y=1.77
+ $X2=0 $Y2=0
cc_520 N_A_423_343#_c_569_n N_A_193_47#_c_914_n 3.18139e-19 $X=2.92 $Y=1.99
+ $X2=0 $Y2=0
cc_521 N_A_423_343#_c_564_n N_A_193_47#_c_914_n 0.0327297f $X=2.932 $Y=1.355
+ $X2=0 $Y2=0
cc_522 N_A_423_343#_c_565_n N_A_193_47#_c_914_n 0.0177671f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_523 N_A_423_343#_c_566_n N_A_193_47#_c_914_n 0.00228465f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_524 N_A_423_343#_c_568_n N_VPWR_c_1434_n 0.0251559f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_525 N_A_423_343#_c_569_n N_VPWR_c_1434_n 0.0405714f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_526 N_A_423_343#_c_564_n N_VPWR_c_1434_n 0.00458578f $X=2.932 $Y=1.355 $X2=0
+ $Y2=0
cc_527 N_A_423_343#_c_569_n N_VPWR_c_1435_n 0.0418939f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_528 N_A_423_343#_c_565_n N_VPWR_c_1435_n 0.00271398f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_529 N_A_423_343#_c_568_n N_VPWR_c_1441_n 0.0046653f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_530 N_A_423_343#_c_569_n N_VPWR_c_1448_n 0.0167964f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_531 N_A_423_343#_M1013_s N_VPWR_c_1432_n 0.00173907f $X=2.795 $Y=1.845 $X2=0
+ $Y2=0
cc_532 N_A_423_343#_c_568_n N_VPWR_c_1432_n 0.00430483f $X=2.19 $Y=1.77 $X2=0
+ $Y2=0
cc_533 N_A_423_343#_c_569_n N_VPWR_c_1432_n 0.00581267f $X=2.92 $Y=1.99 $X2=0
+ $Y2=0
cc_534 N_A_423_343#_c_568_n N_A_299_47#_c_1596_n 0.00159809f $X=2.19 $Y=1.77
+ $X2=0 $Y2=0
cc_535 N_A_423_343#_M1018_g N_A_299_47#_c_1592_n 2.04373e-19 $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_536 N_A_423_343#_M1029_s N_A_299_47#_c_1593_n 6.77802e-19 $X=2.795 $Y=0.235
+ $X2=0 $Y2=0
cc_537 N_A_423_343#_M1018_g N_A_299_47#_c_1593_n 0.00414801f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_538 N_A_423_343#_c_563_n N_A_299_47#_c_1593_n 0.0183276f $X=2.92 $Y=0.51
+ $X2=0 $Y2=0
cc_539 N_A_423_343#_c_565_n N_A_299_47#_c_1593_n 0.0107001f $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_540 N_A_423_343#_c_566_n N_A_299_47#_c_1593_n 9.48498e-19 $X=3.55 $Y=1.01
+ $X2=0 $Y2=0
cc_541 N_A_423_343#_c_567_n N_A_299_47#_c_1593_n 0.00351536f $X=2.932 $Y=1.01
+ $X2=0 $Y2=0
cc_542 N_A_423_343#_M1018_g N_A_299_47#_c_1594_n 0.00155158f $X=3.57 $Y=0.445
+ $X2=0 $Y2=0
cc_543 N_A_423_343#_c_563_n N_VGND_c_1736_n 0.0164318f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_544 N_A_423_343#_M1018_g N_VGND_c_1737_n 0.0113899f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_545 N_A_423_343#_c_563_n N_VGND_c_1737_n 0.0148662f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_546 N_A_423_343#_c_565_n N_VGND_c_1737_n 0.0151977f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_547 N_A_423_343#_c_566_n N_VGND_c_1737_n 0.00159308f $X=3.55 $Y=1.01 $X2=0
+ $Y2=0
cc_548 N_A_423_343#_c_563_n N_VGND_c_1751_n 0.0154917f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_549 N_A_423_343#_M1018_g N_VGND_c_1752_n 0.00505556f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_550 N_A_423_343#_M1029_s N_VGND_c_1754_n 0.00120778f $X=2.795 $Y=0.235 $X2=0
+ $Y2=0
cc_551 N_A_423_343#_M1018_g N_VGND_c_1754_n 0.00379888f $X=3.57 $Y=0.445 $X2=0
+ $Y2=0
cc_552 N_A_423_343#_c_563_n N_VGND_c_1754_n 0.00215984f $X=2.92 $Y=0.51 $X2=0
+ $Y2=0
cc_553 N_DE_M1016_g N_A_791_264#_M1026_g 0.033024f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_554 N_DE_c_654_n N_A_791_264#_c_751_n 0.00334239f $X=3.13 $Y=1.46 $X2=0 $Y2=0
cc_555 N_DE_c_659_n N_A_791_264#_c_751_n 0.00386505f $X=3.495 $Y=1.535 $X2=0
+ $Y2=0
cc_556 N_DE_c_659_n N_A_791_264#_c_752_n 0.00786818f $X=3.495 $Y=1.535 $X2=0
+ $Y2=0
cc_557 N_DE_c_654_n N_A_791_264#_c_741_n 0.00317814f $X=3.13 $Y=1.46 $X2=0 $Y2=0
cc_558 N_DE_c_659_n N_A_193_47#_c_914_n 0.0079741f $X=3.495 $Y=1.535 $X2=0 $Y2=0
cc_559 N_DE_c_661_n N_A_193_47#_c_914_n 0.00255711f $X=3.13 $Y=1.535 $X2=0 $Y2=0
cc_560 DE N_A_193_47#_c_914_n 0.0181093f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_561 N_DE_M1013_g N_VPWR_c_1434_n 0.00292738f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_562 DE N_VPWR_c_1434_n 0.00131185f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_563 N_DE_M1013_g N_VPWR_c_1435_n 0.00567389f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_564 N_DE_c_659_n N_VPWR_c_1435_n 0.00241702f $X=3.495 $Y=1.535 $X2=0 $Y2=0
cc_565 N_DE_M1016_g N_VPWR_c_1435_n 0.00345066f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_566 N_DE_M1013_g N_VPWR_c_1448_n 0.00542953f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_567 N_DE_M1016_g N_VPWR_c_1449_n 0.00585385f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_568 N_DE_M1013_g N_VPWR_c_1432_n 0.00739796f $X=3.13 $Y=2.165 $X2=0 $Y2=0
cc_569 N_DE_M1016_g N_VPWR_c_1432_n 0.00652437f $X=3.57 $Y=2.165 $X2=0 $Y2=0
cc_570 N_DE_M1016_g N_A_299_47#_c_1598_n 0.00208296f $X=3.57 $Y=2.165 $X2=0
+ $Y2=0
cc_571 N_DE_M1004_g N_A_299_47#_c_1593_n 0.00328866f $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_572 N_DE_c_651_n N_A_299_47#_c_1593_n 0.00449574f $X=3.055 $Y=0.925 $X2=0
+ $Y2=0
cc_573 N_DE_M1029_g N_A_299_47#_c_1593_n 0.00212954f $X=3.13 $Y=0.445 $X2=0
+ $Y2=0
cc_574 DE N_A_299_47#_c_1593_n 0.014806f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_575 N_DE_M1004_g N_A_299_47#_c_1595_n 7.72933e-19 $X=2.19 $Y=0.445 $X2=0
+ $Y2=0
cc_576 N_DE_M1004_g N_VGND_c_1736_n 0.0103332f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_577 N_DE_c_651_n N_VGND_c_1736_n 5.49262e-19 $X=3.055 $Y=0.925 $X2=0 $Y2=0
cc_578 N_DE_c_652_n N_VGND_c_1736_n 9.86308e-19 $X=2.455 $Y=0.925 $X2=0 $Y2=0
cc_579 N_DE_M1029_g N_VGND_c_1736_n 0.00200593f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_580 DE N_VGND_c_1736_n 0.0147118f $X=2.13 $Y=0.765 $X2=0 $Y2=0
cc_581 N_DE_M1029_g N_VGND_c_1737_n 0.00765346f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_582 N_DE_M1004_g N_VGND_c_1742_n 0.0046653f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_583 N_DE_M1029_g N_VGND_c_1751_n 0.00505556f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_584 N_DE_M1004_g N_VGND_c_1754_n 0.00313929f $X=2.19 $Y=0.445 $X2=0 $Y2=0
cc_585 N_DE_M1029_g N_VGND_c_1754_n 0.00491778f $X=3.13 $Y=0.445 $X2=0 $Y2=0
cc_586 N_A_791_264#_M1026_g N_A_193_47#_M1009_g 0.00900582f $X=4.08 $Y=2.165
+ $X2=0 $Y2=0
cc_587 N_A_791_264#_c_752_n N_A_193_47#_M1009_g 0.00336172f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_588 N_A_791_264#_c_739_n N_A_193_47#_c_902_n 4.65473e-19 $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_589 N_A_791_264#_c_739_n N_A_193_47#_M1028_g 0.00493455f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_590 N_A_791_264#_c_749_n N_A_193_47#_M1024_g 0.0199779f $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_591 N_A_791_264#_M1020_g N_A_193_47#_c_905_n 3.66194e-19 $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_592 N_A_791_264#_c_739_n N_A_193_47#_c_905_n 0.0311489f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_593 N_A_791_264#_c_739_n N_A_193_47#_c_906_n 0.00343724f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_594 N_A_791_264#_c_751_n N_A_193_47#_c_914_n 0.0212f $X=4.09 $Y=1.485 $X2=0
+ $Y2=0
cc_595 N_A_791_264#_c_752_n N_A_193_47#_c_914_n 0.00192918f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_596 N_A_791_264#_c_739_n N_A_193_47#_c_914_n 0.0309696f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_597 N_A_791_264#_c_740_n N_A_193_47#_c_914_n 0.013239f $X=4.035 $Y=0.85 $X2=0
+ $Y2=0
cc_598 N_A_791_264#_c_741_n N_A_193_47#_c_914_n 3.15466e-19 $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_599 N_A_791_264#_c_739_n N_A_193_47#_c_916_n 0.132905f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_600 N_A_791_264#_c_739_n N_A_193_47#_c_917_n 0.0130915f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_601 N_A_791_264#_c_739_n N_A_193_47#_c_960_n 0.012252f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_602 N_A_791_264#_c_749_n N_A_193_47#_c_907_n 7.03497e-19 $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_603 N_A_791_264#_M1032_g N_A_193_47#_c_908_n 0.00150065f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_604 N_A_791_264#_c_752_n N_A_193_47#_c_908_n 0.00311382f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_605 N_A_791_264#_c_739_n N_A_193_47#_c_908_n 0.00127009f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_606 N_A_791_264#_M1032_g N_A_193_47#_c_909_n 7.03902e-19 $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_607 N_A_791_264#_c_739_n N_A_193_47#_c_909_n 0.0014675f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_608 N_A_791_264#_c_749_n N_A_193_47#_c_921_n 0.0137111f $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_609 N_A_791_264#_c_739_n N_A_1150_159#_M1011_g 0.00577171f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_610 N_A_791_264#_c_739_n N_A_1150_159#_c_1101_n 0.00619242f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_611 N_A_791_264#_c_739_n N_A_1150_159#_c_1103_n 0.0564626f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_612 N_A_791_264#_c_739_n N_A_1150_159#_c_1105_n 0.012477f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_613 N_A_791_264#_c_739_n N_A_1150_159#_c_1107_n 0.0112362f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_614 N_A_791_264#_c_739_n N_A_1150_159#_c_1108_n 0.00300444f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_615 N_A_791_264#_c_739_n N_A_986_413#_c_1236_n 0.00659708f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_616 N_A_791_264#_c_739_n N_A_986_413#_c_1221_n 0.0152331f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_617 N_A_791_264#_c_739_n N_A_986_413#_c_1222_n 0.00619733f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_618 N_A_791_264#_c_737_n N_A_1591_413#_M1012_g 0.00561498f $X=9.715 $Y=0.385
+ $X2=0 $Y2=0
cc_619 N_A_791_264#_c_738_n N_A_1591_413#_M1012_g 0.00477121f $X=9.715 $Y=0.825
+ $X2=0 $Y2=0
cc_620 N_A_791_264#_c_742_n N_A_1591_413#_M1012_g 0.00517962f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_621 N_A_791_264#_c_743_n N_A_1591_413#_M1012_g 0.0052888f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_622 N_A_791_264#_c_749_n N_A_1591_413#_M1027_g 0.00345271f $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_623 N_A_791_264#_c_750_n N_A_1591_413#_M1027_g 0.00613006f $X=9.705 $Y=1.99
+ $X2=0 $Y2=0
cc_624 N_A_791_264#_c_753_n N_A_1591_413#_M1027_g 0.0104703f $X=9.71 $Y=1.717
+ $X2=0 $Y2=0
cc_625 N_A_791_264#_c_743_n N_A_1591_413#_M1027_g 0.00721223f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_626 N_A_791_264#_c_737_n N_A_1591_413#_c_1324_n 5.51494e-19 $X=9.715 $Y=0.385
+ $X2=0 $Y2=0
cc_627 N_A_791_264#_c_742_n N_A_1591_413#_c_1324_n 3.16115e-19 $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_628 N_A_791_264#_c_743_n N_A_1591_413#_M1005_g 4.45214e-19 $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_629 N_A_791_264#_M1020_g N_A_1591_413#_c_1325_n 0.0191523f $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_630 N_A_791_264#_c_748_n N_A_1591_413#_c_1325_n 0.00609226f $X=9.54 $Y=1.717
+ $X2=0 $Y2=0
cc_631 N_A_791_264#_c_753_n N_A_1591_413#_c_1325_n 0.00641947f $X=9.71 $Y=1.717
+ $X2=0 $Y2=0
cc_632 N_A_791_264#_c_738_n N_A_1591_413#_c_1325_n 0.00500691f $X=9.715 $Y=0.825
+ $X2=0 $Y2=0
cc_633 N_A_791_264#_c_739_n N_A_1591_413#_c_1325_n 0.00892528f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_634 N_A_791_264#_c_742_n N_A_1591_413#_c_1325_n 0.00143362f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_635 N_A_791_264#_c_743_n N_A_1591_413#_c_1325_n 0.0170494f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_636 N_A_791_264#_c_743_n N_A_1591_413#_c_1326_n 0.00983534f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_637 N_A_791_264#_M1019_g N_A_1591_413#_c_1339_n 0.00510852f $X=8.87 $Y=2.275
+ $X2=0 $Y2=0
cc_638 N_A_791_264#_M1020_g N_A_1591_413#_c_1342_n 0.00188481f $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_639 N_A_791_264#_c_739_n N_A_1591_413#_c_1342_n 0.00605628f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_640 N_A_791_264#_M1020_g N_A_1591_413#_c_1328_n 0.0088172f $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_641 N_A_791_264#_c_739_n N_A_1591_413#_c_1328_n 0.0223085f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_642 N_A_791_264#_M1019_g N_A_1591_413#_c_1337_n 0.0120201f $X=8.87 $Y=2.275
+ $X2=0 $Y2=0
cc_643 N_A_791_264#_M1020_g N_A_1591_413#_c_1337_n 0.00751613f $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_644 N_A_791_264#_c_748_n N_A_1591_413#_c_1337_n 0.0282373f $X=9.54 $Y=1.717
+ $X2=0 $Y2=0
cc_645 N_A_791_264#_c_749_n N_A_1591_413#_c_1337_n 0.0079118f $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_646 N_A_791_264#_M1020_g N_A_1591_413#_c_1329_n 0.0183255f $X=8.985 $Y=0.445
+ $X2=0 $Y2=0
cc_647 N_A_791_264#_c_748_n N_A_1591_413#_c_1329_n 0.0359416f $X=9.54 $Y=1.717
+ $X2=0 $Y2=0
cc_648 N_A_791_264#_c_749_n N_A_1591_413#_c_1329_n 0.00495398f $X=9.065 $Y=1.74
+ $X2=0 $Y2=0
cc_649 N_A_791_264#_c_739_n N_A_1591_413#_c_1329_n 0.0291683f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_650 N_A_791_264#_c_743_n N_A_1591_413#_c_1329_n 0.0240437f $X=9.785 $Y=0.85
+ $X2=0 $Y2=0
cc_651 N_A_791_264#_M1019_g N_VPWR_c_1439_n 0.00462747f $X=8.87 $Y=2.275 $X2=0
+ $Y2=0
cc_652 N_A_791_264#_c_748_n N_VPWR_c_1439_n 0.0155824f $X=9.54 $Y=1.717 $X2=0
+ $Y2=0
cc_653 N_A_791_264#_c_749_n N_VPWR_c_1439_n 0.00514677f $X=9.065 $Y=1.74 $X2=0
+ $Y2=0
cc_654 N_A_791_264#_c_750_n N_VPWR_c_1439_n 0.0182471f $X=9.705 $Y=1.99 $X2=0
+ $Y2=0
cc_655 N_A_791_264#_c_753_n N_VPWR_c_1440_n 0.0283369f $X=9.71 $Y=1.717 $X2=0
+ $Y2=0
cc_656 N_A_791_264#_c_743_n N_VPWR_c_1440_n 0.00515656f $X=9.785 $Y=0.85 $X2=0
+ $Y2=0
cc_657 N_A_791_264#_M1019_g N_VPWR_c_1443_n 0.00564808f $X=8.87 $Y=2.275 $X2=0
+ $Y2=0
cc_658 N_A_791_264#_c_750_n N_VPWR_c_1445_n 0.0217414f $X=9.705 $Y=1.99 $X2=0
+ $Y2=0
cc_659 N_A_791_264#_M1026_g N_VPWR_c_1449_n 0.00541359f $X=4.08 $Y=2.165 $X2=0
+ $Y2=0
cc_660 N_A_791_264#_M1027_s N_VPWR_c_1432_n 0.00217517f $X=9.58 $Y=1.845 $X2=0
+ $Y2=0
cc_661 N_A_791_264#_M1026_g N_VPWR_c_1432_n 0.00707761f $X=4.08 $Y=2.165 $X2=0
+ $Y2=0
cc_662 N_A_791_264#_M1019_g N_VPWR_c_1432_n 0.0117199f $X=8.87 $Y=2.275 $X2=0
+ $Y2=0
cc_663 N_A_791_264#_c_748_n N_VPWR_c_1432_n 0.0122998f $X=9.54 $Y=1.717 $X2=0
+ $Y2=0
cc_664 N_A_791_264#_c_749_n N_VPWR_c_1432_n 8.92751e-19 $X=9.065 $Y=1.74 $X2=0
+ $Y2=0
cc_665 N_A_791_264#_c_750_n N_VPWR_c_1432_n 0.0128119f $X=9.705 $Y=1.99 $X2=0
+ $Y2=0
cc_666 N_A_791_264#_M1026_g N_A_299_47#_c_1598_n 0.0133737f $X=4.08 $Y=2.165
+ $X2=0 $Y2=0
cc_667 N_A_791_264#_c_751_n N_A_299_47#_c_1598_n 0.00318555f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_668 N_A_791_264#_c_752_n N_A_299_47#_c_1598_n 0.00178853f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_669 N_A_791_264#_M1032_g N_A_299_47#_c_1589_n 0.0013593f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_670 N_A_791_264#_M1026_g N_A_299_47#_c_1589_n 0.0027891f $X=4.08 $Y=2.165
+ $X2=0 $Y2=0
cc_671 N_A_791_264#_c_751_n N_A_299_47#_c_1589_n 0.0237025f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_672 N_A_791_264#_c_752_n N_A_299_47#_c_1589_n 0.00289234f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_673 N_A_791_264#_c_741_n N_A_299_47#_c_1589_n 0.00525839f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_674 N_A_791_264#_M1032_g N_A_299_47#_c_1590_n 0.00517267f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_675 N_A_791_264#_c_751_n N_A_299_47#_c_1590_n 0.00212358f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_676 N_A_791_264#_c_752_n N_A_299_47#_c_1590_n 0.00197416f $X=4.09 $Y=1.485
+ $X2=0 $Y2=0
cc_677 N_A_791_264#_c_739_n N_A_299_47#_c_1590_n 0.00430154f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_678 N_A_791_264#_M1032_g N_A_299_47#_c_1592_n 0.00100352f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_679 N_A_791_264#_c_739_n N_A_299_47#_c_1592_n 0.0250725f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_680 N_A_791_264#_M1032_g N_A_299_47#_c_1593_n 0.00367101f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_681 N_A_791_264#_c_739_n N_A_299_47#_c_1593_n 0.00735691f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_682 N_A_791_264#_c_740_n N_A_299_47#_c_1593_n 0.0273168f $X=4.035 $Y=0.85
+ $X2=0 $Y2=0
cc_683 N_A_791_264#_c_741_n N_A_299_47#_c_1593_n 0.00264974f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_684 N_A_791_264#_M1032_g N_A_299_47#_c_1594_n 0.0148374f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_685 N_A_791_264#_c_739_n N_A_299_47#_c_1594_n 0.0181297f $X=9.64 $Y=0.85
+ $X2=0 $Y2=0
cc_686 N_A_791_264#_c_740_n N_A_299_47#_c_1594_n 0.00238395f $X=4.035 $Y=0.85
+ $X2=0 $Y2=0
cc_687 N_A_791_264#_c_741_n N_A_299_47#_c_1594_n 0.0329237f $X=3.89 $Y=0.85
+ $X2=0 $Y2=0
cc_688 N_A_791_264#_c_742_n N_Q_c_1718_n 0.00151602f $X=9.785 $Y=0.85 $X2=0
+ $Y2=0
cc_689 N_A_791_264#_c_743_n N_Q_c_1718_n 0.0137869f $X=9.785 $Y=0.85 $X2=0 $Y2=0
cc_690 N_A_791_264#_M1032_g N_VGND_c_1737_n 0.00210691f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_691 N_A_791_264#_c_739_n N_VGND_c_1738_n 0.00209284f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_692 N_A_791_264#_c_739_n N_VGND_c_1739_n 0.00448688f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_693 N_A_791_264#_M1020_g N_VGND_c_1740_n 0.010757f $X=8.985 $Y=0.445 $X2=0
+ $Y2=0
cc_694 N_A_791_264#_c_737_n N_VGND_c_1740_n 0.0246268f $X=9.715 $Y=0.385 $X2=0
+ $Y2=0
cc_695 N_A_791_264#_c_739_n N_VGND_c_1740_n 0.00490532f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_696 N_A_791_264#_c_737_n N_VGND_c_1741_n 0.0299916f $X=9.715 $Y=0.385 $X2=0
+ $Y2=0
cc_697 N_A_791_264#_c_742_n N_VGND_c_1741_n 0.00495351f $X=9.785 $Y=0.85 $X2=0
+ $Y2=0
cc_698 N_A_791_264#_M1020_g N_VGND_c_1746_n 0.00544582f $X=8.985 $Y=0.445 $X2=0
+ $Y2=0
cc_699 N_A_791_264#_c_737_n N_VGND_c_1748_n 0.016199f $X=9.715 $Y=0.385 $X2=0
+ $Y2=0
cc_700 N_A_791_264#_M1032_g N_VGND_c_1752_n 0.00571722f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_701 N_A_791_264#_c_741_n N_VGND_c_1752_n 0.00260398f $X=3.89 $Y=0.85 $X2=0
+ $Y2=0
cc_702 N_A_791_264#_M1012_s N_VGND_c_1754_n 0.00169299f $X=9.59 $Y=0.235 $X2=0
+ $Y2=0
cc_703 N_A_791_264#_M1032_g N_VGND_c_1754_n 0.0068705f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_704 N_A_791_264#_M1020_g N_VGND_c_1754_n 0.00524744f $X=8.985 $Y=0.445 $X2=0
+ $Y2=0
cc_705 N_A_791_264#_c_737_n N_VGND_c_1754_n 0.00555624f $X=9.715 $Y=0.385 $X2=0
+ $Y2=0
cc_706 N_A_791_264#_c_739_n N_VGND_c_1754_n 0.249572f $X=9.64 $Y=0.85 $X2=0
+ $Y2=0
cc_707 N_A_791_264#_c_742_n N_VGND_c_1754_n 0.0146996f $X=9.785 $Y=0.85 $X2=0
+ $Y2=0
cc_708 N_A_193_47#_c_902_n N_A_1150_159#_M1001_g 0.0138337f $X=5.355 $Y=1.29
+ $X2=0 $Y2=0
cc_709 N_A_193_47#_c_916_n N_A_1150_159#_M1001_g 0.00185536f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_710 N_A_193_47#_c_908_n N_A_1150_159#_M1001_g 0.00119103f $X=4.88 $Y=1.29
+ $X2=0 $Y2=0
cc_711 N_A_193_47#_M1028_g N_A_1150_159#_M1033_g 0.0189994f $X=5.43 $Y=0.415
+ $X2=0 $Y2=0
cc_712 N_A_193_47#_c_916_n N_A_1150_159#_M1023_g 0.00722181f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_713 N_A_193_47#_c_904_n N_A_1150_159#_M1011_g 0.0181756f $X=7.98 $Y=0.705
+ $X2=0 $Y2=0
cc_714 N_A_193_47#_c_905_n N_A_1150_159#_M1011_g 0.00208129f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_715 N_A_193_47#_c_906_n N_A_1150_159#_c_1101_n 0.0181756f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_716 N_A_193_47#_c_916_n N_A_1150_159#_c_1101_n 0.00123775f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_717 N_A_193_47#_c_907_n N_A_1150_159#_c_1101_n 2.51226e-19 $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_718 N_A_193_47#_c_916_n N_A_1150_159#_c_1102_n 0.00252648f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_719 N_A_193_47#_c_916_n N_A_1150_159#_c_1103_n 0.00787458f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_720 N_A_193_47#_c_916_n N_A_1150_159#_c_1113_n 0.0260184f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_721 N_A_193_47#_c_916_n N_A_1150_159#_c_1105_n 0.0182403f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_722 N_A_193_47#_c_907_n N_A_1150_159#_c_1106_n 0.00478379f $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_723 N_A_193_47#_c_916_n N_A_1150_159#_c_1107_n 7.49207e-19 $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_724 N_A_193_47#_M1028_g N_A_1150_159#_c_1108_n 0.0138337f $X=5.43 $Y=0.415
+ $X2=0 $Y2=0
cc_725 N_A_193_47#_c_916_n N_A_986_413#_M1014_g 0.00174404f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_726 N_A_193_47#_c_916_n N_A_986_413#_c_1219_n 8.02119e-19 $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_727 N_A_193_47#_c_916_n N_A_986_413#_c_1220_n 0.00120348f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_728 N_A_193_47#_M1009_g N_A_986_413#_c_1230_n 0.00390359f $X=4.855 $Y=2.275
+ $X2=0 $Y2=0
cc_729 N_A_193_47#_c_908_n N_A_986_413#_c_1230_n 9.99101e-19 $X=4.88 $Y=1.29
+ $X2=0 $Y2=0
cc_730 N_A_193_47#_c_909_n N_A_986_413#_c_1230_n 7.25987e-19 $X=4.88 $Y=1.35
+ $X2=0 $Y2=0
cc_731 N_A_193_47#_c_902_n N_A_986_413#_c_1236_n 4.77975e-19 $X=5.355 $Y=1.29
+ $X2=0 $Y2=0
cc_732 N_A_193_47#_M1028_g N_A_986_413#_c_1236_n 0.0112915f $X=5.43 $Y=0.415
+ $X2=0 $Y2=0
cc_733 N_A_193_47#_M1028_g N_A_986_413#_c_1221_n 0.00847049f $X=5.43 $Y=0.415
+ $X2=0 $Y2=0
cc_734 N_A_193_47#_c_916_n N_A_986_413#_c_1226_n 0.0041331f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_735 N_A_193_47#_c_902_n N_A_986_413#_c_1222_n 5.3564e-19 $X=5.355 $Y=1.29
+ $X2=0 $Y2=0
cc_736 N_A_193_47#_c_916_n N_A_986_413#_c_1222_n 0.0376331f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_737 N_A_193_47#_M1024_g N_A_1591_413#_c_1339_n 0.00963552f $X=8.3 $Y=2.275
+ $X2=0 $Y2=0
cc_738 N_A_193_47#_c_916_n N_A_1591_413#_c_1339_n 0.00391921f $X=8.16 $Y=1.53
+ $X2=0 $Y2=0
cc_739 N_A_193_47#_c_960_n N_A_1591_413#_c_1339_n 0.00103138f $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_740 N_A_193_47#_c_907_n N_A_1591_413#_c_1339_n 0.0198599f $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_921_n N_A_1591_413#_c_1339_n 0.00303787f $X=8.385 $Y=1.74
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_c_904_n N_A_1591_413#_c_1342_n 0.00459251f $X=7.98 $Y=0.705
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_905_n N_A_1591_413#_c_1342_n 0.0278532f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_744 N_A_193_47#_c_906_n N_A_1591_413#_c_1342_n 0.00108492f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_745 N_A_193_47#_c_905_n N_A_1591_413#_c_1328_n 0.0210561f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_746 N_A_193_47#_M1024_g N_A_1591_413#_c_1337_n 0.00365921f $X=8.3 $Y=2.275
+ $X2=0 $Y2=0
cc_747 N_A_193_47#_c_960_n N_A_1591_413#_c_1337_n 0.00161073f $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_748 N_A_193_47#_c_907_n N_A_1591_413#_c_1337_n 0.0495718f $X=8.305 $Y=1.53
+ $X2=0 $Y2=0
cc_749 N_A_193_47#_c_921_n N_A_1591_413#_c_1337_n 0.00182086f $X=8.385 $Y=1.74
+ $X2=0 $Y2=0
cc_750 N_A_193_47#_c_905_n N_A_1591_413#_c_1330_n 0.0277807f $X=8.09 $Y=0.87
+ $X2=0 $Y2=0
cc_751 N_A_193_47#_c_910_n N_VPWR_c_1433_n 0.012721f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_752 N_A_193_47#_c_914_n N_VPWR_c_1434_n 0.00138291f $X=4.74 $Y=1.53 $X2=0
+ $Y2=0
cc_753 N_A_193_47#_c_914_n N_VPWR_c_1435_n 7.40558e-19 $X=4.74 $Y=1.53 $X2=0
+ $Y2=0
cc_754 N_A_193_47#_c_916_n N_VPWR_c_1436_n 8.15834e-19 $X=8.16 $Y=1.53 $X2=0
+ $Y2=0
cc_755 N_A_193_47#_c_910_n N_VPWR_c_1441_n 0.0120448f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_756 N_A_193_47#_M1024_g N_VPWR_c_1443_n 0.0037981f $X=8.3 $Y=2.275 $X2=0
+ $Y2=0
cc_757 N_A_193_47#_M1009_g N_VPWR_c_1449_n 0.00564445f $X=4.855 $Y=2.275 $X2=0
+ $Y2=0
cc_758 N_A_193_47#_M1009_g N_VPWR_c_1432_n 0.00713447f $X=4.855 $Y=2.275 $X2=0
+ $Y2=0
cc_759 N_A_193_47#_M1024_g N_VPWR_c_1432_n 0.0057367f $X=8.3 $Y=2.275 $X2=0
+ $Y2=0
cc_760 N_A_193_47#_c_910_n N_VPWR_c_1432_n 0.00308197f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_761 N_A_193_47#_c_914_n N_A_299_47#_c_1596_n 0.0010389f $X=4.74 $Y=1.53 $X2=0
+ $Y2=0
cc_762 N_A_193_47#_c_914_n N_A_299_47#_c_1588_n 0.0170784f $X=4.74 $Y=1.53 $X2=0
+ $Y2=0
cc_763 N_A_193_47#_c_915_n N_A_299_47#_c_1588_n 0.00275409f $X=1.245 $Y=1.53
+ $X2=0 $Y2=0
cc_764 N_A_193_47#_c_910_n N_A_299_47#_c_1588_n 0.145237f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_765 N_A_193_47#_M1009_g N_A_299_47#_c_1598_n 0.00734257f $X=4.855 $Y=2.275
+ $X2=0 $Y2=0
cc_766 N_A_193_47#_c_914_n N_A_299_47#_c_1598_n 8.15261e-19 $X=4.74 $Y=1.53
+ $X2=0 $Y2=0
cc_767 N_A_193_47#_M1009_g N_A_299_47#_c_1589_n 0.00499579f $X=4.855 $Y=2.275
+ $X2=0 $Y2=0
cc_768 N_A_193_47#_c_914_n N_A_299_47#_c_1589_n 0.0134484f $X=4.74 $Y=1.53 $X2=0
+ $Y2=0
cc_769 N_A_193_47#_c_917_n N_A_299_47#_c_1589_n 0.00238903f $X=5.03 $Y=1.53
+ $X2=0 $Y2=0
cc_770 N_A_193_47#_c_908_n N_A_299_47#_c_1589_n 0.00273481f $X=4.88 $Y=1.29
+ $X2=0 $Y2=0
cc_771 N_A_193_47#_c_914_n N_A_299_47#_c_1590_n 0.00275532f $X=4.74 $Y=1.53
+ $X2=0 $Y2=0
cc_772 N_A_193_47#_c_909_n N_A_299_47#_c_1590_n 0.0276847f $X=4.88 $Y=1.35 $X2=0
+ $Y2=0
cc_773 N_A_193_47#_c_910_n N_A_299_47#_c_1591_n 0.00796831f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_774 N_A_193_47#_c_910_n N_A_299_47#_c_1595_n 0.0117897f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_775 N_A_193_47#_M1028_g N_VGND_c_1738_n 0.00140802f $X=5.43 $Y=0.415 $X2=0
+ $Y2=0
cc_776 N_A_193_47#_c_904_n N_VGND_c_1739_n 0.00237285f $X=7.98 $Y=0.705 $X2=0
+ $Y2=0
cc_777 N_A_193_47#_c_910_n N_VGND_c_1742_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_778 N_A_193_47#_c_904_n N_VGND_c_1746_n 0.00523869f $X=7.98 $Y=0.705 $X2=0
+ $Y2=0
cc_779 N_A_193_47#_c_905_n N_VGND_c_1746_n 2.78187e-19 $X=8.09 $Y=0.87 $X2=0
+ $Y2=0
cc_780 N_A_193_47#_M1028_g N_VGND_c_1752_n 0.00357877f $X=5.43 $Y=0.415 $X2=0
+ $Y2=0
cc_781 N_A_193_47#_M1017_d N_VGND_c_1754_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_782 N_A_193_47#_M1028_g N_VGND_c_1754_n 0.00553273f $X=5.43 $Y=0.415 $X2=0
+ $Y2=0
cc_783 N_A_193_47#_c_904_n N_VGND_c_1754_n 0.00656556f $X=7.98 $Y=0.705 $X2=0
+ $Y2=0
cc_784 N_A_193_47#_c_905_n N_VGND_c_1754_n 0.00106975f $X=8.09 $Y=0.87 $X2=0
+ $Y2=0
cc_785 N_A_193_47#_c_910_n N_VGND_c_1754_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_786 N_A_1150_159#_c_1103_n N_A_986_413#_c_1216_n 0.00661847f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_787 N_A_1150_159#_c_1105_n N_A_986_413#_c_1216_n 2.83663e-19 $X=7.36 $Y=1.21
+ $X2=0 $Y2=0
cc_788 N_A_1150_159#_c_1106_n N_A_986_413#_c_1216_n 0.00149495f $X=7.36 $Y=1.21
+ $X2=0 $Y2=0
cc_789 N_A_1150_159#_M1001_g N_A_986_413#_M1014_g 0.0142214f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_790 N_A_1150_159#_c_1113_n N_A_986_413#_M1014_g 0.0168148f $X=6.695 $Y=1.88
+ $X2=0 $Y2=0
cc_791 N_A_1150_159#_M1033_g N_A_986_413#_c_1217_n 0.0121471f $X=5.96 $Y=0.445
+ $X2=0 $Y2=0
cc_792 N_A_1150_159#_c_1101_n N_A_986_413#_c_1217_n 0.00145117f $X=7.397
+ $Y=1.045 $X2=0 $Y2=0
cc_793 N_A_1150_159#_c_1103_n N_A_986_413#_c_1217_n 0.00790103f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_794 N_A_1150_159#_c_1104_n N_A_986_413#_c_1217_n 0.0110908f $X=6.765 $Y=0.39
+ $X2=0 $Y2=0
cc_795 N_A_1150_159#_c_1108_n N_A_986_413#_c_1217_n 0.00500472f $X=5.96 $Y=0.93
+ $X2=0 $Y2=0
cc_796 N_A_1150_159#_M1001_g N_A_986_413#_c_1218_n 0.00465771f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_797 N_A_1150_159#_c_1103_n N_A_986_413#_c_1218_n 0.0132603f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_798 N_A_1150_159#_c_1106_n N_A_986_413#_c_1218_n 0.00145117f $X=7.36 $Y=1.21
+ $X2=0 $Y2=0
cc_799 N_A_1150_159#_c_1107_n N_A_986_413#_c_1218_n 2.46982e-19 $X=6.07 $Y=0.93
+ $X2=0 $Y2=0
cc_800 N_A_1150_159#_c_1108_n N_A_986_413#_c_1218_n 0.0049948f $X=5.96 $Y=0.93
+ $X2=0 $Y2=0
cc_801 N_A_1150_159#_M1001_g N_A_986_413#_c_1219_n 0.0173823f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_802 N_A_1150_159#_c_1103_n N_A_986_413#_c_1219_n 0.00455719f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_803 N_A_1150_159#_c_1108_n N_A_986_413#_c_1219_n 5.95332e-19 $X=5.96 $Y=0.93
+ $X2=0 $Y2=0
cc_804 N_A_1150_159#_c_1102_n N_A_986_413#_c_1220_n 0.00149495f $X=7.362
+ $Y=1.375 $X2=0 $Y2=0
cc_805 N_A_1150_159#_c_1103_n N_A_986_413#_c_1220_n 0.00339078f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_806 N_A_1150_159#_c_1113_n N_A_986_413#_c_1220_n 0.0056425f $X=6.695 $Y=1.88
+ $X2=0 $Y2=0
cc_807 N_A_1150_159#_M1001_g N_A_986_413#_c_1230_n 0.00989606f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_808 N_A_1150_159#_M1033_g N_A_986_413#_c_1236_n 0.00266694f $X=5.96 $Y=0.445
+ $X2=0 $Y2=0
cc_809 N_A_1150_159#_M1033_g N_A_986_413#_c_1221_n 0.00424924f $X=5.96 $Y=0.445
+ $X2=0 $Y2=0
cc_810 N_A_1150_159#_c_1107_n N_A_986_413#_c_1221_n 0.0222086f $X=6.07 $Y=0.93
+ $X2=0 $Y2=0
cc_811 N_A_1150_159#_c_1108_n N_A_986_413#_c_1221_n 0.00620582f $X=5.96 $Y=0.93
+ $X2=0 $Y2=0
cc_812 N_A_1150_159#_M1001_g N_A_986_413#_c_1226_n 0.0163963f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_813 N_A_1150_159#_c_1113_n N_A_986_413#_c_1226_n 0.00686804f $X=6.695 $Y=1.88
+ $X2=0 $Y2=0
cc_814 N_A_1150_159#_M1001_g N_A_986_413#_c_1222_n 0.0131936f $X=5.825 $Y=2.275
+ $X2=0 $Y2=0
cc_815 N_A_1150_159#_c_1103_n N_A_986_413#_c_1222_n 0.0417632f $X=6.53 $Y=0.915
+ $X2=0 $Y2=0
cc_816 N_A_1150_159#_c_1107_n N_A_986_413#_c_1222_n 0.0114411f $X=6.07 $Y=0.93
+ $X2=0 $Y2=0
cc_817 N_A_1150_159#_c_1108_n N_A_986_413#_c_1222_n 0.00198791f $X=5.96 $Y=0.93
+ $X2=0 $Y2=0
cc_818 N_A_1150_159#_M1023_g N_A_1591_413#_c_1339_n 5.6946e-19 $X=7.425 $Y=2.275
+ $X2=0 $Y2=0
cc_819 N_A_1150_159#_M1011_g N_A_1591_413#_c_1342_n 6.23163e-19 $X=7.495
+ $Y=0.445 $X2=0 $Y2=0
cc_820 N_A_1150_159#_M1001_g N_VPWR_c_1436_n 0.00644429f $X=5.825 $Y=2.275 $X2=0
+ $Y2=0
cc_821 N_A_1150_159#_c_1113_n N_VPWR_c_1436_n 0.0249957f $X=6.695 $Y=1.88 $X2=0
+ $Y2=0
cc_822 N_A_1150_159#_c_1113_n N_VPWR_c_1437_n 0.0210382f $X=6.695 $Y=1.88 $X2=0
+ $Y2=0
cc_823 N_A_1150_159#_M1023_g N_VPWR_c_1438_n 0.0123787f $X=7.425 $Y=2.275 $X2=0
+ $Y2=0
cc_824 N_A_1150_159#_c_1113_n N_VPWR_c_1438_n 0.0256005f $X=6.695 $Y=1.88 $X2=0
+ $Y2=0
cc_825 N_A_1150_159#_M1023_g N_VPWR_c_1443_n 0.00544582f $X=7.425 $Y=2.275 $X2=0
+ $Y2=0
cc_826 N_A_1150_159#_M1001_g N_VPWR_c_1449_n 0.00375838f $X=5.825 $Y=2.275 $X2=0
+ $Y2=0
cc_827 N_A_1150_159#_M1014_d N_VPWR_c_1432_n 0.00172424f $X=6.56 $Y=1.735 $X2=0
+ $Y2=0
cc_828 N_A_1150_159#_M1001_g N_VPWR_c_1432_n 0.0060313f $X=5.825 $Y=2.275 $X2=0
+ $Y2=0
cc_829 N_A_1150_159#_M1023_g N_VPWR_c_1432_n 0.0052001f $X=7.425 $Y=2.275 $X2=0
+ $Y2=0
cc_830 N_A_1150_159#_c_1113_n N_VPWR_c_1432_n 0.00592003f $X=6.695 $Y=1.88 $X2=0
+ $Y2=0
cc_831 N_A_1150_159#_c_1103_n N_VGND_M1033_d 0.00294965f $X=6.53 $Y=0.915 $X2=0
+ $Y2=0
cc_832 N_A_1150_159#_M1033_g N_VGND_c_1738_n 0.013797f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_833 N_A_1150_159#_c_1104_n N_VGND_c_1738_n 0.02237f $X=6.765 $Y=0.39 $X2=0
+ $Y2=0
cc_834 N_A_1150_159#_c_1107_n N_VGND_c_1738_n 0.0221165f $X=6.07 $Y=0.93 $X2=0
+ $Y2=0
cc_835 N_A_1150_159#_c_1108_n N_VGND_c_1738_n 4.43315e-19 $X=5.96 $Y=0.93 $X2=0
+ $Y2=0
cc_836 N_A_1150_159#_M1011_g N_VGND_c_1739_n 0.0133742f $X=7.495 $Y=0.445 $X2=0
+ $Y2=0
cc_837 N_A_1150_159#_c_1101_n N_VGND_c_1739_n 0.00332209f $X=7.397 $Y=1.045
+ $X2=0 $Y2=0
cc_838 N_A_1150_159#_c_1104_n N_VGND_c_1739_n 0.0237563f $X=6.765 $Y=0.39 $X2=0
+ $Y2=0
cc_839 N_A_1150_159#_c_1105_n N_VGND_c_1739_n 0.00471991f $X=7.36 $Y=1.21 $X2=0
+ $Y2=0
cc_840 N_A_1150_159#_c_1104_n N_VGND_c_1744_n 0.0261692f $X=6.765 $Y=0.39 $X2=0
+ $Y2=0
cc_841 N_A_1150_159#_M1011_g N_VGND_c_1746_n 0.00505556f $X=7.495 $Y=0.445 $X2=0
+ $Y2=0
cc_842 N_A_1150_159#_M1033_g N_VGND_c_1752_n 0.00232377f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_843 N_A_1150_159#_M1022_d N_VGND_c_1754_n 0.00172424f $X=6.63 $Y=0.235 $X2=0
+ $Y2=0
cc_844 N_A_1150_159#_M1033_g N_VGND_c_1754_n 0.00261449f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_845 N_A_1150_159#_M1011_g N_VGND_c_1754_n 0.00494779f $X=7.495 $Y=0.445 $X2=0
+ $Y2=0
cc_846 N_A_1150_159#_c_1103_n N_VGND_c_1754_n 0.00432725f $X=6.53 $Y=0.915 $X2=0
+ $Y2=0
cc_847 N_A_1150_159#_c_1104_n N_VGND_c_1754_n 0.00714477f $X=6.765 $Y=0.39 $X2=0
+ $Y2=0
cc_848 N_A_1150_159#_c_1107_n N_VGND_c_1754_n 0.00255175f $X=6.07 $Y=0.93 $X2=0
+ $Y2=0
cc_849 N_A_1150_159#_c_1108_n N_VGND_c_1754_n 7.19298e-19 $X=5.96 $Y=0.93 $X2=0
+ $Y2=0
cc_850 N_A_986_413#_M1014_g N_VPWR_c_1436_n 0.0032365f $X=6.485 $Y=2.11 $X2=0
+ $Y2=0
cc_851 N_A_986_413#_c_1219_n N_VPWR_c_1436_n 0.00132475f $X=6.41 $Y=1.41 $X2=0
+ $Y2=0
cc_852 N_A_986_413#_c_1226_n N_VPWR_c_1436_n 0.0209688f $X=5.87 $Y=2.175 $X2=0
+ $Y2=0
cc_853 N_A_986_413#_c_1222_n N_VPWR_c_1436_n 0.0108482f $X=5.87 $Y=1.41 $X2=0
+ $Y2=0
cc_854 N_A_986_413#_M1014_g N_VPWR_c_1437_n 0.00541359f $X=6.485 $Y=2.11 $X2=0
+ $Y2=0
cc_855 N_A_986_413#_M1014_g N_VPWR_c_1438_n 0.00292103f $X=6.485 $Y=2.11 $X2=0
+ $Y2=0
cc_856 N_A_986_413#_c_1230_n N_VPWR_c_1449_n 0.0372444f $X=5.785 $Y=2.275 $X2=0
+ $Y2=0
cc_857 N_A_986_413#_M1009_d N_VPWR_c_1432_n 0.00206096f $X=4.93 $Y=2.065 $X2=0
+ $Y2=0
cc_858 N_A_986_413#_M1014_g N_VPWR_c_1432_n 0.00782689f $X=6.485 $Y=2.11 $X2=0
+ $Y2=0
cc_859 N_A_986_413#_c_1230_n N_VPWR_c_1432_n 0.0160193f $X=5.785 $Y=2.275 $X2=0
+ $Y2=0
cc_860 N_A_986_413#_c_1230_n N_A_299_47#_c_1598_n 0.0075195f $X=5.785 $Y=2.275
+ $X2=0 $Y2=0
cc_861 N_A_986_413#_c_1236_n N_A_299_47#_c_1592_n 0.00423578f $X=5.51 $Y=0.41
+ $X2=0 $Y2=0
cc_862 N_A_986_413#_c_1236_n N_A_299_47#_c_1594_n 0.00697085f $X=5.51 $Y=0.41
+ $X2=0 $Y2=0
cc_863 N_A_986_413#_c_1230_n A_1077_413# 0.00553919f $X=5.785 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_864 N_A_986_413#_c_1217_n N_VGND_c_1738_n 0.00570804f $X=6.52 $Y=0.95 $X2=0
+ $Y2=0
cc_865 N_A_986_413#_c_1236_n N_VGND_c_1738_n 0.0181194f $X=5.51 $Y=0.41 $X2=0
+ $Y2=0
cc_866 N_A_986_413#_c_1217_n N_VGND_c_1739_n 0.00214573f $X=6.52 $Y=0.95 $X2=0
+ $Y2=0
cc_867 N_A_986_413#_c_1217_n N_VGND_c_1744_n 0.00435091f $X=6.52 $Y=0.95 $X2=0
+ $Y2=0
cc_868 N_A_986_413#_c_1236_n N_VGND_c_1752_n 0.0393557f $X=5.51 $Y=0.41 $X2=0
+ $Y2=0
cc_869 N_A_986_413#_M1006_d N_VGND_c_1754_n 0.00190253f $X=5.065 $Y=0.235 $X2=0
+ $Y2=0
cc_870 N_A_986_413#_c_1217_n N_VGND_c_1754_n 0.00708984f $X=6.52 $Y=0.95 $X2=0
+ $Y2=0
cc_871 N_A_986_413#_c_1236_n N_VGND_c_1754_n 0.0114791f $X=5.51 $Y=0.41 $X2=0
+ $Y2=0
cc_872 N_A_986_413#_c_1236_n A_1101_47# 0.00436463f $X=5.51 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_873 N_A_986_413#_c_1221_n A_1101_47# 0.00105811f $X=5.595 $Y=1.315 $X2=-0.19
+ $Y2=-0.24
cc_874 N_A_1591_413#_c_1339_n N_VPWR_c_1438_n 0.00551479f $X=8.64 $Y=2.26 $X2=0
+ $Y2=0
cc_875 N_A_1591_413#_M1027_g N_VPWR_c_1439_n 0.00188178f $X=9.925 $Y=2.165 $X2=0
+ $Y2=0
cc_876 N_A_1591_413#_M1027_g N_VPWR_c_1440_n 0.00910498f $X=9.925 $Y=2.165 $X2=0
+ $Y2=0
cc_877 N_A_1591_413#_c_1323_n N_VPWR_c_1440_n 0.00466622f $X=10.335 $Y=1.16
+ $X2=0 $Y2=0
cc_878 N_A_1591_413#_M1005_g N_VPWR_c_1440_n 0.00310362f $X=10.41 $Y=1.985 $X2=0
+ $Y2=0
cc_879 N_A_1591_413#_c_1339_n N_VPWR_c_1443_n 0.0295685f $X=8.64 $Y=2.26 $X2=0
+ $Y2=0
cc_880 N_A_1591_413#_M1027_g N_VPWR_c_1445_n 0.00541359f $X=9.925 $Y=2.165 $X2=0
+ $Y2=0
cc_881 N_A_1591_413#_M1005_g N_VPWR_c_1450_n 0.00557712f $X=10.41 $Y=1.985 $X2=0
+ $Y2=0
cc_882 N_A_1591_413#_M1030_d N_VPWR_c_1432_n 0.00215743f $X=7.955 $Y=2.065 $X2=0
+ $Y2=0
cc_883 N_A_1591_413#_M1027_g N_VPWR_c_1432_n 0.0110723f $X=9.925 $Y=2.165 $X2=0
+ $Y2=0
cc_884 N_A_1591_413#_M1005_g N_VPWR_c_1432_n 0.0110874f $X=10.41 $Y=1.985 $X2=0
+ $Y2=0
cc_885 N_A_1591_413#_c_1339_n N_VPWR_c_1432_n 0.0280716f $X=8.64 $Y=2.26 $X2=0
+ $Y2=0
cc_886 N_A_1591_413#_c_1339_n A_1675_413# 0.00905112f $X=8.64 $Y=2.26 $X2=-0.19
+ $Y2=-0.24
cc_887 N_A_1591_413#_c_1337_n A_1675_413# 0.00123507f $X=8.725 $Y=2.165
+ $X2=-0.19 $Y2=-0.24
cc_888 N_A_1591_413#_M1012_g N_Q_c_1718_n 4.27936e-19 $X=9.925 $Y=0.445 $X2=0
+ $Y2=0
cc_889 N_A_1591_413#_M1027_g N_Q_c_1718_n 6.50973e-19 $X=9.925 $Y=2.165 $X2=0
+ $Y2=0
cc_890 N_A_1591_413#_c_1324_n N_Q_c_1718_n 0.00994181f $X=10.41 $Y=0.995 $X2=0
+ $Y2=0
cc_891 N_A_1591_413#_M1005_g N_Q_c_1718_n 0.0153574f $X=10.41 $Y=1.985 $X2=0
+ $Y2=0
cc_892 N_A_1591_413#_c_1327_n N_Q_c_1718_n 0.0164431f $X=10.41 $Y=1.16 $X2=0
+ $Y2=0
cc_893 N_A_1591_413#_c_1342_n N_VGND_c_1739_n 0.00574753f $X=8.64 $Y=0.432 $X2=0
+ $Y2=0
cc_894 N_A_1591_413#_M1012_g N_VGND_c_1740_n 0.00357154f $X=9.925 $Y=0.445 $X2=0
+ $Y2=0
cc_895 N_A_1591_413#_c_1325_n N_VGND_c_1740_n 0.00151274f $X=9.85 $Y=1.16 $X2=0
+ $Y2=0
cc_896 N_A_1591_413#_c_1342_n N_VGND_c_1740_n 0.0129405f $X=8.64 $Y=0.432 $X2=0
+ $Y2=0
cc_897 N_A_1591_413#_c_1328_n N_VGND_c_1740_n 0.00448678f $X=8.725 $Y=0.995
+ $X2=0 $Y2=0
cc_898 N_A_1591_413#_c_1329_n N_VGND_c_1740_n 0.00691913f $X=9.425 $Y=1.16 $X2=0
+ $Y2=0
cc_899 N_A_1591_413#_M1012_g N_VGND_c_1741_n 0.0069333f $X=9.925 $Y=0.445 $X2=0
+ $Y2=0
cc_900 N_A_1591_413#_c_1323_n N_VGND_c_1741_n 0.00495621f $X=10.335 $Y=1.16
+ $X2=0 $Y2=0
cc_901 N_A_1591_413#_c_1324_n N_VGND_c_1741_n 0.00306265f $X=10.41 $Y=0.995
+ $X2=0 $Y2=0
cc_902 N_A_1591_413#_c_1342_n N_VGND_c_1746_n 0.0312214f $X=8.64 $Y=0.432 $X2=0
+ $Y2=0
cc_903 N_A_1591_413#_M1012_g N_VGND_c_1748_n 0.00543148f $X=9.925 $Y=0.445 $X2=0
+ $Y2=0
cc_904 N_A_1591_413#_c_1324_n N_VGND_c_1753_n 0.00557839f $X=10.41 $Y=0.995
+ $X2=0 $Y2=0
cc_905 N_A_1591_413#_M1003_d N_VGND_c_1754_n 0.00256476f $X=8.055 $Y=0.235 $X2=0
+ $Y2=0
cc_906 N_A_1591_413#_M1012_g N_VGND_c_1754_n 0.00952759f $X=9.925 $Y=0.445 $X2=0
+ $Y2=0
cc_907 N_A_1591_413#_c_1324_n N_VGND_c_1754_n 0.0110878f $X=10.41 $Y=0.995 $X2=0
+ $Y2=0
cc_908 N_A_1591_413#_c_1342_n N_VGND_c_1754_n 0.0125713f $X=8.64 $Y=0.432 $X2=0
+ $Y2=0
cc_909 N_A_1591_413#_c_1342_n A_1717_47# 0.00443949f $X=8.64 $Y=0.432 $X2=-0.19
+ $Y2=-0.24
cc_910 N_A_1591_413#_c_1328_n A_1717_47# 0.00147825f $X=8.725 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_911 N_VPWR_c_1432_n N_A_299_47#_M1021_s 0.00172424f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_912 N_VPWR_c_1432_n N_A_299_47#_M1026_d 0.0063859f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_913 N_VPWR_c_1434_n N_A_299_47#_c_1596_n 0.0192069f $X=2.4 $Y=2 $X2=0 $Y2=0
cc_914 N_VPWR_c_1441_n N_A_299_47#_c_1596_n 0.0280365f $X=2.235 $Y=2.72 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1432_n N_A_299_47#_c_1596_n 0.00771147f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1435_n N_A_299_47#_c_1598_n 0.00729213f $X=3.35 $Y=1.99 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1449_n N_A_299_47#_c_1598_n 0.0219939f $X=6.125 $Y=2.72 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1432_n N_A_299_47#_c_1598_n 0.00669153f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1432_n A_381_369# 0.00302076f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_920 N_VPWR_c_1432_n A_729_369# 0.00517845f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_921 N_VPWR_c_1432_n A_1077_413# 0.00247765f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_922 N_VPWR_c_1432_n A_1500_413# 0.0042834f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_923 N_VPWR_c_1432_n A_1675_413# 0.00357865f $X=10.81 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_924 N_VPWR_c_1432_n N_Q_M1005_d 0.00228626f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_925 N_VPWR_c_1440_n N_Q_c_1718_n 0.0365895f $X=10.2 $Y=1.63 $X2=0 $Y2=0
cc_926 N_VPWR_c_1450_n N_Q_c_1718_n 0.0163462f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_927 N_VPWR_c_1432_n N_Q_c_1718_n 0.0121893f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_928 N_VPWR_c_1440_n N_VGND_c_1741_n 0.00976036f $X=10.2 $Y=1.63 $X2=0 $Y2=0
cc_929 N_A_299_47#_c_1593_n N_VGND_M1004_d 0.00213973f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_930 N_A_299_47#_c_1595_n N_VGND_c_1735_n 0.00316681f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_931 N_A_299_47#_c_1593_n N_VGND_c_1736_n 0.0145222f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_932 N_A_299_47#_c_1595_n N_VGND_c_1736_n 0.0070895f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_933 N_A_299_47#_c_1592_n N_VGND_c_1737_n 5.24197e-19 $X=4.27 $Y=0.51 $X2=0
+ $Y2=0
cc_934 N_A_299_47#_c_1593_n N_VGND_c_1737_n 0.0213503f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_935 N_A_299_47#_c_1594_n N_VGND_c_1737_n 0.0056261f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_936 N_A_299_47#_c_1591_n N_VGND_c_1742_n 6.17783e-19 $X=1.585 $Y=0.51 $X2=0
+ $Y2=0
cc_937 N_A_299_47#_c_1593_n N_VGND_c_1742_n 0.00229575f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_938 N_A_299_47#_c_1595_n N_VGND_c_1742_n 0.0264163f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_939 N_A_299_47#_c_1593_n N_VGND_c_1751_n 0.00219701f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_940 N_A_299_47#_c_1593_n N_VGND_c_1752_n 0.00288773f $X=4.125 $Y=0.51 $X2=0
+ $Y2=0
cc_941 N_A_299_47#_c_1594_n N_VGND_c_1752_n 0.0168081f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_942 N_A_299_47#_M1002_s N_VGND_c_1754_n 0.00110044f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_943 N_A_299_47#_M1032_d N_VGND_c_1754_n 0.00786092f $X=4.155 $Y=0.235 $X2=0
+ $Y2=0
cc_944 N_A_299_47#_c_1591_n N_VGND_c_1754_n 0.305313f $X=1.585 $Y=0.51 $X2=0
+ $Y2=0
cc_945 N_A_299_47#_c_1594_n N_VGND_c_1754_n 0.00257571f $X=4.29 $Y=0.445 $X2=0
+ $Y2=0
cc_946 N_A_299_47#_c_1595_n N_VGND_c_1754_n 0.00373095f $X=1.62 $Y=0.415 $X2=0
+ $Y2=0
cc_947 N_A_299_47#_c_1593_n A_381_47# 0.00879585f $X=4.125 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_948 N_A_299_47#_c_1593_n A_729_47# 0.00632255f $X=4.125 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_949 N_Q_c_1718_n N_VGND_c_1741_n 0.022497f $X=10.63 $Y=0.395 $X2=0 $Y2=0
cc_950 N_Q_c_1718_n N_VGND_c_1753_n 0.0159484f $X=10.63 $Y=0.395 $X2=0 $Y2=0
cc_951 N_Q_M1008_d N_VGND_c_1754_n 0.00229159f $X=10.485 $Y=0.235 $X2=0 $Y2=0
cc_952 N_Q_c_1718_n N_VGND_c_1754_n 0.0121559f $X=10.63 $Y=0.395 $X2=0 $Y2=0
cc_953 N_VGND_c_1754_n A_381_47# 0.00172536f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_954 N_VGND_c_1754_n A_729_47# 0.0025277f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_955 N_VGND_c_1754_n A_1101_47# 0.00379452f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_956 N_VGND_c_1754_n A_1514_47# 0.00481883f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24
cc_957 N_VGND_c_1754_n A_1717_47# 0.00296047f $X=10.81 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a221oi_2.spice
* Created: Thu Aug 27 14:02:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a221oi_2.spice.pex"
.subckt sky130_fd_sc_hd__a221oi_2  VNB VPB C1 B2 B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_C1_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1755 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1001_d N_C1_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1008 N_A_383_47#_M1008_d N_B2_M1008_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1013 N_A_383_47#_M1008_d N_B1_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1014 N_A_383_47#_M1014_d N_B1_M1014_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1019 N_A_383_47#_M1014_d N_B2_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75002.8
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1015 N_A_735_47#_M1015_d N_A2_M1015_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=5.532 M=1 R=4.33333 SA=75003.3
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1009 N_A_735_47#_M1015_d N_A1_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1012 N_A_735_47#_M1012_d N_A1_M1012_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_735_47#_M1012_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_27_297#_M1000_d N_C1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.27 AS=0.135 PD=2.54 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1004 N_A_27_297#_M1004_d N_C1_M1004_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_A_301_297#_M1002_d N_B2_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_297#_M1002_s N_B1_M1003_g N_A_301_297#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1007 N_A_27_297#_M1007_d N_B1_M1007_g N_A_301_297#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1011 N_A_301_297#_M1011_d N_B2_M1011_g N_A_27_297#_M1007_d VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.135 PD=1.35 PS=1.27 NRD=6.8753 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75002 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_301_297#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75001.9
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1005_d N_A1_M1010_g N_A_301_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_301_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1017_d N_A2_M1006_g N_A_301_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.285 PD=1.27 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_45 VNB 0 1.67842e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__a221oi_2.spice.SKY130_FD_SC_HD__A221OI_2.pxi"
*
.ends
*
*

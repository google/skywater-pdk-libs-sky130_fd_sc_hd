* File: sky130_fd_sc_hd__o31ai_1.spice
* Created: Thu Aug 27 14:40:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o31ai_1.pex.spice"
.subckt sky130_fd_sc_hd__o31ai_1  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1007 N_A_109_47#_M1007_d N_A1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_109_47#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1003 N_A_109_47#_M1003_d N_A3_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.08775 PD=1.26 PS=0.92 NRD=1.836 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_109_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.221 AS=0.19825 PD=1.98 PS=1.26 NRD=10.152 NRS=59.076 M=1 R=4.33333
+ SA=75001.8 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 A_109_297# N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1001 A_193_297# N_A2_M1001_g A_109_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A3_M1000_g A_193_297# VPB PHIGHVT L=0.15 W=1 AD=0.3925
+ AS=0.135 PD=1.785 PS=1.27 NRD=99.4653 NRS=15.7403 M=1 R=6.66667 SA=75001
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1 AD=0.3
+ AS=0.3925 PD=2.6 PS=1.785 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
*
.include "sky130_fd_sc_hd__o31ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nand4_4.pxi.spice
* Created: Tue Sep  1 19:16:51 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4_4%D N_D_M1009_g N_D_M1002_g N_D_M1014_g N_D_M1003_g
+ N_D_M1017_g N_D_M1018_g N_D_c_128_n N_D_M1030_g N_D_M1027_g D D D D
+ PM_SKY130_FD_SC_HD__NAND4_4%D
x_PM_SKY130_FD_SC_HD__NAND4_4%C N_C_M1015_g N_C_M1000_g N_C_M1020_g N_C_M1004_g
+ N_C_M1025_g N_C_M1022_g N_C_M1026_g N_C_M1028_g C C C C N_C_c_212_n
+ PM_SKY130_FD_SC_HD__NAND4_4%C
x_PM_SKY130_FD_SC_HD__NAND4_4%B N_B_M1007_g N_B_M1001_g N_B_M1010_g N_B_M1005_g
+ N_B_M1016_g N_B_M1008_g N_B_M1021_g N_B_M1029_g B B B B N_B_c_292_n
+ N_B_c_293_n PM_SKY130_FD_SC_HD__NAND4_4%B
x_PM_SKY130_FD_SC_HD__NAND4_4%A N_A_M1011_g N_A_M1006_g N_A_M1013_g N_A_M1012_g
+ N_A_M1023_g N_A_M1019_g N_A_M1024_g N_A_M1031_g A A A N_A_c_371_n
+ PM_SKY130_FD_SC_HD__NAND4_4%A
x_PM_SKY130_FD_SC_HD__NAND4_4%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1027_s
+ N_VPWR_M1004_s N_VPWR_M1028_s N_VPWR_M1005_s N_VPWR_M1029_s N_VPWR_M1012_s
+ N_VPWR_M1031_s N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n
+ N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n
+ N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n
+ N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n VPWR N_VPWR_c_466_n
+ N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_443_n
+ PM_SKY130_FD_SC_HD__NAND4_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND4_4%Y N_Y_M1011_d N_Y_M1023_d N_Y_M1002_d N_Y_M1018_d
+ N_Y_M1000_d N_Y_M1022_d N_Y_M1001_d N_Y_M1008_d N_Y_M1006_d N_Y_M1019_d
+ N_Y_c_569_n N_Y_c_589_n N_Y_c_570_n N_Y_c_596_n N_Y_c_571_n N_Y_c_601_n
+ N_Y_c_572_n N_Y_c_616_n N_Y_c_573_n N_Y_c_632_n N_Y_c_574_n N_Y_c_639_n
+ N_Y_c_575_n N_Y_c_643_n N_Y_c_659_n N_Y_c_567_n N_Y_c_576_n N_Y_c_577_n
+ N_Y_c_673_n N_Y_c_578_n N_Y_c_579_n N_Y_c_580_n N_Y_c_581_n N_Y_c_582_n
+ N_Y_c_583_n Y PM_SKY130_FD_SC_HD__NAND4_4%Y
x_PM_SKY130_FD_SC_HD__NAND4_4%A_27_47# N_A_27_47#_M1009_d N_A_27_47#_M1014_d
+ N_A_27_47#_M1030_d N_A_27_47#_M1020_s N_A_27_47#_M1026_s N_A_27_47#_c_739_n
+ N_A_27_47#_c_740_n N_A_27_47#_c_741_n N_A_27_47#_c_773_p N_A_27_47#_c_742_n
+ N_A_27_47#_c_776_p N_A_27_47#_c_743_n N_A_27_47#_c_744_n
+ PM_SKY130_FD_SC_HD__NAND4_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4_4%VGND N_VGND_M1009_s N_VGND_M1017_s N_VGND_c_796_n
+ N_VGND_c_797_n VGND N_VGND_c_798_n N_VGND_c_799_n N_VGND_c_800_n
+ N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n PM_SKY130_FD_SC_HD__NAND4_4%VGND
x_PM_SKY130_FD_SC_HD__NAND4_4%A_445_47# N_A_445_47#_M1015_d N_A_445_47#_M1025_d
+ N_A_445_47#_M1007_d N_A_445_47#_M1016_d N_A_445_47#_c_887_n
+ PM_SKY130_FD_SC_HD__NAND4_4%A_445_47#
x_PM_SKY130_FD_SC_HD__NAND4_4%A_803_47# N_A_803_47#_M1007_s N_A_803_47#_M1010_s
+ N_A_803_47#_M1021_s N_A_803_47#_M1013_s N_A_803_47#_M1024_s
+ N_A_803_47#_c_920_n N_A_803_47#_c_921_n N_A_803_47#_c_930_n
+ N_A_803_47#_c_922_n N_A_803_47#_c_923_n N_A_803_47#_c_959_n
+ PM_SKY130_FD_SC_HD__NAND4_4%A_803_47#
cc_1 VNB N_D_M1009_g 0.0228678f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_D_M1014_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_3 VNB N_D_M1003_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_4 VNB N_D_M1017_g 0.0170779f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_5 VNB N_D_M1018_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_6 VNB N_D_c_128_n 0.0851909f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.025
cc_7 VNB N_D_M1030_g 0.0173425f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_D_M1027_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB D 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_10 VNB N_C_M1015_g 0.0176998f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_11 VNB N_C_M1000_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_12 VNB N_C_M1020_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_13 VNB N_C_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_14 VNB N_C_M1025_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_15 VNB N_C_M1022_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_16 VNB N_C_M1026_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_17 VNB N_C_M1028_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_18 VNB C 0.00607228f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_19 VNB N_C_c_212_n 0.0626315f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_20 VNB N_B_M1007_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_B_M1001_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_22 VNB N_B_M1010_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_23 VNB N_B_M1005_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_24 VNB N_B_M1016_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_25 VNB N_B_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_26 VNB N_B_M1021_g 0.0182949f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_27 VNB N_B_M1029_g 4.84968e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_28 VNB B 0.00341134f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_29 VNB N_B_c_292_n 0.0304355f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_30 VNB N_B_c_293_n 0.0588674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_M1011_g 0.0177686f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_32 VNB N_A_M1006_g 4.4822e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_33 VNB N_A_M1013_g 0.0172592f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_34 VNB N_A_M1012_g 4.48029e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_35 VNB N_A_M1023_g 0.0172855f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_36 VNB N_A_M1019_g 4.50014e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_37 VNB N_A_M1024_g 0.0229701f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_38 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_39 VNB N_A_c_371_n 0.0862653f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_40 VNB N_VPWR_c_443_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_567_n 0.00600951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB Y 0.00122711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_739_n 0.015377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_27_47#_c_740_n 0.0029408f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_45 VNB N_A_27_47#_c_741_n 0.0122649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_c_742_n 0.0059349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_c_743_n 0.00271098f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_48 VNB N_A_27_47#_c_744_n 0.00127314f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_49 VNB N_VGND_c_796_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.025
cc_50 VNB N_VGND_c_797_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.295
cc_51 VNB N_VGND_c_798_n 0.0143703f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.025
cc_52 VNB N_VGND_c_799_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_53 VNB N_VGND_c_800_n 0.139841f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.295
cc_54 VNB N_VGND_c_801_n 0.374339f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_55 VNB N_VGND_c_802_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_56 VNB N_VGND_c_803_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_57 VNB N_A_445_47#_c_887_n 0.0269328f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.295
cc_58 VNB N_A_803_47#_c_920_n 0.00263528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_803_47#_c_921_n 0.00294889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_803_47#_c_922_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_61 VNB N_A_803_47#_c_923_n 0.0176798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VPB N_D_M1002_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_63 VPB N_D_M1003_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_64 VPB N_D_M1018_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_65 VPB N_D_c_128_n 0.00817555f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.025
cc_66 VPB N_D_M1027_g 0.0194869f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_67 VPB N_C_M1000_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_68 VPB N_C_M1004_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_69 VPB N_C_M1022_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_70 VPB N_C_M1028_g 0.026721f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_71 VPB N_B_M1001_g 0.026721f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_72 VPB N_B_M1005_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_73 VPB N_B_M1008_g 0.0191843f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_74 VPB N_B_M1029_g 0.0201549f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_75 VPB N_A_M1006_g 0.0195915f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_76 VPB N_A_M1012_g 0.0191504f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_77 VPB N_A_M1019_g 0.0191642f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_78 VPB N_A_M1031_g 0.0263683f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_79 VPB N_A_c_371_n 0.00805825f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_80 VPB N_VPWR_c_444_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_445_n 0.0458771f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_82 VPB N_VPWR_c_446_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.53 $Y2=1.105
cc_83 VPB N_VPWR_c_447_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_448_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_85 VPB N_VPWR_c_449_n 0.00645473f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_86 VPB N_VPWR_c_450_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_451_n 0.00474148f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_88 VPB N_VPWR_c_452_n 0.0187412f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.175
cc_89 VPB N_VPWR_c_453_n 0.00410835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_454_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_455_n 0.0464356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_456_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_457_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_458_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_459_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_460_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_461_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_462_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_463_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_464_n 0.0190595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_465_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_466_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_467_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_468_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_469_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_443_n 0.0430679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_Y_c_569_n 0.00223815f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_108 VPB N_Y_c_570_n 0.00219943f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_109 VPB N_Y_c_571_n 0.0035845f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_110 VPB N_Y_c_572_n 0.00219943f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.16
cc_111 VPB N_Y_c_573_n 0.00857646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_Y_c_574_n 0.00219943f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.175
cc_113 VPB N_Y_c_575_n 0.00828681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_Y_c_576_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_Y_c_577_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_Y_c_578_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_Y_c_579_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_580_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_581_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_Y_c_582_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_Y_c_583_n 0.00162617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB Y 0.00132223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 N_D_M1030_g N_C_M1015_g 0.0233915f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_124 N_D_M1027_g N_C_M1000_g 0.0233915f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_125 N_D_c_128_n C 0.00184043f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_126 D C 0.0118174f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_127 N_D_c_128_n N_C_c_212_n 0.0233915f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_128 N_D_M1002_g N_VPWR_c_445_n 0.0041053f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_129 N_D_c_128_n N_VPWR_c_445_n 0.00562759f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_130 D N_VPWR_c_445_n 0.0194886f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_131 N_D_M1003_g N_VPWR_c_446_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_132 N_D_M1018_g N_VPWR_c_446_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_133 N_D_M1027_g N_VPWR_c_447_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_134 N_D_M1002_g N_VPWR_c_456_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_135 N_D_M1003_g N_VPWR_c_456_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_136 N_D_M1018_g N_VPWR_c_458_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_137 N_D_M1027_g N_VPWR_c_458_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_138 N_D_M1002_g N_VPWR_c_443_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_139 N_D_M1003_g N_VPWR_c_443_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_140 N_D_M1018_g N_VPWR_c_443_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_D_M1027_g N_VPWR_c_443_n 0.00952874f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_D_M1002_g N_Y_c_569_n 0.00331821f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_143 N_D_M1003_g N_Y_c_569_n 0.00149073f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_144 N_D_c_128_n N_Y_c_569_n 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_145 D N_Y_c_569_n 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_146 N_D_M1002_g N_Y_c_589_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_147 N_D_M1003_g N_Y_c_589_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_148 N_D_M1018_g N_Y_c_589_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_149 N_D_M1003_g N_Y_c_570_n 0.0120357f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_150 N_D_M1018_g N_Y_c_570_n 0.0120357f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_151 N_D_c_128_n N_Y_c_570_n 0.0019951f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_152 D N_Y_c_570_n 0.0366837f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_153 N_D_M1003_g N_Y_c_596_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_154 N_D_M1018_g N_Y_c_596_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_155 N_D_M1027_g N_Y_c_596_n 0.00975139f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_156 N_D_M1027_g N_Y_c_571_n 0.0132678f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_157 D N_Y_c_571_n 0.00101487f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_158 N_D_M1027_g N_Y_c_601_n 6.1949e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_159 N_D_M1018_g N_Y_c_578_n 0.00149073f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_160 N_D_c_128_n N_Y_c_578_n 0.00206439f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_161 N_D_M1027_g N_Y_c_578_n 0.00149073f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_162 D N_Y_c_578_n 0.026643f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_163 N_D_M1009_g N_A_27_47#_c_740_n 0.0133188f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_164 N_D_M1014_g N_A_27_47#_c_740_n 0.0125938f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_165 N_D_c_128_n N_A_27_47#_c_740_n 0.00325533f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_166 D N_A_27_47#_c_740_n 0.0487569f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_167 N_D_c_128_n N_A_27_47#_c_741_n 0.00584307f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_168 D N_A_27_47#_c_741_n 0.0194939f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_169 N_D_M1017_g N_A_27_47#_c_742_n 0.0125286f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_170 N_D_c_128_n N_A_27_47#_c_742_n 0.00207461f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_171 N_D_M1030_g N_A_27_47#_c_742_n 0.0136531f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_172 D N_A_27_47#_c_742_n 0.0376402f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_173 N_D_c_128_n N_A_27_47#_c_744_n 0.00213429f $X=1.73 $Y=1.025 $X2=0 $Y2=0
cc_174 D N_A_27_47#_c_744_n 0.0138109f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_175 N_D_M1009_g N_VGND_c_796_n 0.00856801f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_176 N_D_M1014_g N_VGND_c_796_n 0.00685342f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_177 N_D_M1017_g N_VGND_c_796_n 5.54209e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_178 N_D_M1014_g N_VGND_c_797_n 5.54209e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_179 N_D_M1017_g N_VGND_c_797_n 0.00685342f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_180 N_D_M1030_g N_VGND_c_797_n 0.00803842f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_181 N_D_M1009_g N_VGND_c_798_n 0.00341689f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_182 N_D_M1014_g N_VGND_c_799_n 0.00341689f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_183 N_D_M1017_g N_VGND_c_799_n 0.00341689f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_184 N_D_M1030_g N_VGND_c_800_n 0.00341689f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_185 N_D_M1009_g N_VGND_c_801_n 0.0050171f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_186 N_D_M1014_g N_VGND_c_801_n 0.0040262f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_187 N_D_M1017_g N_VGND_c_801_n 0.0040262f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_188 N_D_M1030_g N_VGND_c_801_n 0.00405445f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_189 C B 0.0121822f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_190 N_C_c_212_n B 8.71733e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_191 C N_B_c_292_n 8.07044e-19 $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_192 N_C_c_212_n N_B_c_292_n 0.00741568f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_193 N_C_M1000_g N_VPWR_c_447_n 0.00146448f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_194 N_C_M1004_g N_VPWR_c_448_n 0.00146448f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_195 N_C_M1022_g N_VPWR_c_448_n 0.00146448f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_196 N_C_M1028_g N_VPWR_c_449_n 0.0033532f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 N_C_M1000_g N_VPWR_c_460_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_198 N_C_M1004_g N_VPWR_c_460_n 0.00541359f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_199 N_C_M1022_g N_VPWR_c_466_n 0.00541359f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_200 N_C_M1028_g N_VPWR_c_466_n 0.00541359f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_201 N_C_M1000_g N_VPWR_c_443_n 0.00952874f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_202 N_C_M1004_g N_VPWR_c_443_n 0.00950154f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_203 N_C_M1022_g N_VPWR_c_443_n 0.00950154f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_204 N_C_M1028_g N_VPWR_c_443_n 0.0108276f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_205 N_C_M1000_g N_Y_c_596_n 6.1949e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_206 N_C_M1000_g N_Y_c_571_n 0.0119784f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_207 C N_Y_c_571_n 0.0149743f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_208 N_C_M1000_g N_Y_c_601_n 0.00975139f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_209 N_C_M1004_g N_Y_c_601_n 0.00975139f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_210 N_C_M1022_g N_Y_c_601_n 6.1949e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_211 N_C_M1004_g N_Y_c_572_n 0.0120357f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_212 N_C_M1022_g N_Y_c_572_n 0.0120357f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_213 C N_Y_c_572_n 0.0366837f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_214 N_C_c_212_n N_Y_c_572_n 0.0019951f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_215 N_C_M1004_g N_Y_c_616_n 6.1949e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_216 N_C_M1022_g N_Y_c_616_n 0.00975139f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_217 N_C_M1028_g N_Y_c_616_n 0.0145598f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_218 N_C_M1028_g N_Y_c_573_n 0.0147646f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_219 C N_Y_c_573_n 0.0126419f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_220 N_C_M1000_g N_Y_c_579_n 0.00149073f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_221 N_C_M1004_g N_Y_c_579_n 0.00149073f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_222 C N_Y_c_579_n 0.026643f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_223 N_C_c_212_n N_Y_c_579_n 0.00206439f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_224 N_C_M1022_g N_Y_c_580_n 0.00149073f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_225 N_C_M1028_g N_Y_c_580_n 0.00149073f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_226 C N_Y_c_580_n 0.026643f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_227 N_C_c_212_n N_Y_c_580_n 0.00206439f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_228 N_C_M1015_g N_A_27_47#_c_742_n 4.48192e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_229 C N_A_27_47#_c_742_n 0.00297817f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_230 N_C_M1015_g N_A_27_47#_c_743_n 0.0123469f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_231 N_C_M1020_g N_A_27_47#_c_743_n 0.00912735f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_232 N_C_M1025_g N_A_27_47#_c_743_n 0.00918728f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_233 N_C_M1026_g N_A_27_47#_c_743_n 0.00918728f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_234 C N_A_27_47#_c_743_n 0.00381697f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_235 N_C_M1015_g N_VGND_c_797_n 0.00128815f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_236 N_C_M1015_g N_VGND_c_800_n 0.00357877f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_237 N_C_M1020_g N_VGND_c_800_n 0.00357877f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_238 N_C_M1025_g N_VGND_c_800_n 0.00357877f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_239 N_C_M1026_g N_VGND_c_800_n 0.00357877f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_240 N_C_M1015_g N_VGND_c_801_n 0.0052923f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_241 N_C_M1020_g N_VGND_c_801_n 0.00522516f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_242 N_C_M1025_g N_VGND_c_801_n 0.00522516f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_243 N_C_M1026_g N_VGND_c_801_n 0.00655123f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_244 N_C_M1015_g N_A_445_47#_c_887_n 0.0036194f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_245 N_C_M1020_g N_A_445_47#_c_887_n 0.0107009f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_246 N_C_M1025_g N_A_445_47#_c_887_n 0.0107009f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_247 N_C_M1026_g N_A_445_47#_c_887_n 0.0138053f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_248 C N_A_445_47#_c_887_n 0.0987339f $X=3.37 $Y=1.105 $X2=0 $Y2=0
cc_249 N_C_c_212_n N_A_445_47#_c_887_n 0.00622382f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B_M1021_g N_A_M1011_g 0.0153812f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B_M1029_g N_A_M1006_g 0.0153812f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_252 B N_A_c_371_n 7.96788e-19 $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_253 N_B_c_293_n N_A_c_371_n 0.0153812f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B_M1001_g N_VPWR_c_449_n 0.0033532f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B_M1005_g N_VPWR_c_450_n 0.00146448f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_256 N_B_M1008_g N_VPWR_c_450_n 0.00268723f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_257 N_B_M1029_g N_VPWR_c_451_n 0.00487512f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_258 N_B_M1001_g N_VPWR_c_462_n 0.00541359f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_259 N_B_M1005_g N_VPWR_c_462_n 0.00541359f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B_M1008_g N_VPWR_c_464_n 0.00541359f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_261 N_B_M1029_g N_VPWR_c_464_n 0.00541359f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_262 N_B_M1001_g N_VPWR_c_443_n 0.0108276f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_263 N_B_M1005_g N_VPWR_c_443_n 0.00950154f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B_M1008_g N_VPWR_c_443_n 0.00950154f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B_M1029_g N_VPWR_c_443_n 0.00975716f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B_M1001_g N_Y_c_573_n 0.0147646f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_267 B N_Y_c_573_n 0.0400987f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_268 N_B_c_292_n N_Y_c_573_n 0.00729564f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B_M1001_g N_Y_c_632_n 0.0145598f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B_M1005_g N_Y_c_632_n 0.00975139f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B_M1008_g N_Y_c_632_n 6.1949e-19 $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B_M1005_g N_Y_c_574_n 0.0120357f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B_M1008_g N_Y_c_574_n 0.0120357f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_274 B N_Y_c_574_n 0.0366837f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_275 N_B_c_293_n N_Y_c_574_n 0.0019951f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B_M1005_g N_Y_c_639_n 6.1949e-19 $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B_M1008_g N_Y_c_639_n 0.00975139f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B_M1029_g N_Y_c_639_n 0.0105476f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B_M1029_g N_Y_c_575_n 0.0161923f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B_M1029_g N_Y_c_643_n 6.30012e-19 $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_281 N_B_M1001_g N_Y_c_581_n 0.00149073f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_282 N_B_M1005_g N_Y_c_581_n 0.00149073f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_283 B N_Y_c_581_n 0.026643f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_284 N_B_c_293_n N_Y_c_581_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B_M1008_g N_Y_c_582_n 0.00149073f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_286 N_B_M1029_g N_Y_c_582_n 0.00149073f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_287 B N_Y_c_582_n 0.026643f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_288 N_B_c_293_n N_Y_c_582_n 0.00206439f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B_M1021_g Y 0.00263367f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_290 B Y 0.00580225f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_291 N_B_M1007_g N_VGND_c_800_n 0.00357877f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_292 N_B_M1010_g N_VGND_c_800_n 0.00357877f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_293 N_B_M1016_g N_VGND_c_800_n 0.00357877f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_294 N_B_M1021_g N_VGND_c_800_n 0.00357877f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_295 N_B_M1007_g N_VGND_c_801_n 0.00655123f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_296 N_B_M1010_g N_VGND_c_801_n 0.00522516f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_297 N_B_M1016_g N_VGND_c_801_n 0.00522516f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_298 N_B_M1021_g N_VGND_c_801_n 0.00539297f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_299 N_B_M1007_g N_A_445_47#_c_887_n 0.0138053f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_300 N_B_M1010_g N_A_445_47#_c_887_n 0.0107009f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_301 N_B_M1016_g N_A_445_47#_c_887_n 0.0107009f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_302 N_B_M1021_g N_A_445_47#_c_887_n 0.00385251f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_303 B N_A_445_47#_c_887_n 0.126473f $X=5.23 $Y=1.105 $X2=0 $Y2=0
cc_304 N_B_c_292_n N_A_445_47#_c_887_n 0.00758649f $X=4.275 $Y=1.16 $X2=0 $Y2=0
cc_305 N_B_c_293_n N_A_445_47#_c_887_n 0.00622382f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_306 N_B_M1007_g N_A_803_47#_c_920_n 0.00918728f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_307 N_B_M1010_g N_A_803_47#_c_920_n 0.00918728f $X=4.77 $Y=0.56 $X2=0 $Y2=0
cc_308 N_B_M1016_g N_A_803_47#_c_920_n 0.00918728f $X=5.19 $Y=0.56 $X2=0 $Y2=0
cc_309 N_B_M1021_g N_A_803_47#_c_920_n 0.0129875f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_310 N_B_M1021_g N_A_803_47#_c_921_n 0.00410771f $X=5.61 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A_M1006_g N_VPWR_c_451_n 0.00488266f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A_M1006_g N_VPWR_c_452_n 0.00541359f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_313 N_A_M1012_g N_VPWR_c_452_n 0.00541359f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A_M1012_g N_VPWR_c_453_n 0.00268723f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A_M1019_g N_VPWR_c_453_n 0.00146448f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_M1031_g N_VPWR_c_455_n 0.00410837f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_317 A N_VPWR_c_455_n 0.0190809f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_318 N_A_c_371_n N_VPWR_c_455_n 0.00550986f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_M1019_g N_VPWR_c_467_n 0.00541359f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_M1031_g N_VPWR_c_467_n 0.00541359f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_M1006_g N_VPWR_c_443_n 0.00973207f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_M1012_g N_VPWR_c_443_n 0.00950154f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_M1019_g N_VPWR_c_443_n 0.00950154f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_324 N_A_M1031_g N_VPWR_c_443_n 0.0104557f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A_M1006_g N_Y_c_639_n 6.38575e-19 $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_M1006_g N_Y_c_575_n 0.0134006f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A_M1006_g N_Y_c_643_n 0.0104002f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_M1012_g N_Y_c_643_n 0.00975139f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_M1019_g N_Y_c_643_n 6.1949e-19 $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_M1011_g N_Y_c_659_n 0.00404754f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A_M1013_g N_Y_c_567_n 0.0110353f $X=6.51 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_M1023_g N_Y_c_567_n 0.0107009f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_333 N_A_M1024_g N_Y_c_567_n 0.00376463f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_334 A N_Y_c_567_n 0.0615297f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_335 N_A_c_371_n N_Y_c_567_n 0.00566081f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_M1012_g N_Y_c_576_n 0.0120357f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_M1019_g N_Y_c_576_n 0.0120357f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_338 A N_Y_c_576_n 0.0366837f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_339 N_A_c_371_n N_Y_c_576_n 0.0019951f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_M1019_g N_Y_c_577_n 0.00149073f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_M1031_g N_Y_c_577_n 0.00331821f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_342 A N_Y_c_577_n 0.026643f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_343 N_A_c_371_n N_Y_c_577_n 0.00206439f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_M1012_g N_Y_c_673_n 6.1949e-19 $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A_M1019_g N_Y_c_673_n 0.00975139f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A_M1031_g N_Y_c_673_n 0.00902485f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A_M1006_g N_Y_c_583_n 0.00281972f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A_M1012_g N_Y_c_583_n 0.00180793f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A_c_371_n N_Y_c_583_n 0.00156621f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A_M1011_g Y 0.0031541f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A_M1006_g Y 0.00395599f $X=6.09 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A_M1013_g Y 0.00255229f $X=6.51 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A_M1012_g Y 0.00319572f $X=6.51 $Y=1.985 $X2=0 $Y2=0
cc_354 A Y 0.0147921f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_355 N_A_c_371_n Y 0.0160797f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A_M1011_g N_VGND_c_800_n 0.00357877f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_M1013_g N_VGND_c_800_n 0.00357877f $X=6.51 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_M1023_g N_VGND_c_800_n 0.00357877f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_M1024_g N_VGND_c_800_n 0.00357877f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_M1011_g N_VGND_c_801_n 0.00539297f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_M1013_g N_VGND_c_801_n 0.00522516f $X=6.51 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_M1023_g N_VGND_c_801_n 0.00522516f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_M1024_g N_VGND_c_801_n 0.00617937f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_M1011_g N_A_803_47#_c_921_n 0.0040054f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_M1011_g N_A_803_47#_c_930_n 0.0121869f $X=6.09 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_M1013_g N_A_803_47#_c_930_n 0.00918728f $X=6.51 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_M1023_g N_A_803_47#_c_930_n 0.00918728f $X=6.93 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_M1024_g N_A_803_47#_c_930_n 0.0108017f $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_369 A N_A_803_47#_c_930_n 0.00362591f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_370 N_A_M1024_g N_A_803_47#_c_923_n 4.62114e-19 $X=7.35 $Y=0.56 $X2=0 $Y2=0
cc_371 A N_A_803_47#_c_923_n 0.0190063f $X=7.5 $Y=1.105 $X2=0 $Y2=0
cc_372 N_A_c_371_n N_A_803_47#_c_923_n 0.00569691f $X=7.35 $Y=1.16 $X2=0 $Y2=0
cc_373 N_VPWR_c_443_n N_Y_M1002_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_443_n N_Y_M1018_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_c_443_n N_Y_M1000_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_443_n N_Y_M1022_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_377 N_VPWR_c_443_n N_Y_M1001_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_443_n N_Y_M1008_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_c_443_n N_Y_M1006_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_443_n N_Y_M1019_d 0.00215201f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_445_n N_Y_c_569_n 0.0108343f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_382 N_VPWR_c_456_n N_Y_c_589_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_443_n N_Y_c_589_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_M1003_s N_Y_c_570_n 0.00167154f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_385 N_VPWR_c_446_n N_Y_c_570_n 0.0129161f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_386 N_VPWR_c_458_n N_Y_c_596_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_443_n N_Y_c_596_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1027_s N_Y_c_571_n 0.00167154f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_447_n N_Y_c_571_n 0.0129161f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_390 N_VPWR_c_460_n N_Y_c_601_n 0.0189039f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_443_n N_Y_c_601_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_M1004_s N_Y_c_572_n 0.00167154f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_393 N_VPWR_c_448_n N_Y_c_572_n 0.0129161f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_394 N_VPWR_c_466_n N_Y_c_616_n 0.0189039f $X=3.535 $Y=2.72 $X2=0 $Y2=0
cc_395 N_VPWR_c_443_n N_Y_c_616_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_M1028_s N_Y_c_573_n 0.0115037f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_397 N_VPWR_c_449_n N_Y_c_573_n 0.0559698f $X=4.14 $Y=2 $X2=0 $Y2=0
cc_398 N_VPWR_c_462_n N_Y_c_632_n 0.0189039f $X=4.895 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_443_n N_Y_c_632_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_M1005_s N_Y_c_574_n 0.00167154f $X=4.845 $Y=1.485 $X2=0 $Y2=0
cc_401 N_VPWR_c_450_n N_Y_c_574_n 0.0129161f $X=4.98 $Y=2 $X2=0 $Y2=0
cc_402 N_VPWR_c_451_n N_Y_c_639_n 0.0402652f $X=5.855 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_464_n N_Y_c_639_n 0.0189039f $X=5.77 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_443_n N_Y_c_639_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1029_s N_Y_c_575_n 0.00368964f $X=5.685 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_c_451_n N_Y_c_575_n 0.0139097f $X=5.855 $Y=2 $X2=0 $Y2=0
cc_407 N_VPWR_c_451_n N_Y_c_643_n 0.0418431f $X=5.855 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_452_n N_Y_c_643_n 0.0189039f $X=6.635 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_443_n N_Y_c_643_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_M1012_s N_Y_c_576_n 0.00167154f $X=6.585 $Y=1.485 $X2=0 $Y2=0
cc_411 N_VPWR_c_453_n N_Y_c_576_n 0.0129161f $X=6.72 $Y=2 $X2=0 $Y2=0
cc_412 N_VPWR_c_455_n N_Y_c_577_n 0.010839f $X=7.56 $Y=1.66 $X2=0 $Y2=0
cc_413 N_VPWR_c_467_n N_Y_c_673_n 0.0189039f $X=7.475 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_443_n N_Y_c_673_n 0.0122217f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_c_445_n N_A_27_47#_c_741_n 5.83538e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_416 N_VPWR_c_455_n N_A_803_47#_c_923_n 7.91944e-19 $X=7.56 $Y=1.66 $X2=0
+ $Y2=0
cc_417 N_Y_c_571_n N_A_27_47#_c_742_n 0.00983243f $X=2.195 $Y=1.555 $X2=0 $Y2=0
cc_418 N_Y_M1011_d N_VGND_c_801_n 0.00216833f $X=6.165 $Y=0.235 $X2=0 $Y2=0
cc_419 N_Y_M1023_d N_VGND_c_801_n 0.00216833f $X=7.005 $Y=0.235 $X2=0 $Y2=0
cc_420 N_Y_c_573_n N_A_445_47#_c_887_n 0.0110045f $X=4.395 $Y=1.555 $X2=0 $Y2=0
cc_421 N_Y_c_567_n N_A_803_47#_M1013_s 0.00162409f $X=7.14 $Y=0.74 $X2=0 $Y2=0
cc_422 N_Y_c_575_n N_A_803_47#_c_921_n 0.00644161f $X=6.11 $Y=1.555 $X2=0 $Y2=0
cc_423 N_Y_c_659_n N_A_803_47#_c_921_n 0.0196757f $X=6.29 $Y=0.78 $X2=0 $Y2=0
cc_424 N_Y_M1011_d N_A_803_47#_c_930_n 0.00304831f $X=6.165 $Y=0.235 $X2=0 $Y2=0
cc_425 N_Y_M1023_d N_A_803_47#_c_930_n 0.0030596f $X=7.005 $Y=0.235 $X2=0 $Y2=0
cc_426 N_Y_c_659_n N_A_803_47#_c_930_n 0.00938106f $X=6.29 $Y=0.78 $X2=0 $Y2=0
cc_427 N_Y_c_567_n N_A_803_47#_c_930_n 0.0513693f $X=7.14 $Y=0.74 $X2=0 $Y2=0
cc_428 N_Y_c_567_n N_A_803_47#_c_923_n 0.01117f $X=7.14 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A_27_47#_c_740_n N_VGND_M1009_s 0.00162029f $X=1.015 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_430 N_A_27_47#_c_742_n N_VGND_M1017_s 0.00162029f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_431 N_A_27_47#_c_740_n N_VGND_c_796_n 0.0164771f $X=1.015 $Y=0.78 $X2=0 $Y2=0
cc_432 N_A_27_47#_c_742_n N_VGND_c_797_n 0.0164771f $X=1.855 $Y=0.78 $X2=0 $Y2=0
cc_433 N_A_27_47#_c_739_n N_VGND_c_798_n 0.0175846f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_740_n N_VGND_c_798_n 0.00237003f $X=1.015 $Y=0.78 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_c_740_n N_VGND_c_799_n 0.00237003f $X=1.015 $Y=0.78 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_773_p N_VGND_c_799_n 0.0113595f $X=1.1 $Y=0.655 $X2=0 $Y2=0
cc_437 N_A_27_47#_c_742_n N_VGND_c_799_n 0.00237003f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_742_n N_VGND_c_800_n 0.00237003f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_776_p N_VGND_c_800_n 0.0114305f $X=2.025 $Y=0.37 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_743_n N_VGND_c_800_n 0.0994545f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_441 N_A_27_47#_M1009_d N_VGND_c_801_n 0.00229009f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_M1014_d N_VGND_c_801_n 0.00254582f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_M1030_d N_VGND_c_801_n 0.00236502f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_M1020_s N_VGND_c_801_n 0.00215227f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1026_s N_VGND_c_801_n 0.00209344f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_739_n N_VGND_c_801_n 0.00973192f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_740_n N_VGND_c_801_n 0.00989142f $X=1.015 $Y=0.78 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_773_p N_VGND_c_801_n 0.0064623f $X=1.1 $Y=0.655 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_742_n N_VGND_c_801_n 0.00989142f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_776_p N_VGND_c_801_n 0.00653924f $X=2.025 $Y=0.37 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_743_n N_VGND_c_801_n 0.063033f $X=3.62 $Y=0.4 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_743_n N_A_445_47#_M1015_d 0.0030596f $X=3.62 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_453 N_A_27_47#_c_743_n N_A_445_47#_M1025_d 0.0030596f $X=3.62 $Y=0.4 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1020_s N_A_445_47#_c_887_n 0.00162409f $X=2.645 $Y=0.235
+ $X2=0 $Y2=0
cc_455 N_A_27_47#_M1026_s N_A_445_47#_c_887_n 0.00312742f $X=3.485 $Y=0.235
+ $X2=0 $Y2=0
cc_456 N_A_27_47#_c_742_n N_A_445_47#_c_887_n 0.0113394f $X=1.855 $Y=0.78 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_743_n N_A_445_47#_c_887_n 0.0842925f $X=3.62 $Y=0.4 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_743_n N_A_803_47#_c_920_n 0.0197363f $X=3.62 $Y=0.4 $X2=0
+ $Y2=0
cc_459 N_VGND_c_801_n N_A_445_47#_M1015_d 0.00216833f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_460 N_VGND_c_801_n N_A_445_47#_M1025_d 0.00216833f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_801_n N_A_445_47#_M1007_d 0.00216833f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_801_n N_A_445_47#_M1016_d 0.00216833f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_800_n N_A_445_47#_c_887_n 0.00342407f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_801_n N_A_445_47#_c_887_n 0.0114501f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_c_801_n N_A_803_47#_M1007_s 0.00209344f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_466 N_VGND_c_801_n N_A_803_47#_M1010_s 0.00215227f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_801_n N_A_803_47#_M1021_s 0.00263396f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_801_n N_A_803_47#_M1013_s 0.00215227f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_801_n N_A_803_47#_M1024_s 0.00209324f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_800_n N_A_803_47#_c_920_n 0.101456f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_801_n N_A_803_47#_c_920_n 0.0642748f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_472 N_VGND_c_800_n N_A_803_47#_c_930_n 0.0847971f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_801_n N_A_803_47#_c_930_n 0.0545231f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_800_n N_A_803_47#_c_922_n 0.0176918f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_801_n N_A_803_47#_c_922_n 0.00980895f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_800_n N_A_803_47#_c_959_n 0.0119155f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_c_801_n N_A_803_47#_c_959_n 0.00653933f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_478 N_A_445_47#_c_887_n N_A_803_47#_M1007_s 0.00312742f $X=5.4 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_479 N_A_445_47#_c_887_n N_A_803_47#_M1010_s 0.00162409f $X=5.4 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A_445_47#_M1007_d N_A_803_47#_c_920_n 0.0030596f $X=4.425 $Y=0.235
+ $X2=0 $Y2=0
cc_481 N_A_445_47#_M1016_d N_A_803_47#_c_920_n 0.0030596f $X=5.265 $Y=0.235
+ $X2=0 $Y2=0
cc_482 N_A_445_47#_c_887_n N_A_803_47#_c_920_n 0.0842925f $X=5.4 $Y=0.74 $X2=0
+ $Y2=0
cc_483 N_A_445_47#_c_887_n N_A_803_47#_c_921_n 0.0168798f $X=5.4 $Y=0.74 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__or4b_1.spice.SKY130_FD_SC_HD__OR4B_1.pxi
* Created: Thu Aug 27 14:44:21 2020
* 
x_PM_SKY130_FD_SC_HD__OR4B_1%D_N N_D_N_M1002_g N_D_N_M1007_g D_N D_N
+ N_D_N_c_76_n PM_SKY130_FD_SC_HD__OR4B_1%D_N
x_PM_SKY130_FD_SC_HD__OR4B_1%A_109_53# N_A_109_53#_M1002_d N_A_109_53#_M1007_d
+ N_A_109_53#_M1005_g N_A_109_53#_M1000_g N_A_109_53#_c_101_n
+ N_A_109_53#_c_105_n N_A_109_53#_c_102_n N_A_109_53#_c_103_n
+ PM_SKY130_FD_SC_HD__OR4B_1%A_109_53#
x_PM_SKY130_FD_SC_HD__OR4B_1%C N_C_M1004_g N_C_M1009_g C C N_C_c_142_n
+ PM_SKY130_FD_SC_HD__OR4B_1%C
x_PM_SKY130_FD_SC_HD__OR4B_1%B N_B_c_180_n N_B_M1010_g N_B_M1003_g N_B_c_178_n
+ N_B_c_179_n B B B B N_B_c_182_n PM_SKY130_FD_SC_HD__OR4B_1%B
x_PM_SKY130_FD_SC_HD__OR4B_1%A N_A_M1006_g N_A_M1011_g A N_A_c_218_n N_A_c_219_n
+ PM_SKY130_FD_SC_HD__OR4B_1%A
x_PM_SKY130_FD_SC_HD__OR4B_1%A_215_297# N_A_215_297#_M1005_d
+ N_A_215_297#_M1003_d N_A_215_297#_M1000_s N_A_215_297#_M1008_g
+ N_A_215_297#_M1001_g N_A_215_297#_c_268_n N_A_215_297#_c_340_p
+ N_A_215_297#_c_259_n N_A_215_297#_c_260_n N_A_215_297#_c_348_p
+ N_A_215_297#_c_261_n N_A_215_297#_c_304_n N_A_215_297#_c_269_n
+ N_A_215_297#_c_270_n N_A_215_297#_c_262_n N_A_215_297#_c_271_n
+ N_A_215_297#_c_263_n N_A_215_297#_c_264_n N_A_215_297#_c_265_n
+ N_A_215_297#_c_266_n PM_SKY130_FD_SC_HD__OR4B_1%A_215_297#
x_PM_SKY130_FD_SC_HD__OR4B_1%VPWR N_VPWR_M1007_s N_VPWR_M1011_d N_VPWR_c_358_n
+ N_VPWR_c_359_n N_VPWR_c_360_n VPWR N_VPWR_c_361_n N_VPWR_c_362_n
+ N_VPWR_c_357_n N_VPWR_c_364_n PM_SKY130_FD_SC_HD__OR4B_1%VPWR
x_PM_SKY130_FD_SC_HD__OR4B_1%X N_X_M1008_d N_X_M1001_d N_X_c_400_n N_X_c_402_n
+ N_X_c_401_n X PM_SKY130_FD_SC_HD__OR4B_1%X
x_PM_SKY130_FD_SC_HD__OR4B_1%VGND N_VGND_M1002_s N_VGND_M1005_s N_VGND_M1004_d
+ N_VGND_M1006_d N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n
+ N_VGND_c_422_n VGND N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ PM_SKY130_FD_SC_HD__OR4B_1%VGND
cc_1 VNB N_D_N_M1002_g 0.0365462f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB D_N 0.0235541f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_N_c_76_n 0.0396061f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_109_53#_M1005_g 0.0324971f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB N_A_109_53#_c_101_n 0.0137682f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_109_53#_c_102_n 0.0124493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_109_53#_c_103_n 0.0351157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_C_M1004_g 0.025648f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_9 VNB C 0.0071247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_C_c_142_n 0.0181144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_M1010_g 0.0178172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_178_n 0.013575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B_c_179_n 0.0105451f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_14 VNB N_A_M1006_g 0.0265609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_15 VNB N_A_c_218_n 0.0203331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_c_219_n 0.00298835f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_17 VNB N_A_215_297#_c_259_n 0.00408712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_215_297#_c_260_n 0.00318069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_215_297#_c_261_n 0.00106516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_297#_c_262_n 0.00206408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_215_297#_c_263_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_297#_c_264_n 0.0234012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_215_297#_c_265_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_297#_c_266_n 0.0197196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_357_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_400_n 0.0137601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_401_n 0.0241563f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_VGND_c_418_n 0.010416f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_29 VNB N_VGND_c_419_n 0.0171418f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_30 VNB N_VGND_c_420_n 0.00617292f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=0.85
cc_31 VNB N_VGND_c_421_n 7.9456e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_422_n 6.33941e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_423_n 0.0164253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_424_n 0.0133917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_425_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_426_n 0.0166241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_427_n 0.217992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_428_n 0.00531134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_429_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_430_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_D_N_M1007_g 0.0293008f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_42 VPB D_N 0.00399928f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_43 VPB N_D_N_c_76_n 0.0102869f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_44 VPB N_A_109_53#_M1000_g 0.023679f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_45 VPB N_A_109_53#_c_105_n 0.0120604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_109_53#_c_102_n 0.0082693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_109_53#_c_103_n 0.00901831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_C_M1009_g 0.0166456f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_49 VPB C 0.00184565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_C_c_142_n 0.00438963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_B_c_180_n 0.0369467f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.475
cc_52 VPB N_B_M1010_g 0.0240989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_B_c_182_n 0.0545817f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_M1011_g 0.0211368f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_55 VPB N_A_c_218_n 0.0040133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_c_219_n 0.0015525f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_57 VPB N_A_215_297#_M1001_g 0.0244726f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_58 VPB N_A_215_297#_c_268_n 0.00562978f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_59 VPB N_A_215_297#_c_269_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_215_297#_c_270_n 0.0074033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_215_297#_c_271_n 0.00130803f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_215_297#_c_264_n 0.00544454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_358_n 0.0114263f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_64 VPB N_VPWR_c_359_n 0.0547557f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_65 VPB N_VPWR_c_360_n 0.0125184f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_66 VPB N_VPWR_c_361_n 0.0590127f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_67 VPB N_VPWR_c_362_n 0.0177135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_357_n 0.0690193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_364_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_X_c_402_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_71 VPB N_X_c_401_n 0.00880472f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_72 VPB X 0.032187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 N_D_N_M1002_g N_A_109_53#_c_101_n 0.00816837f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_74 D_N N_A_109_53#_c_101_n 0.0185539f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_D_N_M1007_g N_A_109_53#_c_105_n 0.00756693f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_76 D_N N_A_109_53#_c_102_n 0.0276279f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_77 N_D_N_c_76_n N_A_109_53#_c_102_n 0.00409125f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_78 D_N N_A_109_53#_c_103_n 2.0259e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_79 N_D_N_c_76_n N_A_109_53#_c_103_n 0.00634274f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_80 N_D_N_M1007_g N_A_215_297#_c_270_n 0.00126316f $X=0.47 $Y=1.695 $X2=0
+ $Y2=0
cc_81 N_D_N_M1007_g N_VPWR_c_359_n 0.0120555f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_82 D_N N_VPWR_c_359_n 0.020736f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_83 N_D_N_c_76_n N_VPWR_c_359_n 0.00200083f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_84 N_D_N_M1007_g N_VPWR_c_361_n 0.00261702f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_85 N_D_N_M1007_g N_VPWR_c_357_n 0.00336774f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_86 N_D_N_M1002_g N_VGND_c_419_n 0.0104139f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_87 D_N N_VGND_c_419_n 0.0268998f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_88 N_D_N_c_76_n N_VGND_c_419_n 0.00122319f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_89 N_D_N_M1002_g N_VGND_c_420_n 0.00259868f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_90 N_D_N_M1002_g N_VGND_c_423_n 0.00442511f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_91 N_D_N_M1002_g N_VGND_c_427_n 0.00889084f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_92 D_N N_VGND_c_427_n 0.00135692f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_93 N_A_109_53#_M1005_g N_C_M1004_g 0.0197432f $X=1.41 $Y=0.475 $X2=0 $Y2=0
cc_94 N_A_109_53#_M1000_g N_C_M1009_g 0.0259588f $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_95 N_A_109_53#_c_102_n C 0.0205853f $X=1.165 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_109_53#_c_103_n C 0.0093658f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_109_53#_c_102_n N_C_c_142_n 2.26856e-19 $X=1.165 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_109_53#_c_103_n N_C_c_142_n 0.0208217f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_109_53#_M1000_g N_B_c_182_n 0.00441071f $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_100 N_A_109_53#_c_105_n N_B_c_182_n 0.0162027f $X=0.68 $Y=1.72 $X2=0 $Y2=0
cc_101 N_A_109_53#_M1000_g N_A_215_297#_c_268_n 0.0118251f $X=1.41 $Y=1.695
+ $X2=0 $Y2=0
cc_102 N_A_109_53#_M1005_g N_A_215_297#_c_260_n 0.00522712f $X=1.41 $Y=0.475
+ $X2=0 $Y2=0
cc_103 N_A_109_53#_M1000_g N_A_215_297#_c_270_n 0.00723013f $X=1.41 $Y=1.695
+ $X2=0 $Y2=0
cc_104 N_A_109_53#_c_105_n N_A_215_297#_c_270_n 0.0313054f $X=0.68 $Y=1.72 $X2=0
+ $Y2=0
cc_105 N_A_109_53#_c_102_n N_A_215_297#_c_270_n 0.0176028f $X=1.165 $Y=1.16
+ $X2=0 $Y2=0
cc_106 N_A_109_53#_c_103_n N_A_215_297#_c_270_n 0.00736963f $X=1.41 $Y=1.16
+ $X2=0 $Y2=0
cc_107 N_A_109_53#_c_105_n N_VPWR_c_359_n 0.014125f $X=0.68 $Y=1.72 $X2=0 $Y2=0
cc_108 N_A_109_53#_c_105_n N_VPWR_c_357_n 0.00106784f $X=0.68 $Y=1.72 $X2=0
+ $Y2=0
cc_109 N_A_109_53#_M1005_g N_VGND_c_420_n 0.0111676f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_110 N_A_109_53#_c_101_n N_VGND_c_420_n 0.0207055f $X=0.68 $Y=0.5 $X2=0 $Y2=0
cc_111 N_A_109_53#_c_102_n N_VGND_c_420_n 0.00902763f $X=1.165 $Y=1.16 $X2=0
+ $Y2=0
cc_112 N_A_109_53#_c_103_n N_VGND_c_420_n 0.00612453f $X=1.41 $Y=1.16 $X2=0
+ $Y2=0
cc_113 N_A_109_53#_M1005_g N_VGND_c_421_n 5.20066e-19 $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_114 N_A_109_53#_c_101_n N_VGND_c_423_n 0.0128191f $X=0.68 $Y=0.5 $X2=0 $Y2=0
cc_115 N_A_109_53#_M1005_g N_VGND_c_424_n 0.00442511f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_116 N_A_109_53#_M1005_g N_VGND_c_427_n 0.0079095f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_117 N_A_109_53#_c_101_n N_VGND_c_427_n 0.00912835f $X=0.68 $Y=0.5 $X2=0 $Y2=0
cc_118 N_C_M1009_g N_B_M1010_g 0.0443586f $X=1.885 $Y=1.695 $X2=0 $Y2=0
cc_119 C N_B_M1010_g 0.0187585f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_120 N_C_c_142_n N_B_M1010_g 0.0213084f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_121 N_C_M1004_g N_B_c_178_n 0.0136769f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_122 N_C_M1004_g N_B_c_179_n 0.0137915f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_123 N_C_M1009_g N_B_c_182_n 0.00439246f $X=1.885 $Y=1.695 $X2=0 $Y2=0
cc_124 C N_A_M1011_g 0.00101963f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_125 C N_A_c_218_n 2.93432e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_126 C N_A_c_219_n 0.0279535f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_127 N_C_M1009_g N_A_215_297#_c_268_n 0.00926379f $X=1.885 $Y=1.695 $X2=0
+ $Y2=0
cc_128 C N_A_215_297#_c_268_n 0.0427505f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_129 N_C_c_142_n N_A_215_297#_c_268_n 3.54678e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_130 N_C_M1004_g N_A_215_297#_c_259_n 0.0109295f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_131 C N_A_215_297#_c_259_n 0.0414766f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_132 N_C_c_142_n N_A_215_297#_c_259_n 0.00187025f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_133 C N_A_215_297#_c_260_n 0.0152593f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_134 N_C_c_142_n N_A_215_297#_c_260_n 9.23324e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_135 N_C_M1009_g N_A_215_297#_c_270_n 9.66796e-19 $X=1.885 $Y=1.695 $X2=0
+ $Y2=0
cc_136 C N_A_215_297#_c_271_n 0.00739975f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_137 C A_297_297# 0.00283158f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_138 C A_392_297# 0.00111992f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_139 N_C_M1004_g N_VGND_c_420_n 5.57841e-19 $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_140 N_C_M1004_g N_VGND_c_421_n 0.00693276f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_141 N_C_M1004_g N_VGND_c_424_n 0.00322006f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_142 N_C_M1004_g N_VGND_c_427_n 0.00396803f $X=1.865 $Y=0.475 $X2=0 $Y2=0
cc_143 N_B_M1010_g N_A_M1006_g 0.00366469f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_144 N_B_c_178_n N_A_M1006_g 0.0187531f $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_145 N_B_M1010_g N_A_M1011_g 0.0271408f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_146 N_B_c_182_n N_A_M1011_g 8.96507e-19 $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_147 N_B_M1010_g N_A_c_218_n 0.0172254f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_148 N_B_M1010_g N_A_c_219_n 0.0020271f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_149 N_B_c_180_n N_A_215_297#_c_268_n 0.0011988f $X=2.25 $Y=2.145 $X2=0 $Y2=0
cc_150 N_B_M1010_g N_A_215_297#_c_268_n 0.0113982f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_151 N_B_c_182_n N_A_215_297#_c_268_n 0.084547f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_152 N_B_c_178_n N_A_215_297#_c_259_n 0.00683722f $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_153 N_B_c_179_n N_A_215_297#_c_259_n 0.00840807f $X=2.267 $Y=0.91 $X2=0 $Y2=0
cc_154 N_B_c_182_n N_A_215_297#_c_270_n 0.0260771f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_155 N_B_M1010_g N_A_215_297#_c_271_n 0.0045878f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_156 N_B_c_182_n N_A_215_297#_c_271_n 0.0136891f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_157 N_B_c_182_n N_VPWR_c_359_n 0.0240471f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_158 N_B_c_180_n N_VPWR_c_360_n 7.25512e-19 $X=2.25 $Y=2.145 $X2=0 $Y2=0
cc_159 N_B_M1010_g N_VPWR_c_360_n 0.00255415f $X=2.25 $Y=1.695 $X2=0 $Y2=0
cc_160 N_B_c_182_n N_VPWR_c_360_n 0.02518f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_161 N_B_c_180_n N_VPWR_c_361_n 0.00735836f $X=2.25 $Y=2.145 $X2=0 $Y2=0
cc_162 N_B_c_182_n N_VPWR_c_361_n 0.103458f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_163 N_B_c_180_n N_VPWR_c_357_n 0.0106117f $X=2.25 $Y=2.145 $X2=0 $Y2=0
cc_164 N_B_c_182_n N_VPWR_c_357_n 0.0748203f $X=2.295 $Y=2.28 $X2=0 $Y2=0
cc_165 N_B_c_178_n N_VGND_c_421_n 0.00679416f $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_166 N_B_c_178_n N_VGND_c_422_n 5.25642e-19 $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_167 N_B_c_178_n N_VGND_c_425_n 0.00322006f $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_168 N_B_c_178_n N_VGND_c_427_n 0.00390029f $X=2.267 $Y=0.76 $X2=0 $Y2=0
cc_169 N_A_M1011_g N_A_215_297#_M1001_g 0.0189405f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_170 N_A_M1011_g N_A_215_297#_c_268_n 2.08355e-19 $X=2.705 $Y=1.695 $X2=0
+ $Y2=0
cc_171 N_A_c_219_n N_A_215_297#_c_268_n 0.00230038f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_M1006_g N_A_215_297#_c_261_n 0.0116406f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_173 N_A_c_218_n N_A_215_297#_c_261_n 0.00220162f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_219_n N_A_215_297#_c_261_n 0.0166868f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_M1011_g N_A_215_297#_c_304_n 0.0112156f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_176 N_A_c_219_n N_A_215_297#_c_304_n 0.00969518f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_M1011_g N_A_215_297#_c_269_n 0.0034529f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_178 N_A_c_218_n N_A_215_297#_c_262_n 5.77159e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_219_n N_A_215_297#_c_262_n 0.0128912f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_M1011_g N_A_215_297#_c_271_n 0.00985088f $X=2.705 $Y=1.695 $X2=0
+ $Y2=0
cc_181 N_A_c_218_n N_A_215_297#_c_271_n 0.00156816f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_219_n N_A_215_297#_c_271_n 0.0112207f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_c_218_n N_A_215_297#_c_263_n 0.00186332f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_c_219_n N_A_215_297#_c_263_n 0.0259797f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_218_n N_A_215_297#_c_264_n 0.0202671f $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_219_n N_A_215_297#_c_264_n 3.58533e-19 $X=2.69 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_M1006_g N_A_215_297#_c_265_n 0.0034529f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_188 N_A_M1006_g N_A_215_297#_c_266_n 0.0172443f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_189 N_A_M1011_g N_VPWR_c_360_n 0.00293484f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_190 N_A_M1011_g N_VPWR_c_361_n 0.00264561f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_191 N_A_M1011_g N_VPWR_c_357_n 0.00333991f $X=2.705 $Y=1.695 $X2=0 $Y2=0
cc_192 N_A_M1006_g N_VGND_c_421_n 5.2354e-19 $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_193 N_A_M1006_g N_VGND_c_422_n 0.00709299f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_194 N_A_M1006_g N_VGND_c_425_n 0.00322006f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_195 N_A_M1006_g N_VGND_c_427_n 0.00390029f $X=2.705 $Y=0.475 $X2=0 $Y2=0
cc_196 N_A_215_297#_c_304_n N_VPWR_M1011_d 0.00526233f $X=2.98 $Y=1.58 $X2=0
+ $Y2=0
cc_197 N_A_215_297#_c_270_n N_VPWR_c_359_n 0.00105998f $X=1.2 $Y=1.685 $X2=0
+ $Y2=0
cc_198 N_A_215_297#_M1001_g N_VPWR_c_360_n 0.00485906f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_215_297#_c_304_n N_VPWR_c_360_n 0.0190361f $X=2.98 $Y=1.58 $X2=0
+ $Y2=0
cc_200 N_A_215_297#_c_271_n N_VPWR_c_360_n 0.00605542f $X=2.575 $Y=1.58 $X2=0
+ $Y2=0
cc_201 N_A_215_297#_c_264_n N_VPWR_c_360_n 2.11345e-19 $X=3.17 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_215_297#_M1001_g N_VPWR_c_362_n 0.00585385f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_215_297#_M1001_g N_VPWR_c_357_n 0.0128443f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_215_297#_c_268_n A_297_297# 0.0021725f $X=2.49 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_205 N_A_215_297#_c_268_n A_392_297# 0.00107627f $X=2.49 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_215_297#_c_268_n A_465_297# 0.00315317f $X=2.49 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_207 N_A_215_297#_c_271_n A_465_297# 0.00424971f $X=2.575 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_208 N_A_215_297#_M1001_g N_X_c_401_n 0.00349311f $X=3.195 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_215_297#_c_261_n N_X_c_401_n 0.0035218f $X=2.98 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_215_297#_c_269_n N_X_c_401_n 0.00841221f $X=3.065 $Y=1.495 $X2=0
+ $Y2=0
cc_211 N_A_215_297#_c_263_n N_X_c_401_n 0.024459f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_215_297#_c_264_n N_X_c_401_n 0.00753248f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_215_297#_c_265_n N_X_c_401_n 0.00836618f $X=3.117 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_215_297#_c_266_n N_X_c_401_n 0.00441003f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_215_297#_c_259_n N_VGND_M1004_d 0.00160115f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_216 N_A_215_297#_c_261_n N_VGND_M1006_d 0.00482895f $X=2.98 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A_215_297#_c_265_n N_VGND_M1006_d 6.98847e-19 $X=3.117 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_215_297#_c_340_p N_VGND_c_420_n 0.0182384f $X=1.65 $Y=0.47 $X2=0
+ $Y2=0
cc_219 N_A_215_297#_c_259_n N_VGND_c_421_n 0.0160613f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_215_297#_c_261_n N_VGND_c_422_n 0.020701f $X=2.98 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_215_297#_c_264_n N_VGND_c_422_n 2.33671e-19 $X=3.17 $Y=1.16 $X2=0
+ $Y2=0
cc_222 N_A_215_297#_c_266_n N_VGND_c_422_n 0.0132447f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_215_297#_c_340_p N_VGND_c_424_n 0.00873683f $X=1.65 $Y=0.47 $X2=0
+ $Y2=0
cc_224 N_A_215_297#_c_259_n N_VGND_c_424_n 0.00237039f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_215_297#_c_259_n N_VGND_c_425_n 0.00232396f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_215_297#_c_348_p N_VGND_c_425_n 0.00846569f $X=2.495 $Y=0.47 $X2=0
+ $Y2=0
cc_227 N_A_215_297#_c_261_n N_VGND_c_425_n 0.00232396f $X=2.98 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_A_215_297#_c_261_n N_VGND_c_426_n 3.34073e-19 $X=2.98 $Y=0.74 $X2=0
+ $Y2=0
cc_229 N_A_215_297#_c_266_n N_VGND_c_426_n 0.00524631f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_215_297#_c_340_p N_VGND_c_427_n 0.00625157f $X=1.65 $Y=0.47 $X2=0
+ $Y2=0
cc_231 N_A_215_297#_c_259_n N_VGND_c_427_n 0.00984491f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_215_297#_c_348_p N_VGND_c_427_n 0.00625722f $X=2.495 $Y=0.47 $X2=0
+ $Y2=0
cc_233 N_A_215_297#_c_261_n N_VGND_c_427_n 0.00637905f $X=2.98 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_215_297#_c_266_n N_VGND_c_427_n 0.00951738f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_357_n N_X_M1001_d 0.00399469f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_362_n X 0.0190559f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_357_n X 0.0105137f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_238 N_X_c_400_n N_VGND_c_426_n 0.00892672f $X=3.51 $Y=0.587 $X2=0 $Y2=0
cc_239 N_X_M1008_d N_VGND_c_427_n 0.00416042f $X=3.27 $Y=0.235 $X2=0 $Y2=0
cc_240 N_X_c_400_n N_VGND_c_427_n 0.00941771f $X=3.51 $Y=0.587 $X2=0 $Y2=0

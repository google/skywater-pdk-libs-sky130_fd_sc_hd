* File: sky130_fd_sc_hd__inv_4.spice.SKY130_FD_SC_HD__INV_4.pxi
* Created: Thu Aug 27 14:22:46 2020
* 
x_PM_SKY130_FD_SC_HD__INV_4%A N_A_c_39_n N_A_M1002_g N_A_M1000_g N_A_c_40_n
+ N_A_M1003_g N_A_M1001_g N_A_c_41_n N_A_M1004_g N_A_M1005_g N_A_c_42_n
+ N_A_M1006_g N_A_M1007_g A A A A N_A_c_44_n N_A_c_45_n
+ PM_SKY130_FD_SC_HD__INV_4%A
x_PM_SKY130_FD_SC_HD__INV_4%VPWR N_VPWR_M1000_s N_VPWR_M1001_s N_VPWR_M1007_s
+ N_VPWR_c_117_n N_VPWR_c_118_n N_VPWR_c_119_n N_VPWR_c_120_n N_VPWR_c_121_n
+ VPWR N_VPWR_c_122_n N_VPWR_c_123_n N_VPWR_c_124_n N_VPWR_c_116_n
+ PM_SKY130_FD_SC_HD__INV_4%VPWR
x_PM_SKY130_FD_SC_HD__INV_4%Y N_Y_M1002_s N_Y_M1004_s N_Y_M1000_d N_Y_M1005_d
+ N_Y_c_156_n N_Y_c_159_n N_Y_c_163_n N_Y_c_151_n N_Y_c_152_n N_Y_c_174_n
+ N_Y_c_177_n Y Y Y N_Y_c_187_n PM_SKY130_FD_SC_HD__INV_4%Y
x_PM_SKY130_FD_SC_HD__INV_4%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_M1006_d
+ N_VGND_c_217_n N_VGND_c_218_n N_VGND_c_219_n N_VGND_c_220_n N_VGND_c_221_n
+ VGND N_VGND_c_222_n N_VGND_c_223_n N_VGND_c_224_n N_VGND_c_225_n
+ PM_SKY130_FD_SC_HD__INV_4%VGND
cc_1 VNB N_A_c_39_n 0.0218814f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_c_40_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_c_41_n 0.0157835f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.995
cc_4 VNB N_A_c_42_n 0.0191475f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=0.995
cc_5 VNB A 0.00932659f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.105
cc_6 VNB N_A_c_44_n 0.0338038f $X=-0.19 $Y=-0.24 $X2=0.445 $Y2=1.16
cc_7 VNB N_A_c_45_n 0.0604092f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_8 VNB N_VPWR_c_116_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.16
cc_9 VNB N_Y_c_151_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_152_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=0.995
cc_11 VNB Y 0.0330601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_217_n 0.0114137f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_13 VNB N_VGND_c_218_n 0.0170366f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.985
cc_14 VNB N_VGND_c_219_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=0.56
cc_15 VNB N_VGND_c_220_n 0.0115482f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.325
cc_16 VNB N_VGND_c_221_n 0.0166667f $X=-0.19 $Y=-0.24 $X2=1.36 $Y2=1.985
cc_17 VNB N_VGND_c_222_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=0.56
cc_18 VNB N_VGND_c_223_n 0.0166866f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_19 VNB N_VGND_c_224_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_20 VNB N_VGND_c_225_n 0.144872f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_21 VPB N_A_M1000_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_22 VPB N_A_M1001_g 0.0185065f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.985
cc_23 VPB N_A_M1005_g 0.0184996f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.985
cc_24 VPB N_A_M1007_g 0.0218766f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.985
cc_25 VPB A 7.73822e-19 $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.105
cc_26 VPB N_A_c_44_n 0.0114928f $X=-0.19 $Y=1.305 $X2=0.445 $Y2=1.16
cc_27 VPB N_A_c_45_n 0.0100156f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_28 VPB N_VPWR_c_117_n 0.0114158f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.56
cc_29 VPB N_VPWR_c_118_n 0.0427864f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.985
cc_30 VPB N_VPWR_c_119_n 0.00358901f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.325
cc_31 VPB N_VPWR_c_120_n 0.0121106f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.985
cc_32 VPB N_VPWR_c_121_n 0.00438892f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=0.995
cc_33 VPB N_VPWR_c_122_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.985
cc_34 VPB N_VPWR_c_123_n 0.017949f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_35 VPB N_VPWR_c_124_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_36 VPB N_VPWR_c_116_n 0.0480032f $X=-0.19 $Y=1.305 $X2=1.36 $Y2=1.16
cc_37 VPB Y 0.00964194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB Y 0.0100741f $X=-0.19 $Y=1.305 $X2=0.445 $Y2=1.16
cc_39 N_A_M1000_g N_VPWR_c_118_n 0.00322031f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_40 A N_VPWR_c_118_n 0.0211311f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_41 N_A_c_44_n N_VPWR_c_118_n 0.00610847f $X=0.445 $Y=1.16 $X2=0 $Y2=0
cc_42 N_A_M1001_g N_VPWR_c_119_n 0.00146448f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_43 N_A_M1005_g N_VPWR_c_119_n 0.00146448f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_44 N_A_M1007_g N_VPWR_c_121_n 0.0031902f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_VPWR_c_122_n 0.00541359f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_VPWR_c_122_n 0.00541359f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_VPWR_c_123_n 0.00541359f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_48 N_A_M1007_g N_VPWR_c_123_n 0.00541359f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_VPWR_c_116_n 0.0105004f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_M1001_g N_VPWR_c_116_n 0.00950154f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_51 N_A_M1005_g N_VPWR_c_116_n 0.00950154f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A_M1007_g N_VPWR_c_116_n 0.0105004f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_53 N_A_c_39_n N_Y_c_156_n 0.0125306f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_c_40_n N_Y_c_156_n 0.0076511f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_55 N_A_c_41_n N_Y_c_156_n 5.48633e-19 $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A_M1000_g N_Y_c_159_n 0.00229676f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_Y_c_159_n 8.84614e-19 $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_58 A N_Y_c_159_n 0.0213676f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_c_45_n N_Y_c_159_n 0.00209661f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_Y_c_163_n 0.00902485f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_Y_c_163_n 0.00973632f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_Y_c_163_n 6.21474e-19 $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_c_40_n N_Y_c_151_n 0.00870364f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_c_41_n N_Y_c_151_n 0.00870364f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_65 A N_Y_c_151_n 0.0608989f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A_c_45_n N_Y_c_151_n 0.00222133f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_c_39_n N_Y_c_152_n 0.0110654f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A_c_40_n N_Y_c_152_n 0.00301106f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_69 A N_Y_c_152_n 0.0269421f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_45_n N_Y_c_152_n 0.00230339f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_40_n N_Y_c_174_n 5.49422e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_c_41_n N_Y_c_174_n 0.00777159f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_42_n N_Y_c_174_n 0.0125136f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A_M1001_g N_Y_c_177_n 5.61575e-19 $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1005_g N_Y_c_177_n 0.00950901f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1007_g N_Y_c_177_n 0.0249522f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_77 N_A_c_41_n Y 0.00314333f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_c_42_n Y 0.037092f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_79 A Y 0.0204697f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_c_45_n Y 0.00222133f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1005_g Y 0.00128027f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_M1007_g Y 0.0155463f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_c_45_n Y 0.00202298f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_M1001_g N_Y_c_187_n 0.0107189f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_Y_c_187_n 0.0107189f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_86 A N_Y_c_187_n 0.0516972f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_c_45_n N_Y_c_187_n 0.00201785f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_c_39_n N_VGND_c_218_n 0.00322031f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_89 A N_VGND_c_218_n 0.00872088f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_44_n N_VGND_c_218_n 0.00522062f $X=0.445 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_c_40_n N_VGND_c_219_n 0.00146448f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_c_41_n N_VGND_c_219_n 0.00146448f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_42_n N_VGND_c_221_n 0.00321269f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_c_39_n N_VGND_c_222_n 0.00541359f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_c_40_n N_VGND_c_222_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_c_41_n N_VGND_c_223_n 0.0042235f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_42_n N_VGND_c_223_n 0.0042235f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_c_39_n N_VGND_c_225_n 0.0105004f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_40_n N_VGND_c_225_n 0.0057163f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_c_41_n N_VGND_c_225_n 0.00573094f $X=1.36 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_42_n N_VGND_c_225_n 0.0067298f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_102 N_VPWR_c_116_n N_Y_M1000_d 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_103 N_VPWR_c_116_n N_Y_M1005_d 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_104 N_VPWR_c_122_n N_Y_c_163_n 0.0189039f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_105 N_VPWR_c_116_n N_Y_c_163_n 0.0122217f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_106 N_VPWR_c_123_n N_Y_c_177_n 0.0189039f $X=1.905 $Y=2.72 $X2=0 $Y2=0
cc_107 N_VPWR_c_116_n N_Y_c_177_n 0.0122217f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_108 N_VPWR_M1007_s Y 6.41575e-19 $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_109 N_VPWR_M1007_s Y 0.00505197f $X=1.855 $Y=1.485 $X2=0 $Y2=0
cc_110 N_VPWR_c_121_n Y 0.0074969f $X=1.99 $Y=2.34 $X2=0 $Y2=0
cc_111 N_VPWR_M1001_s N_Y_c_187_n 0.00311483f $X=1.015 $Y=1.485 $X2=0 $Y2=0
cc_112 N_VPWR_c_119_n N_Y_c_187_n 0.0126919f $X=1.15 $Y=2 $X2=0 $Y2=0
cc_113 N_Y_c_151_n N_VGND_M1003_d 0.001659f $X=1.405 $Y=0.815 $X2=0 $Y2=0
cc_114 Y N_VGND_M1006_d 0.00283816f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_115 N_Y_c_151_n N_VGND_c_219_n 0.0116647f $X=1.405 $Y=0.815 $X2=0 $Y2=0
cc_116 Y N_VGND_c_220_n 2.30187e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_117 Y N_VGND_c_221_n 0.0186601f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_118 N_Y_c_156_n N_VGND_c_222_n 0.0188551f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_119 N_Y_c_151_n N_VGND_c_222_n 0.00198695f $X=1.405 $Y=0.815 $X2=0 $Y2=0
cc_120 N_Y_c_151_n N_VGND_c_223_n 0.00400646f $X=1.405 $Y=0.815 $X2=0 $Y2=0
cc_121 N_Y_c_174_n N_VGND_c_223_n 0.0185141f $X=1.57 $Y=0.42 $X2=0 $Y2=0
cc_122 N_Y_M1002_s N_VGND_c_225_n 0.00215201f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_123 N_Y_M1004_s N_VGND_c_225_n 0.00215201f $X=1.435 $Y=0.235 $X2=0 $Y2=0
cc_124 N_Y_c_156_n N_VGND_c_225_n 0.0122069f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_125 N_Y_c_151_n N_VGND_c_225_n 0.0122828f $X=1.405 $Y=0.815 $X2=0 $Y2=0
cc_126 N_Y_c_174_n N_VGND_c_225_n 0.0121046f $X=1.57 $Y=0.42 $X2=0 $Y2=0
cc_127 Y N_VGND_c_225_n 0.00139502f $X=1.985 $Y=0.765 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__o311a_2.spice.pex
* Created: Thu Aug 27 14:39:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O311A_2%A_91_21# 1 2 3 10 12 15 17 19 22 26 27 29 30
+ 32 33 34 36 38 39 40 42 43 45 50
c110 26 0 1.7983e-19 $X=1.16 $Y=1.16
r111 56 58 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.53 $Y=1.16
+ $X2=0.95 $Y2=1.16
r112 50 52 15.3743 $w=5.83e-07 $l=4.25e-07 $layer=LI1_cond $X=3.762 $Y=0.4
+ $X2=3.762 $Y2=0.825
r113 43 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.91 $Y=1.58
+ $X2=3.555 $Y2=1.58
r114 43 45 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=3.91 $Y=1.665
+ $X2=3.91 $Y2=1.815
r115 42 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=1.495
+ $X2=3.555 $Y2=1.58
r116 42 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.555 $Y=1.495
+ $X2=3.555 $Y2=0.825
r117 39 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=1.58
+ $X2=3.555 $Y2=1.58
r118 39 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.47 $Y=1.58
+ $X2=3.175 $Y2=1.58
r119 36 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=2.295
+ $X2=3.01 $Y2=2.38
r120 36 38 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.01 $Y=2.295
+ $X2=3.01 $Y2=1.68
r121 35 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.01 $Y=1.665
+ $X2=3.175 $Y2=1.58
r122 35 38 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.01 $Y=1.665
+ $X2=3.01 $Y2=1.68
r123 33 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=2.38
+ $X2=3.01 $Y2=2.38
r124 33 34 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.845 $Y=2.38
+ $X2=1.81 $Y2=2.38
r125 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.725 $Y=2.295
+ $X2=1.81 $Y2=2.38
r126 31 32 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.725 $Y=1.665
+ $X2=1.725 $Y2=2.295
r127 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.64 $Y=1.58
+ $X2=1.725 $Y2=1.665
r128 29 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.64 $Y=1.58
+ $X2=1.245 $Y2=1.58
r129 27 58 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=0.95 $Y2=1.16
r130 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.16 $X2=1.16 $Y2=1.16
r131 24 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.16 $Y=1.495
+ $X2=1.245 $Y2=1.58
r132 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.16 $Y=1.495
+ $X2=1.16 $Y2=1.16
r133 20 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.325
+ $X2=0.95 $Y2=1.16
r134 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.95 $Y=1.325
+ $X2=0.95 $Y2=1.985
r135 17 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=1.16
r136 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=0.56
r137 13 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.16
r138 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.53 $Y=1.325
+ $X2=0.53 $Y2=1.985
r139 10 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=0.995
+ $X2=0.53 $Y2=1.16
r140 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.53 $Y=0.995
+ $X2=0.53 $Y2=0.56
r141 3 45 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=1.485 $X2=3.88 $Y2=1.815
r142 2 48 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.485 $X2=3.01 $Y2=2.36
r143 2 38 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.485 $X2=3.01 $Y2=1.68
r144 1 50 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.745
+ $Y=0.235 $X2=3.88 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%A1 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.16
+ $X2=1.665 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.16
+ $X2=1.665 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.16 $X2=1.665 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.725 $Y=1.985
+ $X2=1.725 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.725 $Y=0.56
+ $X2=1.725 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%A2 3 6 8 9 10 15 16 17
c36 16 0 5.25348e-20 $X=2.165 $Y=1.16
r37 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=1.16
+ $X2=2.165 $Y2=1.325
r38 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=1.16
+ $X2=2.165 $Y2=0.995
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.16 $X2=2.165 $Y2=1.16
r40 9 10 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.115 $Y=1.53
+ $X2=2.115 $Y2=1.87
r41 9 29 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.115 $Y=1.53
+ $X2=2.115 $Y2=1.325
r42 8 29 5.12956 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.085 $Y=1.19
+ $X2=2.085 $Y2=1.325
r43 8 16 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.085 $Y=1.19 $X2=2.085
+ $Y2=1.16
r44 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.225 $Y=1.985
+ $X2=2.225 $Y2=1.325
r45 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.225 $Y=0.56
+ $X2=2.225 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%A3 3 6 8 9 10 15 16 17
r35 15 18 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=1.325
r36 15 17 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=0.995
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.16 $X2=2.645 $Y2=1.16
r38 9 10 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.557 $Y=1.53
+ $X2=2.557 $Y2=1.87
r39 9 29 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=2.557 $Y=1.53
+ $X2=2.557 $Y2=1.325
r40 8 29 5.81314 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.585 $Y=1.19
+ $X2=2.585 $Y2=1.325
r41 8 16 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.585 $Y=1.19 $X2=2.585
+ $Y2=1.16
r42 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.795 $Y=1.985
+ $X2=2.795 $Y2=1.325
r43 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.795 $Y=0.56
+ $X2=2.795 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%B1 3 7 8 11 12 13
r35 11 14 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.232 $Y=1.16
+ $X2=3.232 $Y2=1.325
r36 11 13 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.232 $Y=1.16
+ $X2=3.232 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.215
+ $Y=1.16 $X2=3.215 $Y2=1.16
r38 8 12 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.985 $Y=1.16
+ $X2=3.215 $Y2=1.16
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.56 $X2=3.31
+ $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.22 $Y=1.985
+ $X2=3.22 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%C1 1 3 6 8 13
r26 10 13 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.67 $Y=1.16
+ $X2=3.895 $Y2=1.16
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=1.16 $X2=3.895 $Y2=1.16
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.325
+ $X2=3.67 $Y2=1.16
r29 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.325 $X2=3.67
+ $Y2=1.985
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.995
+ $X2=3.67 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.67 $Y=0.995 $X2=3.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%VPWR 1 2 3 10 12 16 20 24 26 28 38 39 45 48
c58 2 0 1.27295e-19 $X=1.025 $Y=1.485
r59 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 39 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 36 48 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.477 $Y2=2.72
r64 36 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 32 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r68 32 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r69 31 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 29 45 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.272 $Y2=2.72
r72 29 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.61 $Y2=2.72
r73 28 48 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.36 $Y=2.72
+ $X2=3.477 $Y2=2.72
r74 28 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.36 $Y=2.72 $X2=2.99
+ $Y2=2.72
r75 26 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 26 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 22 48 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.477 $Y=2.635
+ $X2=3.477 $Y2=2.72
r78 22 24 31.1405 $w=2.33e-07 $l=6.35e-07 $layer=LI1_cond $X=3.477 $Y=2.635
+ $X2=3.477 $Y2=2
r79 18 45 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.272 $Y=2.635
+ $X2=1.272 $Y2=2.72
r80 18 20 17.9431 $w=3.93e-07 $l=6.15e-07 $layer=LI1_cond $X=1.272 $Y=2.635
+ $X2=1.272 $Y2=2.02
r81 17 42 4.4818 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=2.72 $X2=0.19
+ $Y2=2.72
r82 16 45 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=1.272 $Y2=2.72
r83 16 17 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=0.38 $Y2=2.72
r84 12 15 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.232 $Y=1.66
+ $X2=0.232 $Y2=2.34
r85 10 42 2.99573 $w=2.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.232 $Y=2.635
+ $X2=0.19 $Y2=2.72
r86 10 15 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.232 $Y=2.635
+ $X2=0.232 $Y2=2.34
r87 3 24 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=3.295
+ $Y=1.485 $X2=3.445 $Y2=2
r88 2 20 300 $w=1.7e-07 $l=6.56258e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=1.485 $X2=1.295 $Y2=2.02
r89 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r90 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%X 1 2 7 8 9 10 11 12 13 21
r22 13 42 4.22021 $w=3.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.727 $Y=2.21
+ $X2=0.727 $Y2=2.34
r23 12 13 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.727 $Y=1.87
+ $X2=0.727 $Y2=2.21
r24 12 36 6.81727 $w=3.53e-07 $l=2.1e-07 $layer=LI1_cond $X=0.727 $Y=1.87
+ $X2=0.727 $Y2=1.66
r25 11 36 4.22021 $w=3.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.727 $Y=1.53
+ $X2=0.727 $Y2=1.66
r26 11 32 6.97958 $w=3.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.727 $Y=1.53
+ $X2=0.727 $Y2=1.315
r27 10 21 2.04183 $w=2.6e-07 $l=1.91413e-07 $layer=LI1_cond $X=0.727 $Y=1.155
+ $X2=0.55 $Y2=1.185
r28 10 25 4.39111 $w=3.15e-07 $l=1.78885e-07 $layer=LI1_cond $X=0.727 $Y=1.155
+ $X2=0.687 $Y2=0.995
r29 10 32 4.39111 $w=3.15e-07 $l=1.6e-07 $layer=LI1_cond $X=0.727 $Y=1.155
+ $X2=0.727 $Y2=1.315
r30 9 25 6.07652 $w=2.73e-07 $l=1.45e-07 $layer=LI1_cond $X=0.687 $Y=0.85
+ $X2=0.687 $Y2=0.995
r31 8 9 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=0.687 $Y=0.51
+ $X2=0.687 $Y2=0.85
r32 7 21 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.235 $Y=1.185
+ $X2=0.55 $Y2=1.185
r33 2 42 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.74 $Y2=2.34
r34 2 36 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.74 $Y2=1.66
r35 1 8 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.235 $X2=0.74 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r56 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r57 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r59 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r60 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r61 36 39 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r62 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 34 49 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.487
+ $Y2=0
r64 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.99
+ $Y2=0
r65 33 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r66 33 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r67 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r68 30 46 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.33
+ $Y2=0
r69 30 32 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=2.07
+ $Y2=0
r70 29 49 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=2.487
+ $Y2=0
r71 29 32 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=2.07
+ $Y2=0
r72 28 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r73 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r74 25 43 4.4818 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r75 25 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.69
+ $Y2=0
r76 24 46 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.33
+ $Y2=0
r77 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.69
+ $Y2=0
r78 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r79 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r80 18 49 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0
r81 18 20 8.45125 $w=3.73e-07 $l=2.75e-07 $layer=LI1_cond $X=2.487 $Y=0.085
+ $X2=2.487 $Y2=0.36
r82 14 46 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=0.085
+ $X2=1.33 $Y2=0
r83 14 16 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.33 $Y=0.085
+ $X2=1.33 $Y2=0.36
r84 10 43 2.99573 $w=2.95e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.232 $Y=0.085
+ $X2=0.19 $Y2=0
r85 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.232 $Y=0.085
+ $X2=0.232 $Y2=0.38
r86 3 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.235 $X2=2.51 $Y2=0.36
r87 2 16 45.5 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_NDIFF $count=4 $X=1.025
+ $Y=0.235 $X2=1.5 $Y2=0.36
r88 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O311A_2%A_360_47# 1 2 9 11 12 13 15
r21 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.655
+ $X2=3.055 $Y2=0.74
r22 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.055 $Y=0.655
+ $X2=3.055 $Y2=0.4
r23 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0.74
+ $X2=3.055 $Y2=0.74
r24 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.89 $Y=0.74
+ $X2=2.12 $Y2=0.74
r25 7 12 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=1.977 $Y=0.655
+ $X2=2.12 $Y2=0.74
r26 7 9 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=1.977 $Y=0.655
+ $X2=1.977 $Y2=0.56
r27 2 18 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.055 $Y2=0.74
r28 2 15 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.055 $Y2=0.4
r29 1 9 182 $w=1.7e-07 $l=4.01092e-07 $layer=licon1_NDIFF $count=1 $X=1.8
+ $Y=0.235 $X2=1.97 $Y2=0.56
.ends


* File: sky130_fd_sc_hd__a21bo_4.spice.SKY130_FD_SC_HD__A21BO_4.pxi
* Created: Thu Aug 27 14:00:16 2020
* 
x_PM_SKY130_FD_SC_HD__A21BO_4%B1_N N_B1_N_M1021_g N_B1_N_M1017_g B1_N
+ N_B1_N_c_98_n N_B1_N_c_99_n PM_SKY130_FD_SC_HD__A21BO_4%B1_N
x_PM_SKY130_FD_SC_HD__A21BO_4%A_205_21# N_A_205_21#_M1014_d N_A_205_21#_M1002_s
+ N_A_205_21#_M1000_s N_A_205_21#_c_129_n N_A_205_21#_M1005_g
+ N_A_205_21#_M1006_g N_A_205_21#_c_130_n N_A_205_21#_M1007_g
+ N_A_205_21#_M1009_g N_A_205_21#_c_131_n N_A_205_21#_M1008_g
+ N_A_205_21#_M1010_g N_A_205_21#_c_132_n N_A_205_21#_M1019_g
+ N_A_205_21#_M1018_g N_A_205_21#_c_210_p N_A_205_21#_c_133_n
+ N_A_205_21#_c_149_p N_A_205_21#_c_244_p N_A_205_21#_c_134_n
+ N_A_205_21#_c_154_p N_A_205_21#_c_135_n N_A_205_21#_c_136_n
+ N_A_205_21#_c_151_p N_A_205_21#_c_183_p PM_SKY130_FD_SC_HD__A21BO_4%A_205_21#
x_PM_SKY130_FD_SC_HD__A21BO_4%A_42_47# N_A_42_47#_M1021_s N_A_42_47#_M1017_s
+ N_A_42_47#_c_268_n N_A_42_47#_M1014_g N_A_42_47#_M1000_g N_A_42_47#_c_269_n
+ N_A_42_47#_M1020_g N_A_42_47#_M1003_g N_A_42_47#_c_270_n N_A_42_47#_c_277_n
+ N_A_42_47#_c_278_n N_A_42_47#_c_279_n N_A_42_47#_c_271_n N_A_42_47#_c_272_n
+ N_A_42_47#_c_281_n N_A_42_47#_c_273_n PM_SKY130_FD_SC_HD__A21BO_4%A_42_47#
x_PM_SKY130_FD_SC_HD__A21BO_4%A2 N_A2_M1015_g N_A2_M1004_g N_A2_M1013_g
+ N_A2_M1016_g N_A2_c_372_n N_A2_c_373_n N_A2_c_374_n N_A2_c_375_n N_A2_c_376_n
+ N_A2_c_377_n N_A2_c_417_p A2 N_A2_c_378_n N_A2_c_379_n N_A2_c_420_p A2
+ PM_SKY130_FD_SC_HD__A21BO_4%A2
x_PM_SKY130_FD_SC_HD__A21BO_4%A1 N_A1_c_451_n N_A1_M1002_g N_A1_M1001_g
+ N_A1_c_452_n N_A1_M1012_g N_A1_M1011_g A1 N_A1_c_453_n
+ PM_SKY130_FD_SC_HD__A21BO_4%A1
x_PM_SKY130_FD_SC_HD__A21BO_4%VPWR N_VPWR_M1017_d N_VPWR_M1009_s N_VPWR_M1018_s
+ N_VPWR_M1015_s N_VPWR_M1011_d N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n
+ VPWR N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_496_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n
+ PM_SKY130_FD_SC_HD__A21BO_4%VPWR
x_PM_SKY130_FD_SC_HD__A21BO_4%X N_X_M1005_s N_X_M1008_s N_X_M1006_d N_X_M1010_d
+ N_X_c_604_n N_X_c_605_n X N_X_c_617_n X N_X_c_618_n
+ PM_SKY130_FD_SC_HD__A21BO_4%X
x_PM_SKY130_FD_SC_HD__A21BO_4%A_603_297# N_A_603_297#_M1000_d
+ N_A_603_297#_M1003_d N_A_603_297#_M1001_s N_A_603_297#_M1016_d
+ N_A_603_297#_c_646_n N_A_603_297#_c_647_n N_A_603_297#_c_682_n
+ N_A_603_297#_c_643_n N_A_603_297#_c_644_n N_A_603_297#_c_645_n
+ N_A_603_297#_c_693_n PM_SKY130_FD_SC_HD__A21BO_4%A_603_297#
x_PM_SKY130_FD_SC_HD__A21BO_4%VGND N_VGND_M1021_d N_VGND_M1007_d N_VGND_M1019_d
+ N_VGND_M1020_s N_VGND_M1013_d N_VGND_c_696_n N_VGND_c_697_n N_VGND_c_698_n
+ N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n
+ N_VGND_c_704_n VGND N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n
+ N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n PM_SKY130_FD_SC_HD__A21BO_4%VGND
cc_1 VNB B1_N 0.00528546f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_2 VNB N_B1_N_c_98_n 0.0259538f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.16
cc_3 VNB N_B1_N_c_99_n 0.0195714f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=0.995
cc_4 VNB N_A_205_21#_c_129_n 0.0150161f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.16
cc_5 VNB N_A_205_21#_c_130_n 0.0159846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_205_21#_c_131_n 0.016003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_205_21#_c_132_n 0.0193863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_205_21#_c_133_n 0.00241062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_205_21#_c_134_n 0.00192199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_205_21#_c_135_n 0.0107246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_205_21#_c_136_n 0.0724083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_42_47#_c_268_n 0.0190644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_42_47#_c_269_n 0.0165854f $X=-0.19 $Y=-0.24 $X2=0.665 $Y2=1.325
cc_14 VNB N_A_42_47#_c_270_n 0.0234483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_42_47#_c_271_n 0.0053415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_42_47#_c_272_n 0.0255593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_42_47#_c_273_n 0.0445355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_372_n 4.44522e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_373_n 0.00795453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_374_n 0.0101098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_375_n 0.0271516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_c_376_n 0.0185455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A2_c_377_n 0.00539737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A2_c_378_n 0.0161936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A2_c_379_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A1_c_451_n 0.0158558f $X=-0.19 $Y=-0.24 $X2=0.67 $Y2=0.995
cc_27 VNB N_A1_c_452_n 0.0162494f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_28 VNB N_A1_c_453_n 0.0320785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_496_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.00419828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_696_n 3.99187e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_697_n 0.0122657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_698_n 3.21528e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_699_n 0.0136763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_700_n 0.00215534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_701_n 0.012531f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_702_n 0.0327763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_703_n 0.0196166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_704_n 0.0044932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_705_n 0.0381373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_706_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_707_n 0.0161586f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_708_n 0.0183347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_709_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_710_n 0.298366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_B1_N_M1017_g 0.0222711f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_47 VPB B1_N 0.00277322f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_48 VPB N_B1_N_c_98_n 0.00478302f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=1.16
cc_49 VPB N_A_205_21#_M1006_g 0.0171979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_205_21#_M1009_g 0.0185175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_205_21#_M1010_g 0.0185456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_205_21#_M1018_g 0.021555f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_205_21#_c_134_n 0.00225717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_205_21#_c_135_n 0.00105623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_205_21#_c_136_n 0.0153173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_42_47#_M1000_g 0.0229436f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=1.16
cc_57 VPB N_A_42_47#_M1003_g 0.0187512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_42_47#_c_270_n 0.0249593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_42_47#_c_277_n 0.00347844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_42_47#_c_278_n 0.00576583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_42_47#_c_279_n 0.0125667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_42_47#_c_271_n 0.00142271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_42_47#_c_281_n 0.0334843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_42_47#_c_273_n 0.0103646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_M1015_g 0.0179332f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=0.56
cc_66 VPB N_A2_M1016_g 0.0244532f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=0.995
cc_67 VPB N_A2_c_372_n 0.00149191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A2_c_375_n 0.00506794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A2_c_376_n 0.00468017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB A2 0.00153697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A1_M1001_g 0.0183773f $X=-0.19 $Y=1.305 $X2=0.67 $Y2=1.985
cc_72 VPB N_A1_M1011_g 0.0183773f $X=-0.19 $Y=1.305 $X2=0.665 $Y2=0.995
cc_73 VPB A1 0.00282525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A1_c_453_n 0.00450322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_497_n 3.99129e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_498_n 0.0122674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_499_n 3.08203e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_500_n 0.00553251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_501_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_502_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_503_n 0.0190371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_504_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_505_n 0.0121314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_506_n 0.0362233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_507_n 0.0117235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_508_n 0.0174547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_496_n 0.056194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_510_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_511_n 0.00516648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_512_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_513_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB X 0.00278331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_603_297#_c_643_n 0.00330706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_603_297#_c_644_n 0.00767904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_603_297#_c_645_n 0.021001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 N_B1_N_c_99_n N_A_205_21#_c_129_n 0.0242787f $X=0.665 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_N_M1017_g N_A_205_21#_M1006_g 0.0435088f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_98 B1_N N_A_205_21#_c_136_n 0.00198219f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B1_N_c_98_n N_A_205_21#_c_136_n 0.0196742f $X=0.665 $Y=1.16 $X2=0 $Y2=0
cc_100 B1_N N_A_42_47#_M1017_s 0.00193083f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B1_N_M1017_g N_A_42_47#_c_270_n 0.00430887f $X=0.67 $Y=1.985 $X2=0
+ $Y2=0
cc_102 B1_N N_A_42_47#_c_270_n 0.0495468f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B1_N_c_98_n N_A_42_47#_c_270_n 0.00248191f $X=0.665 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_N_c_99_n N_A_42_47#_c_270_n 0.00225981f $X=0.665 $Y=0.995 $X2=0
+ $Y2=0
cc_105 N_B1_N_M1017_g N_A_42_47#_c_277_n 0.0102245f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_106 B1_N N_A_42_47#_c_277_n 0.00836872f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_107 B1_N N_A_42_47#_c_272_n 0.00334456f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B1_N_c_98_n N_A_42_47#_c_272_n 2.09046e-19 $X=0.665 $Y=1.16 $X2=0 $Y2=0
cc_109 B1_N N_A_42_47#_c_281_n 0.00330765f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_110 B1_N N_VPWR_M1017_d 0.0015924f $X=0.605 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 N_B1_N_M1017_g N_VPWR_c_497_n 0.0078488f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B1_N_M1017_g N_VPWR_c_503_n 0.00351072f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_113 N_B1_N_M1017_g N_VPWR_c_496_n 0.00514525f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B1_N_M1017_g X 5.09615e-19 $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_115 B1_N X 0.0429209f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B1_N_c_98_n X 0.00107591f $X=0.665 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_N_c_99_n X 0.00135281f $X=0.665 $Y=0.995 $X2=0 $Y2=0
cc_118 B1_N N_VGND_c_696_n 0.00292457f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B1_N_c_99_n N_VGND_c_696_n 0.00887116f $X=0.665 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B1_N_c_99_n N_VGND_c_703_n 0.00447018f $X=0.665 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_N_c_99_n N_VGND_c_710_n 0.0088013f $X=0.665 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_205_21#_c_133_n N_A_42_47#_c_268_n 0.00322808f $X=2.725 $Y=0.995
+ $X2=0 $Y2=0
cc_123 N_A_205_21#_c_149_p N_A_42_47#_c_268_n 0.0152399f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_124 N_A_205_21#_c_134_n N_A_42_47#_c_268_n 0.00141413f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_125 N_A_205_21#_c_151_p N_A_42_47#_c_268_n 2.88686e-19 $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_126 N_A_205_21#_c_134_n N_A_42_47#_M1000_g 0.00111632f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_127 N_A_205_21#_c_134_n N_A_42_47#_c_269_n 0.00260329f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_128 N_A_205_21#_c_154_p N_A_42_47#_c_269_n 0.0146368f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_129 N_A_205_21#_c_134_n N_A_42_47#_M1003_g 0.0017889f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_130 N_A_205_21#_M1006_g N_A_42_47#_c_277_n 0.0114959f $X=1.1 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_205_21#_M1009_g N_A_42_47#_c_277_n 0.0115486f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_205_21#_M1010_g N_A_42_47#_c_277_n 0.0115486f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_205_21#_M1018_g N_A_42_47#_c_277_n 0.0138783f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_205_21#_c_135_n N_A_42_47#_c_277_n 0.00232617f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_205_21#_c_136_n N_A_42_47#_c_277_n 0.0013386f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_205_21#_M1018_g N_A_42_47#_c_278_n 0.0108833f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_205_21#_M1018_g N_A_42_47#_c_279_n 0.00629266f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_205_21#_c_134_n N_A_42_47#_c_279_n 0.0117881f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_139 N_A_205_21#_c_135_n N_A_42_47#_c_279_n 0.0088738f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_205_21#_c_151_p N_A_42_47#_c_279_n 0.00593425f $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_141 N_A_205_21#_M1018_g N_A_42_47#_c_271_n 7.46305e-19 $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_205_21#_c_149_p N_A_42_47#_c_271_n 0.01709f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_143 N_A_205_21#_c_134_n N_A_42_47#_c_271_n 0.0256547f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_144 N_A_205_21#_c_135_n N_A_42_47#_c_271_n 0.0212365f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_205_21#_c_136_n N_A_42_47#_c_271_n 0.00172781f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_205_21#_c_151_p N_A_42_47#_c_271_n 0.0010056f $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_147 N_A_205_21#_c_149_p N_A_42_47#_c_273_n 0.00114071f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_148 N_A_205_21#_c_134_n N_A_42_47#_c_273_n 0.0188095f $X=3.56 $Y=1.62 $X2=0
+ $Y2=0
cc_149 N_A_205_21#_c_135_n N_A_42_47#_c_273_n 8.52775e-19 $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_205_21#_c_136_n N_A_42_47#_c_273_n 0.00654167f $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_205_21#_c_134_n N_A2_c_372_n 0.00447131f $X=3.56 $Y=1.62 $X2=0 $Y2=0
cc_152 N_A_205_21#_c_134_n N_A2_c_376_n 4.5982e-19 $X=3.56 $Y=1.62 $X2=0 $Y2=0
cc_153 N_A_205_21#_c_154_p N_A2_c_376_n 0.00231315f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_154 N_A_205_21#_c_134_n N_A2_c_377_n 0.0111268f $X=3.56 $Y=1.62 $X2=0 $Y2=0
cc_155 N_A_205_21#_c_154_p N_A2_c_377_n 0.0246715f $X=4.685 $Y=0.755 $X2=0 $Y2=0
cc_156 N_A_205_21#_c_154_p N_A2_c_378_n 0.0115203f $X=4.685 $Y=0.755 $X2=0 $Y2=0
cc_157 N_A_205_21#_c_183_p N_A2_c_379_n 0.00126506f $X=4.82 $Y=0.57 $X2=0 $Y2=0
cc_158 N_A_205_21#_c_154_p N_A1_c_451_n 0.011299f $X=4.685 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_205_21#_c_183_p N_A1_c_452_n 0.00875304f $X=4.82 $Y=0.57 $X2=0 $Y2=0
cc_160 N_A_205_21#_c_154_p A1 0.00681644f $X=4.685 $Y=0.755 $X2=0 $Y2=0
cc_161 N_A_205_21#_c_183_p A1 0.0167857f $X=4.82 $Y=0.57 $X2=0 $Y2=0
cc_162 N_A_205_21#_c_183_p N_A1_c_453_n 0.0021041f $X=4.82 $Y=0.57 $X2=0 $Y2=0
cc_163 N_A_205_21#_M1006_g N_VPWR_c_497_n 0.0076143f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_205_21#_M1009_g N_VPWR_c_497_n 0.00104385f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_205_21#_M1006_g N_VPWR_c_498_n 0.00351072f $X=1.1 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_205_21#_M1009_g N_VPWR_c_498_n 0.00351072f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_205_21#_M1006_g N_VPWR_c_499_n 0.00104385f $X=1.1 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_205_21#_M1009_g N_VPWR_c_499_n 0.00765006f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_205_21#_M1010_g N_VPWR_c_499_n 0.00762255f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_205_21#_M1018_g N_VPWR_c_499_n 0.00104065f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A_205_21#_M1010_g N_VPWR_c_500_n 0.00105243f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_205_21#_M1018_g N_VPWR_c_500_n 0.0089652f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A_205_21#_M1010_g N_VPWR_c_505_n 0.00351072f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_205_21#_M1018_g N_VPWR_c_505_n 0.00337001f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_175 N_A_205_21#_M1000_s N_VPWR_c_496_n 0.00224997f $X=3.425 $Y=1.485 $X2=0
+ $Y2=0
cc_176 N_A_205_21#_M1006_g N_VPWR_c_496_n 0.00411677f $X=1.1 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_205_21#_M1009_g N_VPWR_c_496_n 0.00411677f $X=1.53 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_205_21#_M1010_g N_VPWR_c_496_n 0.00411677f $X=1.96 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_205_21#_M1018_g N_VPWR_c_496_n 0.00397572f $X=2.39 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_205_21#_c_129_n N_X_c_604_n 0.00611988f $X=1.1 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_205_21#_c_130_n N_X_c_605_n 0.00972932f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_205_21#_c_131_n N_X_c_605_n 0.00972932f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_205_21#_c_132_n N_X_c_605_n 0.00326174f $X=2.39 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_205_21#_c_210_p N_X_c_605_n 0.0491543f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_205_21#_c_136_n N_X_c_605_n 0.00796547f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_205_21#_c_151_p N_X_c_605_n 0.00946301f $X=3.01 $Y=0.707 $X2=0 $Y2=0
cc_187 N_A_205_21#_c_129_n X 0.00420563f $X=1.1 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_205_21#_M1006_g X 0.0055312f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_205_21#_c_130_n X 0.00403073f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_205_21#_M1009_g X 0.0052446f $X=1.53 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_205_21#_c_210_p X 0.0255555f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_205_21#_c_136_n X 0.011804f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_205_21#_M1006_g N_X_c_617_n 0.0051775f $X=1.1 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_205_21#_M1009_g N_X_c_618_n 0.00901837f $X=1.53 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_205_21#_M1010_g N_X_c_618_n 0.00901837f $X=1.96 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_205_21#_M1018_g N_X_c_618_n 0.00603797f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_205_21#_c_210_p N_X_c_618_n 0.0415672f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_205_21#_c_135_n N_X_c_618_n 0.00222822f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_205_21#_c_136_n N_X_c_618_n 0.00756104f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_205_21#_M1018_g N_A_603_297#_c_646_n 0.00263244f $X=2.39 $Y=1.985
+ $X2=0 $Y2=0
cc_201 N_A_205_21#_M1000_s N_A_603_297#_c_647_n 0.00425956f $X=3.425 $Y=1.485
+ $X2=0 $Y2=0
cc_202 N_A_205_21#_c_134_n N_A_603_297#_c_647_n 0.00668159f $X=3.56 $Y=1.62
+ $X2=0 $Y2=0
cc_203 N_A_205_21#_c_134_n N_A_603_297#_c_643_n 0.00231527f $X=3.56 $Y=1.62
+ $X2=0 $Y2=0
cc_204 N_A_205_21#_c_154_p N_A_603_297#_c_643_n 0.00440519f $X=4.685 $Y=0.755
+ $X2=0 $Y2=0
cc_205 N_A_205_21#_c_133_n N_VGND_M1019_d 0.00318132f $X=2.725 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_205_21#_c_149_p N_VGND_M1019_d 0.00498018f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_207 N_A_205_21#_c_151_p N_VGND_M1019_d 0.0139699f $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_208 N_A_205_21#_c_154_p N_VGND_M1020_s 0.00540394f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_209 N_A_205_21#_c_129_n N_VGND_c_696_n 0.0076133f $X=1.1 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_205_21#_c_130_n N_VGND_c_696_n 0.00104439f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_205_21#_c_129_n N_VGND_c_697_n 0.00350947f $X=1.1 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_205_21#_c_130_n N_VGND_c_697_n 0.00351072f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_205_21#_c_129_n N_VGND_c_698_n 0.00104385f $X=1.1 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_205_21#_c_130_n N_VGND_c_698_n 0.00765006f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_205_21#_c_131_n N_VGND_c_698_n 0.00802115f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_205_21#_c_132_n N_VGND_c_698_n 0.00109177f $X=2.39 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_205_21#_c_149_p N_VGND_c_699_n 0.00289974f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_218 N_A_205_21#_c_244_p N_VGND_c_699_n 0.0113958f $X=3.56 $Y=0.42 $X2=0 $Y2=0
cc_219 N_A_205_21#_c_154_p N_VGND_c_699_n 0.00278663f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_220 N_A_205_21#_c_154_p N_VGND_c_700_n 0.0133243f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_221 N_A_205_21#_c_183_p N_VGND_c_700_n 0.00138436f $X=4.82 $Y=0.57 $X2=0
+ $Y2=0
cc_222 N_A_205_21#_c_154_p N_VGND_c_705_n 0.00696372f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_223 N_A_205_21#_c_183_p N_VGND_c_705_n 0.00778691f $X=4.82 $Y=0.57 $X2=0
+ $Y2=0
cc_224 N_A_205_21#_c_131_n N_VGND_c_707_n 0.00351072f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_205_21#_c_132_n N_VGND_c_707_n 0.00558173f $X=2.39 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_205_21#_c_132_n N_VGND_c_708_n 0.00729481f $X=2.39 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_205_21#_c_135_n N_VGND_c_708_n 0.004019f $X=2.445 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_205_21#_c_136_n N_VGND_c_708_n 3.74016e-19 $X=2.445 $Y=1.16 $X2=0
+ $Y2=0
cc_229 N_A_205_21#_c_151_p N_VGND_c_708_n 0.0443671f $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_230 N_A_205_21#_M1014_d N_VGND_c_710_n 0.00250439f $X=3.425 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_A_205_21#_M1002_s N_VGND_c_710_n 0.00237222f $X=4.685 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_205_21#_c_129_n N_VGND_c_710_n 0.00411477f $X=1.1 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_205_21#_c_130_n N_VGND_c_710_n 0.00411677f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_205_21#_c_131_n N_VGND_c_710_n 0.00411677f $X=1.96 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_205_21#_c_132_n N_VGND_c_710_n 0.0112602f $X=2.39 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_205_21#_c_149_p N_VGND_c_710_n 0.00470987f $X=3.475 $Y=0.7 $X2=0
+ $Y2=0
cc_237 N_A_205_21#_c_244_p N_VGND_c_710_n 0.00646998f $X=3.56 $Y=0.42 $X2=0
+ $Y2=0
cc_238 N_A_205_21#_c_154_p N_VGND_c_710_n 0.0189434f $X=4.685 $Y=0.755 $X2=0
+ $Y2=0
cc_239 N_A_205_21#_c_151_p N_VGND_c_710_n 0.0029858f $X=3.01 $Y=0.707 $X2=0
+ $Y2=0
cc_240 N_A_205_21#_c_183_p N_VGND_c_710_n 0.00961573f $X=4.82 $Y=0.57 $X2=0
+ $Y2=0
cc_241 N_A_205_21#_c_154_p A_861_47# 0.00492452f $X=4.685 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_242 N_A_42_47#_M1003_g N_A2_M1015_g 0.0258569f $X=3.77 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_42_47#_c_273_n N_A2_c_372_n 5.67187e-19 $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_42_47#_c_273_n N_A2_c_376_n 0.0221136f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_42_47#_c_273_n N_A2_c_377_n 0.00236109f $X=3.77 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_42_47#_c_269_n N_A2_c_378_n 0.0234488f $X=3.77 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_42_47#_c_277_n N_VPWR_M1017_d 0.00737383f $X=2.7 $Y=2.02 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_42_47#_c_277_n N_VPWR_M1009_s 0.00337117f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_249 N_A_42_47#_c_277_n N_VPWR_M1018_s 0.00871732f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_250 N_A_42_47#_c_278_n N_VPWR_M1018_s 0.00584651f $X=2.785 $Y=1.935 $X2=0
+ $Y2=0
cc_251 N_A_42_47#_c_279_n N_VPWR_M1018_s 7.69051e-19 $X=3.15 $Y=1.355 $X2=0
+ $Y2=0
cc_252 N_A_42_47#_c_277_n N_VPWR_c_497_n 0.0159085f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_253 N_A_42_47#_c_277_n N_VPWR_c_498_n 0.00846546f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_254 N_A_42_47#_c_277_n N_VPWR_c_499_n 0.0159085f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_255 N_A_42_47#_M1000_g N_VPWR_c_500_n 0.00443811f $X=3.35 $Y=1.985 $X2=0
+ $Y2=0
cc_256 N_A_42_47#_c_277_n N_VPWR_c_500_n 0.0212685f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_257 N_A_42_47#_M1003_g N_VPWR_c_501_n 0.00156191f $X=3.77 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_A_42_47#_c_277_n N_VPWR_c_503_n 0.00243617f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_259 N_A_42_47#_c_281_n N_VPWR_c_503_n 0.0310956f $X=0.335 $Y=2.02 $X2=0 $Y2=0
cc_260 N_A_42_47#_c_277_n N_VPWR_c_505_n 0.00839568f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_261 N_A_42_47#_M1000_g N_VPWR_c_506_n 0.00375019f $X=3.35 $Y=1.985 $X2=0
+ $Y2=0
cc_262 N_A_42_47#_M1003_g N_VPWR_c_506_n 0.00375019f $X=3.77 $Y=1.985 $X2=0
+ $Y2=0
cc_263 N_A_42_47#_c_277_n N_VPWR_c_506_n 0.00208183f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_264 N_A_42_47#_M1017_s N_VPWR_c_496_n 0.00228189f $X=0.33 $Y=1.485 $X2=0
+ $Y2=0
cc_265 N_A_42_47#_M1000_g N_VPWR_c_496_n 0.00669207f $X=3.35 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_A_42_47#_M1003_g N_VPWR_c_496_n 0.00534325f $X=3.77 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_A_42_47#_c_277_n N_VPWR_c_496_n 0.0394466f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_268 N_A_42_47#_c_281_n N_VPWR_c_496_n 0.0175664f $X=0.335 $Y=2.02 $X2=0 $Y2=0
cc_269 N_A_42_47#_c_277_n N_X_M1006_d 0.00444184f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_270 N_A_42_47#_c_277_n N_X_M1010_d 0.00450788f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_271 N_A_42_47#_c_270_n X 0.00358572f $X=0.217 $Y=1.795 $X2=0 $Y2=0
cc_272 N_A_42_47#_c_277_n N_X_c_617_n 0.0114206f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_273 N_A_42_47#_c_277_n N_X_c_618_n 0.0625887f $X=2.7 $Y=2.02 $X2=0 $Y2=0
cc_274 N_A_42_47#_c_278_n N_X_c_618_n 0.00873749f $X=2.785 $Y=1.935 $X2=0 $Y2=0
cc_275 N_A_42_47#_c_279_n N_A_603_297#_M1000_d 0.0033706f $X=3.15 $Y=1.355
+ $X2=-0.19 $Y2=-0.24
cc_276 N_A_42_47#_c_277_n N_A_603_297#_c_646_n 0.0132907f $X=2.7 $Y=2.02 $X2=0
+ $Y2=0
cc_277 N_A_42_47#_c_278_n N_A_603_297#_c_646_n 0.0166633f $X=2.785 $Y=1.935
+ $X2=0 $Y2=0
cc_278 N_A_42_47#_c_279_n N_A_603_297#_c_646_n 0.013188f $X=3.15 $Y=1.355 $X2=0
+ $Y2=0
cc_279 N_A_42_47#_M1000_g N_A_603_297#_c_647_n 0.0126862f $X=3.35 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_42_47#_M1003_g N_A_603_297#_c_647_n 0.0132272f $X=3.77 $Y=1.985 $X2=0
+ $Y2=0
cc_281 N_A_42_47#_M1003_g N_A_603_297#_c_643_n 5.54179e-19 $X=3.77 $Y=1.985
+ $X2=0 $Y2=0
cc_282 N_A_42_47#_c_268_n N_VGND_c_699_n 0.00393283f $X=3.35 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_42_47#_c_269_n N_VGND_c_699_n 0.00430182f $X=3.77 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_42_47#_c_269_n N_VGND_c_700_n 0.00165199f $X=3.77 $Y=0.995 $X2=0
+ $Y2=0
cc_285 N_A_42_47#_c_272_n N_VGND_c_703_n 0.030397f $X=0.375 $Y=0.36 $X2=0 $Y2=0
cc_286 N_A_42_47#_c_268_n N_VGND_c_708_n 0.00719299f $X=3.35 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_42_47#_c_269_n N_VGND_c_708_n 5.25906e-19 $X=3.77 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_42_47#_M1021_s N_VGND_c_710_n 0.00507005f $X=0.21 $Y=0.235 $X2=0
+ $Y2=0
cc_289 N_A_42_47#_c_268_n N_VGND_c_710_n 0.00445457f $X=3.35 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_42_47#_c_269_n N_VGND_c_710_n 0.00577464f $X=3.77 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_42_47#_c_272_n N_VGND_c_710_n 0.016639f $X=0.375 $Y=0.36 $X2=0 $Y2=0
cc_292 N_A2_c_378_n N_A1_c_451_n 0.0514295f $X=4.19 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_293 N_A2_M1015_g N_A1_M1001_g 0.0445633f $X=4.19 $Y=1.985 $X2=0 $Y2=0
cc_294 A2 N_A1_M1001_g 0.0122471f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_295 N_A2_c_379_n N_A1_c_452_n 0.0340804f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A2_M1016_g N_A1_M1011_g 0.0340804f $X=5.45 $Y=1.985 $X2=0 $Y2=0
cc_297 A2 N_A1_M1011_g 0.0149047f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_298 N_A2_c_372_n A1 0.00636853f $X=4.332 $Y=1.595 $X2=0 $Y2=0
cc_299 N_A2_c_373_n A1 0.0139635f $X=5.39 $Y=1.172 $X2=0 $Y2=0
cc_300 N_A2_c_375_n A1 4.42976e-19 $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A2_c_376_n A1 2.96815e-19 $X=4.19 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A2_c_377_n A1 0.0214745f $X=4.332 $Y=1.142 $X2=0 $Y2=0
cc_303 A2 A1 0.0224776f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_304 N_A2_c_372_n N_A1_c_453_n 0.00572537f $X=4.332 $Y=1.595 $X2=0 $Y2=0
cc_305 N_A2_c_373_n N_A1_c_453_n 0.00224079f $X=5.39 $Y=1.172 $X2=0 $Y2=0
cc_306 N_A2_c_375_n N_A1_c_453_n 0.0340804f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A2_c_376_n N_A1_c_453_n 0.0214987f $X=4.19 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A2_c_377_n N_A1_c_453_n 0.00180338f $X=4.332 $Y=1.142 $X2=0 $Y2=0
cc_309 A2 N_A1_c_453_n 0.00626189f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_310 N_A2_c_372_n N_VPWR_M1015_s 0.00122884f $X=4.332 $Y=1.595 $X2=0 $Y2=0
cc_311 N_A2_c_417_p N_VPWR_M1015_s 0.00106536f $X=4.42 $Y=1.68 $X2=0 $Y2=0
cc_312 A2 N_VPWR_M1015_s 0.00278226f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_313 A2 N_VPWR_M1011_d 0.0040068f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_314 N_A2_c_420_p N_VPWR_M1011_d 0.00107749f $X=5.305 $Y=1.595 $X2=0 $Y2=0
cc_315 N_A2_M1015_g N_VPWR_c_501_n 0.00827071f $X=4.19 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A2_M1016_g N_VPWR_c_502_n 0.0143014f $X=5.45 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A2_M1015_g N_VPWR_c_506_n 0.00337001f $X=4.19 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A2_M1016_g N_VPWR_c_508_n 0.00337001f $X=5.45 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A2_M1015_g N_VPWR_c_496_n 0.00397658f $X=4.19 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A2_M1016_g N_VPWR_c_496_n 0.00499407f $X=5.45 $Y=1.985 $X2=0 $Y2=0
cc_321 A2 N_A_603_297#_M1001_s 0.00336344f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_322 N_A2_M1015_g N_A_603_297#_c_643_n 5.08146e-19 $X=4.19 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A2_c_372_n N_A_603_297#_c_643_n 0.00626654f $X=4.332 $Y=1.595 $X2=0
+ $Y2=0
cc_324 N_A2_c_376_n N_A_603_297#_c_643_n 2.22737e-19 $X=4.19 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A2_c_377_n N_A_603_297#_c_643_n 0.00336061f $X=4.332 $Y=1.142 $X2=0
+ $Y2=0
cc_326 N_A2_M1015_g N_A_603_297#_c_644_n 0.0112565f $X=4.19 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A2_M1016_g N_A_603_297#_c_644_n 0.0112871f $X=5.45 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A2_c_374_n N_A_603_297#_c_644_n 0.00359651f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A2_c_377_n N_A_603_297#_c_644_n 0.00354175f $X=4.332 $Y=1.142 $X2=0
+ $Y2=0
cc_330 N_A2_c_417_p N_A_603_297#_c_644_n 0.00916418f $X=4.42 $Y=1.68 $X2=0 $Y2=0
cc_331 A2 N_A_603_297#_c_644_n 0.03995f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_332 N_A2_c_420_p N_A_603_297#_c_644_n 0.00906061f $X=5.305 $Y=1.595 $X2=0
+ $Y2=0
cc_333 N_A2_M1016_g N_A_603_297#_c_645_n 5.62971e-19 $X=5.45 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A2_c_374_n N_A_603_297#_c_645_n 0.0108014f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A2_c_375_n N_A_603_297#_c_645_n 0.00179227f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_336 A2 N_A_603_297#_c_645_n 0.00526012f $X=5.22 $Y=1.445 $X2=0 $Y2=0
cc_337 N_A2_c_378_n N_VGND_c_700_n 0.00902354f $X=4.19 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A2_c_374_n N_VGND_c_702_n 0.0110232f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A2_c_375_n N_VGND_c_702_n 0.00235636f $X=5.51 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A2_c_379_n N_VGND_c_702_n 0.0047742f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A2_c_378_n N_VGND_c_705_n 0.00343403f $X=4.19 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A2_c_379_n N_VGND_c_705_n 0.00585385f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A2_c_378_n N_VGND_c_710_n 0.00397751f $X=4.19 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A2_c_379_n N_VGND_c_710_n 0.011573f $X=5.51 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A1_M1001_g N_VPWR_c_501_n 0.00772604f $X=4.61 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A1_M1011_g N_VPWR_c_501_n 0.0010441f $X=5.03 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A1_M1001_g N_VPWR_c_502_n 0.0010441f $X=4.61 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A1_M1011_g N_VPWR_c_502_n 0.00772604f $X=5.03 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A1_M1001_g N_VPWR_c_507_n 0.00337001f $X=4.61 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A1_M1011_g N_VPWR_c_507_n 0.00337001f $X=5.03 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A1_M1001_g N_VPWR_c_496_n 0.00394833f $X=4.61 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A1_M1011_g N_VPWR_c_496_n 0.00394833f $X=5.03 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A1_M1001_g N_A_603_297#_c_644_n 0.00933951f $X=4.61 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A1_M1011_g N_A_603_297#_c_644_n 0.00933951f $X=5.03 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A1_c_451_n N_VGND_c_700_n 0.00206539f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A1_c_451_n N_VGND_c_705_n 0.00430182f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A1_c_452_n N_VGND_c_705_n 0.00573486f $X=5.03 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A1_c_451_n N_VGND_c_710_n 0.00588392f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A1_c_452_n N_VGND_c_710_n 0.010515f $X=5.03 $Y=0.995 $X2=0 $Y2=0
cc_360 N_VPWR_c_496_n N_X_M1006_d 0.00318969f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_361 N_VPWR_c_496_n N_X_M1010_d 0.00318969f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_362 N_VPWR_M1009_s N_X_c_618_n 0.00368438f $X=1.605 $Y=1.485 $X2=0 $Y2=0
cc_363 N_VPWR_c_496_n N_A_603_297#_M1000_d 0.00355556f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_364 N_VPWR_c_496_n N_A_603_297#_M1003_d 0.00238517f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_496_n N_A_603_297#_M1001_s 0.00307577f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_496_n N_A_603_297#_M1016_d 0.00297225f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_506_n N_A_603_297#_c_647_n 0.0230995f $X=4.235 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_496_n N_A_603_297#_c_647_n 0.0218411f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_500_n N_A_603_297#_c_682_n 0.00628485f $X=2.6 $Y=2.36 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_506_n N_A_603_297#_c_682_n 0.00755661f $X=4.235 $Y=2.72 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_496_n N_A_603_297#_c_682_n 0.00625935f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_372 N_VPWR_M1015_s N_A_603_297#_c_644_n 0.00320647f $X=4.265 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_VPWR_M1011_d N_A_603_297#_c_644_n 0.00323836f $X=5.105 $Y=1.485 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_501_n N_A_603_297#_c_644_n 0.0158599f $X=4.4 $Y=2.36 $X2=0 $Y2=0
cc_375 N_VPWR_c_502_n N_A_603_297#_c_644_n 0.0158599f $X=5.24 $Y=2.36 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_506_n N_A_603_297#_c_644_n 0.00255672f $X=4.235 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_507_n N_A_603_297#_c_644_n 0.00811322f $X=5.075 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_508_n N_A_603_297#_c_644_n 0.00755572f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_496_n N_A_603_297#_c_644_n 0.0327416f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_506_n N_A_603_297#_c_693_n 0.0075927f $X=4.235 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_496_n N_A_603_297#_c_693_n 0.00655231f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_X_c_605_n N_VGND_M1007_d 0.00338318f $X=2.175 $Y=0.7 $X2=0 $Y2=0
cc_383 N_X_c_604_n N_VGND_c_696_n 0.00184492f $X=1.235 $Y=0.7 $X2=0 $Y2=0
cc_384 N_X_c_604_n N_VGND_c_697_n 0.00298323f $X=1.235 $Y=0.7 $X2=0 $Y2=0
cc_385 N_X_c_605_n N_VGND_c_697_n 0.00569019f $X=2.175 $Y=0.7 $X2=0 $Y2=0
cc_386 N_X_c_605_n N_VGND_c_698_n 0.0159085f $X=2.175 $Y=0.7 $X2=0 $Y2=0
cc_387 N_X_c_605_n N_VGND_c_707_n 0.00676299f $X=2.175 $Y=0.7 $X2=0 $Y2=0
cc_388 N_X_M1005_s N_VGND_c_710_n 0.00318884f $X=1.175 $Y=0.235 $X2=0 $Y2=0
cc_389 N_X_M1008_s N_VGND_c_710_n 0.00318969f $X=2.035 $Y=0.235 $X2=0 $Y2=0
cc_390 N_X_c_604_n N_VGND_c_710_n 0.00528066f $X=1.235 $Y=0.7 $X2=0 $Y2=0
cc_391 N_X_c_605_n N_VGND_c_710_n 0.0224517f $X=2.175 $Y=0.7 $X2=0 $Y2=0
cc_392 N_A_603_297#_c_645_n N_VGND_c_702_n 0.00477372f $X=5.66 $Y=1.63 $X2=0
+ $Y2=0
cc_393 N_VGND_c_710_n A_861_47# 0.00280308f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_394 N_VGND_c_710_n A_1021_47# 0.0115413f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__and2_4.spice
* Created: Thu Aug 27 14:07:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2_4.pex.spice"
.subckt sky130_fd_sc_hd__and2_4  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_110_47# N_A_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.65 AD=0.138125
+ AS=0.06825 PD=1.075 PS=0.86 NRD=12.912 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.138125 PD=0.93 PS=1.075 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75001.1 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1002_d N_A_27_47#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1007_d N_A_27_47#_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1007_d N_A_27_47#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.18525 PD=0.93 PS=1.87 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_27_47#_M1006_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_B_M1010_g N_A_27_47#_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1775 AS=0.14 PD=1.355 PS=1.28 NRD=6.8753 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.1775 PD=1.28 PS=1.355 NRD=0 NRS=7.8603 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1001_d N_A_27_47#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1009_d N_A_27_47#_M1009_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1011 N_X_M1009_d N_A_27_47#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__and2_4.pxi.spice"
*
.ends
*
*

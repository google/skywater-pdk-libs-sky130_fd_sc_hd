* File: sky130_fd_sc_hd__nand2b_1.pxi.spice
* Created: Thu Aug 27 14:29:04 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2B_1%A_N N_A_N_c_44_n N_A_N_M1005_g N_A_N_M1002_g A_N
+ N_A_N_c_46_n PM_SKY130_FD_SC_HD__NAND2B_1%A_N
x_PM_SKY130_FD_SC_HD__NAND2B_1%B N_B_M1001_g N_B_M1004_g B N_B_c_71_n N_B_c_72_n
+ N_B_c_73_n PM_SKY130_FD_SC_HD__NAND2B_1%B
x_PM_SKY130_FD_SC_HD__NAND2B_1%A_27_93# N_A_27_93#_M1005_s N_A_27_93#_M1002_s
+ N_A_27_93#_M1000_g N_A_27_93#_M1003_g N_A_27_93#_c_105_n N_A_27_93#_c_119_n
+ N_A_27_93#_c_106_n N_A_27_93#_c_112_n N_A_27_93#_c_107_n N_A_27_93#_c_113_n
+ N_A_27_93#_c_108_n N_A_27_93#_c_109_n N_A_27_93#_c_110_n
+ PM_SKY130_FD_SC_HD__NAND2B_1%A_27_93#
x_PM_SKY130_FD_SC_HD__NAND2B_1%VPWR N_VPWR_M1002_d N_VPWR_M1003_d N_VPWR_c_177_n
+ N_VPWR_c_178_n VPWR N_VPWR_c_179_n N_VPWR_c_180_n N_VPWR_c_181_n
+ N_VPWR_c_176_n N_VPWR_c_183_n N_VPWR_c_184_n PM_SKY130_FD_SC_HD__NAND2B_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND2B_1%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_209_n N_Y_c_206_n
+ N_Y_c_213_n Y Y Y Y Y N_Y_c_208_n N_Y_c_211_n PM_SKY130_FD_SC_HD__NAND2B_1%Y
x_PM_SKY130_FD_SC_HD__NAND2B_1%VGND N_VGND_M1005_d N_VGND_c_249_n VGND
+ N_VGND_c_250_n N_VGND_c_251_n N_VGND_c_252_n N_VGND_c_253_n
+ PM_SKY130_FD_SC_HD__NAND2B_1%VGND
cc_1 VNB N_A_N_c_44_n 0.0236738f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A_N 0.00877746f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_46_n 0.0368982f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_c_71_n 0.022463f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_5 VNB N_B_c_72_n 0.0041123f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_6 VNB N_B_c_73_n 0.0182088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_93#_c_105_n 0.0059118f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_8 VNB N_A_27_93#_c_106_n 0.00178328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_93#_c_107_n 0.0166306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_93#_c_108_n 0.0036436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_93#_c_109_n 0.0278957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_93#_c_110_n 0.0191722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_176_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_206_n 0.00485257f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_15 VNB Y 0.0455434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_208_n 0.0184737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_249_n 0.00801986f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.695
cc_18 VNB N_VGND_c_250_n 0.0183065f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_19 VNB N_VGND_c_251_n 0.0363115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_252_n 0.152786f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_253_n 0.00507625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A_N_M1002_g 0.029585f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_23 VPB A_N 5.16752e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_24 VPB N_A_N_c_46_n 0.00895315f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_25 VPB N_B_M1004_g 0.0221673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_26 VPB N_B_c_71_n 0.00558773f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_27 VPB N_B_c_72_n 0.00147512f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_28 VPB N_A_27_93#_M1003_g 0.021892f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_29 VPB N_A_27_93#_c_112_n 0.00171533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_27_93#_c_113_n 0.0145655f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_27_93#_c_108_n 4.62603e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_93#_c_109_n 0.00698897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_177_n 0.022765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_178_n 0.00441684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_179_n 0.0206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_180_n 0.017296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_181_n 0.0190186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_176_n 0.0666901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_183_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_184_n 0.00410458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_Y_c_209_n 0.00459592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB Y 0.0323363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_Y_c_211_n 0.0146213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 N_A_N_M1002_g N_B_M1004_g 0.0220676f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_45 N_A_N_c_46_n N_B_c_71_n 0.0219809f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_46 A_N N_B_c_72_n 0.0196625f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A_N_c_46_n N_B_c_72_n 0.00178196f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_48 N_A_N_c_44_n N_B_c_73_n 0.0195264f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_N_c_44_n N_A_27_93#_c_105_n 0.0118035f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_50 A_N N_A_27_93#_c_105_n 0.00570078f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_51 N_A_N_c_46_n N_A_27_93#_c_105_n 8.62652e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_N_M1002_g N_A_27_93#_c_119_n 0.0140831f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_53 A_N N_A_27_93#_c_119_n 0.00381374f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_N_c_44_n N_A_27_93#_c_107_n 2.09932e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_55 A_N N_A_27_93#_c_107_n 0.021146f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_N_c_46_n N_A_27_93#_c_107_n 0.00627216f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_57 A_N N_A_27_93#_c_113_n 0.0192164f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_N_c_46_n N_A_27_93#_c_113_n 0.00585749f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_N_M1002_g N_VPWR_c_177_n 0.00385831f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_60 N_A_N_M1002_g N_VPWR_c_179_n 0.00327927f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_61 N_A_N_M1002_g N_VPWR_c_176_n 0.00417489f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_62 N_A_N_c_44_n N_VGND_c_249_n 0.00409614f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_N_c_44_n N_VGND_c_250_n 0.00399957f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_64 N_A_N_c_44_n N_VGND_c_252_n 0.00512902f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_65 N_B_M1004_g N_A_27_93#_M1003_g 0.0294511f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_66 N_B_c_71_n N_A_27_93#_c_105_n 0.0044365f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_72_n N_A_27_93#_c_105_n 0.034861f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B_c_73_n N_A_27_93#_c_105_n 0.0120784f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B_M1004_g N_A_27_93#_c_119_n 0.0143681f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_70 N_B_c_71_n N_A_27_93#_c_119_n 0.00268559f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B_c_72_n N_A_27_93#_c_119_n 0.0290592f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B_c_71_n N_A_27_93#_c_106_n 0.0016389f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B_c_73_n N_A_27_93#_c_106_n 0.00171329f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_74 N_B_M1004_g N_A_27_93#_c_112_n 0.00308989f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_75 N_B_c_71_n N_A_27_93#_c_108_n 0.00104254f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B_c_72_n N_A_27_93#_c_108_n 0.0197295f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B_c_71_n N_A_27_93#_c_109_n 0.0206034f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_c_72_n N_A_27_93#_c_109_n 2.71194e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B_c_73_n N_A_27_93#_c_110_n 0.041822f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_M1004_g N_VPWR_c_177_n 0.00321269f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_VPWR_c_180_n 0.00541359f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_VPWR_c_176_n 0.0108548f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_83 N_B_c_73_n N_Y_c_206_n 8.42228e-19 $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_M1004_g N_Y_c_213_n 0.00747675f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_85 N_B_c_73_n N_VGND_c_249_n 0.0118162f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B_c_73_n N_VGND_c_251_n 0.00350562f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_87 N_B_c_73_n N_VGND_c_252_n 0.00421399f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_27_93#_c_119_n N_VPWR_M1002_d 0.0046614f $X=1.255 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_27_93#_c_119_n N_VPWR_c_177_n 0.0179802f $X=1.255 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_27_93#_M1003_g N_VPWR_c_178_n 0.00319321f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A_27_93#_M1003_g N_VPWR_c_180_n 0.00422241f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A_27_93#_M1003_g N_VPWR_c_176_n 0.00704983f $X=1.375 $Y=1.985 $X2=0
+ $Y2=0
cc_93 N_A_27_93#_c_119_n N_Y_M1004_d 0.00454608f $X=1.255 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_27_93#_M1003_g N_Y_c_209_n 0.0108103f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_119_n N_Y_c_209_n 0.00676409f $X=1.255 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_27_93#_c_108_n N_Y_c_209_n 0.00534441f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_27_93#_c_109_n N_Y_c_209_n 0.00293952f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_27_93#_c_105_n N_Y_c_206_n 3.29472e-19 $X=1.255 $Y=0.82 $X2=0 $Y2=0
cc_99 N_A_27_93#_c_108_n N_Y_c_206_n 0.00534677f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_93#_c_109_n N_Y_c_206_n 0.00321342f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_27_93#_c_110_n N_Y_c_206_n 0.00597897f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_27_93#_M1003_g N_Y_c_213_n 0.011689f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_27_93#_c_119_n N_Y_c_213_n 0.017199f $X=1.255 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_27_93#_M1003_g Y 0.0112918f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_27_93#_c_105_n Y 0.00795379f $X=1.255 $Y=0.82 $X2=0 $Y2=0
cc_106 N_A_27_93#_c_119_n Y 0.00795379f $X=1.255 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A_27_93#_c_106_n Y 0.00717412f $X=1.34 $Y=1.075 $X2=0 $Y2=0
cc_108 N_A_27_93#_c_112_n Y 0.00717868f $X=1.34 $Y=1.495 $X2=0 $Y2=0
cc_109 N_A_27_93#_c_108_n Y 0.0200873f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_27_93#_c_109_n Y 0.003939f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_27_93#_c_110_n Y 0.0100732f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_27_93#_c_105_n N_VGND_M1005_d 0.00240251f $X=1.255 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_113 N_A_27_93#_c_105_n N_VGND_c_249_n 0.0176343f $X=1.255 $Y=0.82 $X2=0 $Y2=0
cc_114 N_A_27_93#_c_110_n N_VGND_c_249_n 0.00199413f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_A_27_93#_c_105_n N_VGND_c_250_n 0.00248202f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_116 N_A_27_93#_c_107_n N_VGND_c_250_n 0.00625139f $X=0.26 $Y=0.69 $X2=0 $Y2=0
cc_117 N_A_27_93#_c_105_n N_VGND_c_251_n 0.00629344f $X=1.255 $Y=0.82 $X2=0
+ $Y2=0
cc_118 N_A_27_93#_c_110_n N_VGND_c_251_n 0.00422832f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_119 N_A_27_93#_c_105_n N_VGND_c_252_n 0.0192375f $X=1.255 $Y=0.82 $X2=0 $Y2=0
cc_120 N_A_27_93#_c_107_n N_VGND_c_252_n 0.00852335f $X=0.26 $Y=0.69 $X2=0 $Y2=0
cc_121 N_A_27_93#_c_110_n N_VGND_c_252_n 0.00726488f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_27_93#_c_105_n A_206_47# 0.00302426f $X=1.255 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_123 N_VPWR_c_176_n N_Y_M1004_d 0.00215201f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_124 N_VPWR_M1003_d N_Y_c_209_n 0.00807619f $X=1.45 $Y=1.485 $X2=0 $Y2=0
cc_125 N_VPWR_c_178_n N_Y_c_209_n 0.0161606f $X=1.585 $Y=2.34 $X2=0 $Y2=0
cc_126 N_VPWR_c_180_n N_Y_c_209_n 0.0020257f $X=1.5 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_181_n N_Y_c_209_n 0.0013052f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_128 N_VPWR_c_176_n N_Y_c_209_n 0.00698115f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_180_n N_Y_c_213_n 0.0188215f $X=1.5 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_c_176_n N_Y_c_213_n 0.0121968f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_131 N_VPWR_c_181_n N_Y_c_211_n 0.00639875f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_132 N_VPWR_c_176_n N_Y_c_211_n 0.0104802f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_133 N_Y_c_206_n N_VGND_c_249_n 0.00934352f $X=1.8 $Y=0.4 $X2=0 $Y2=0
cc_134 N_Y_c_206_n N_VGND_c_251_n 0.0232267f $X=1.8 $Y=0.4 $X2=0 $Y2=0
cc_135 N_Y_c_208_n N_VGND_c_251_n 0.0265272f $X=1.985 $Y=0.545 $X2=0 $Y2=0
cc_136 N_Y_M1000_d N_VGND_c_252_n 0.00209344f $X=1.45 $Y=0.235 $X2=0 $Y2=0
cc_137 N_Y_c_206_n N_VGND_c_252_n 0.0141089f $X=1.8 $Y=0.4 $X2=0 $Y2=0
cc_138 N_Y_c_208_n N_VGND_c_252_n 0.0142494f $X=1.985 $Y=0.545 $X2=0 $Y2=0
cc_139 N_VGND_c_252_n A_206_47# 0.00354994f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24

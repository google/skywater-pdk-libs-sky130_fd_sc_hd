* File: sky130_fd_sc_hd__xor2_4.spice.pex
* Created: Thu Aug 27 14:49:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XOR2_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 58 59 60 62 63 68 71 72 84 92
c229 60 0 1.39671e-19 $X=2.8 $Y=1.53
r230 89 90 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.465 $Y=1.16
+ $X2=6.885 $Y2=1.16
r231 82 84 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.615 $Y=1.16
+ $X2=1.745 $Y2=1.16
r232 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.615
+ $Y=1.16 $X2=1.615 $Y2=1.16
r233 80 82 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.325 $Y=1.16
+ $X2=1.615 $Y2=1.16
r234 79 80 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=1.325 $Y2=1.16
r235 77 79 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.905 $Y2=1.16
r236 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r237 74 77 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.485 $Y=1.16
+ $X2=0.595 $Y2=1.16
r238 72 83 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=1.615 $Y2=1.175
r239 72 78 30.7773 $w=1.98e-07 $l=5.55e-07 $layer=LI1_cond $X=1.15 $Y=1.175
+ $X2=0.595 $Y2=1.175
r240 71 83 56.2864 $w=1.98e-07 $l=1.015e-06 $layer=LI1_cond $X=2.63 $Y=1.175
+ $X2=1.615 $Y2=1.175
r241 69 92 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.19 $Y=1.16
+ $X2=7.305 $Y2=1.16
r242 69 90 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=7.19 $Y=1.16
+ $X2=6.885 $Y2=1.16
r243 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.19
+ $Y=1.16 $X2=7.19 $Y2=1.16
r244 66 89 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=6.17 $Y=1.16
+ $X2=6.465 $Y2=1.16
r245 66 86 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.17 $Y=1.16
+ $X2=6.045 $Y2=1.16
r246 65 68 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=6.17 $Y=1.175
+ $X2=7.19 $Y2=1.175
r247 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.17
+ $Y=1.16 $X2=6.17 $Y2=1.16
r248 63 65 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=6.165 $Y=1.175
+ $X2=6.17 $Y2=1.175
r249 61 63 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=6.08 $Y=1.275
+ $X2=6.165 $Y2=1.175
r250 61 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.08 $Y=1.275
+ $X2=6.08 $Y2=1.445
r251 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.995 $Y=1.53
+ $X2=6.08 $Y2=1.445
r252 59 60 208.444 $w=1.68e-07 $l=3.195e-06 $layer=LI1_cond $X=5.995 $Y=1.53
+ $X2=2.8 $Y2=1.53
r253 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.715 $Y=1.445
+ $X2=2.8 $Y2=1.53
r254 57 71 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.715 $Y=1.275
+ $X2=2.63 $Y2=1.175
r255 57 58 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.715 $Y=1.275
+ $X2=2.715 $Y2=1.445
r256 53 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.305 $Y=1.325
+ $X2=7.305 $Y2=1.16
r257 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.305 $Y=1.325
+ $X2=7.305 $Y2=1.985
r258 50 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.305 $Y=0.995
+ $X2=7.305 $Y2=1.16
r259 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.305 $Y=0.995
+ $X2=7.305 $Y2=0.56
r260 46 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.885 $Y=1.325
+ $X2=6.885 $Y2=1.16
r261 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.885 $Y=1.325
+ $X2=6.885 $Y2=1.985
r262 43 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.885 $Y=0.995
+ $X2=6.885 $Y2=1.16
r263 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.885 $Y=0.995
+ $X2=6.885 $Y2=0.56
r264 39 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.325
+ $X2=6.465 $Y2=1.16
r265 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.465 $Y=1.325
+ $X2=6.465 $Y2=1.985
r266 36 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=0.995
+ $X2=6.465 $Y2=1.16
r267 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.465 $Y=0.995
+ $X2=6.465 $Y2=0.56
r268 32 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=1.325
+ $X2=6.045 $Y2=1.16
r269 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.045 $Y=1.325
+ $X2=6.045 $Y2=1.985
r270 29 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.045 $Y=0.995
+ $X2=6.045 $Y2=1.16
r271 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.045 $Y=0.995
+ $X2=6.045 $Y2=0.56
r272 25 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.16
r273 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.985
r274 22 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=1.16
r275 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=0.56
r276 18 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.16
r277 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.985
r278 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=1.16
r279 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=0.56
r280 11 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r281 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r282 8 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r283 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r284 4 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r285 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.985
r286 1 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r287 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 33
+ 36 38 40 43 45 47 50 52 54 57 63 77 79
c154 13 0 1.56361e-19 $X=2.585 $Y=1.985
r155 78 79 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.205 $Y=1.16
+ $X2=5.625 $Y2=1.16
r156 76 78 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=4.835 $Y=1.16
+ $X2=5.205 $Y2=1.16
r157 76 77 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.835
+ $Y=1.16 $X2=4.835 $Y2=1.16
r158 74 76 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.785 $Y=1.16
+ $X2=4.835 $Y2=1.16
r159 73 74 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.365 $Y=1.16
+ $X2=4.785 $Y2=1.16
r160 70 72 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.135 $Y=1.16
+ $X2=3.425 $Y2=1.16
r161 70 71 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.135
+ $Y=1.16 $X2=3.135 $Y2=1.16
r162 68 70 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=3.005 $Y=1.16
+ $X2=3.135 $Y2=1.16
r163 67 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.585 $Y=1.16
+ $X2=3.005 $Y2=1.16
r164 65 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.165 $Y=1.16
+ $X2=2.585 $Y2=1.16
r165 63 77 51.2955 $w=1.98e-07 $l=9.25e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=4.835 $Y2=1.175
r166 63 71 42.9773 $w=1.98e-07 $l=7.75e-07 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.135 $Y2=1.175
r167 55 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=1.325
+ $X2=5.625 $Y2=1.16
r168 55 57 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.625 $Y=1.325
+ $X2=5.625 $Y2=1.985
r169 52 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=0.995
+ $X2=5.625 $Y2=1.16
r170 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.625 $Y=0.995
+ $X2=5.625 $Y2=0.56
r171 48 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.325
+ $X2=5.205 $Y2=1.16
r172 48 50 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.205 $Y=1.325
+ $X2=5.205 $Y2=1.985
r173 45 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=0.995
+ $X2=5.205 $Y2=1.16
r174 45 47 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.205 $Y=0.995
+ $X2=5.205 $Y2=0.56
r175 41 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=1.325
+ $X2=4.785 $Y2=1.16
r176 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.785 $Y=1.325
+ $X2=4.785 $Y2=1.985
r177 38 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.785 $Y=0.995
+ $X2=4.785 $Y2=1.16
r178 38 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.785 $Y=0.995
+ $X2=4.785 $Y2=0.56
r179 34 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.325
+ $X2=4.365 $Y2=1.16
r180 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.365 $Y=1.325
+ $X2=4.365 $Y2=1.985
r181 31 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.365 $Y2=1.16
r182 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.365 $Y2=0.56
r183 30 72 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.5 $Y=1.16
+ $X2=3.425 $Y2=1.16
r184 29 73 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=1.16
+ $X2=4.365 $Y2=1.16
r185 29 30 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=4.29 $Y=1.16 $X2=3.5
+ $Y2=1.16
r186 25 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.325
+ $X2=3.425 $Y2=1.16
r187 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.425 $Y=1.325
+ $X2=3.425 $Y2=1.985
r188 22 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.16
r189 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=0.56
r190 18 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.005 $Y=1.325
+ $X2=3.005 $Y2=1.16
r191 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.005 $Y=1.325
+ $X2=3.005 $Y2=1.985
r192 15 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=1.16
r193 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=0.56
r194 11 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.325
+ $X2=2.585 $Y2=1.16
r195 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.585 $Y=1.325
+ $X2=2.585 $Y2=1.985
r196 8 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.585 $Y2=1.16
r197 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.585 $Y=0.995
+ $X2=2.585 $Y2=0.56
r198 4 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.16
r199 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.165 $Y=1.325
+ $X2=2.165 $Y2=1.985
r200 1 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=1.16
r201 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.165 $Y=0.995
+ $X2=2.165 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%A_112_47# 1 2 3 4 5 6 19 21 24 26 28 31 33 35
+ 38 40 42 45 48 49 50 53 55 59 61 65 69 71 75 80 82 83 88 91 92 93 94 95 96 97
+ 101 106 107 108 114 115 123
c271 108 0 2.96032e-19 $X=2.215 $Y=1.53
c272 107 0 4.26736e-19 $X=7.445 $Y=1.53
c273 33 0 2.9244e-20 $X=9.095 $Y=0.995
c274 26 0 1.37821e-19 $X=8.675 $Y=0.995
r275 117 119 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.255 $Y=1.16
+ $X2=8.675 $Y2=1.16
r276 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=1.53
+ $X2=7.59 $Y2=1.53
r277 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=1.53
+ $X2=2.07 $Y2=1.53
r278 108 110 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=1.53
+ $X2=2.07 $Y2=1.53
r279 107 114 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=1.53
+ $X2=7.59 $Y2=1.53
r280 107 108 6.47276 $w=1.4e-07 $l=5.23e-06 $layer=MET1_cond $X=7.445 $Y=1.53
+ $X2=2.215 $Y2=1.53
r281 101 104 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.215 $Y=1.87
+ $X2=3.215 $Y2=1.96
r282 96 99 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.375 $Y=1.87
+ $X2=2.375 $Y2=1.96
r283 96 97 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=1.87
+ $X2=2.375 $Y2=1.785
r284 95 111 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=1.53
+ $X2=2.07 $Y2=1.53
r285 91 111 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=0.255 $Y=1.53
+ $X2=2.07 $Y2=1.53
r286 89 123 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=9.385 $Y=1.16
+ $X2=9.515 $Y2=1.16
r287 89 121 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=9.385 $Y=1.16
+ $X2=9.095 $Y2=1.16
r288 88 89 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.385
+ $Y=1.16 $X2=9.385 $Y2=1.16
r289 86 121 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=8.705 $Y=1.16
+ $X2=9.095 $Y2=1.16
r290 86 119 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.705 $Y=1.16
+ $X2=8.675 $Y2=1.16
r291 85 88 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=8.705 $Y=1.175
+ $X2=9.385 $Y2=1.175
r292 85 86 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=1.16 $X2=8.705 $Y2=1.16
r293 83 106 5.8268 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=8.64 $Y=1.175
+ $X2=8.54 $Y2=1.175
r294 83 85 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=8.64 $Y=1.175
+ $X2=8.705 $Y2=1.175
r295 82 106 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=7.71 $Y=1.19
+ $X2=8.54 $Y2=1.19
r296 80 115 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.625 $Y=1.445
+ $X2=7.625 $Y2=1.53
r297 79 82 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.625 $Y=1.275
+ $X2=7.71 $Y2=1.19
r298 79 80 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.625 $Y=1.275
+ $X2=7.625 $Y2=1.445
r299 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.215 $Y=0.725
+ $X2=3.215 $Y2=0.39
r300 72 94 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0.815
+ $X2=2.375 $Y2=0.815
r301 71 73 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.05 $Y=0.815
+ $X2=3.215 $Y2=0.725
r302 71 72 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.05 $Y=0.815
+ $X2=2.54 $Y2=0.815
r303 70 96 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.5 $Y=1.87
+ $X2=2.375 $Y2=1.87
r304 69 101 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=1.87
+ $X2=3.215 $Y2=1.87
r305 69 70 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.09 $Y=1.87 $X2=2.5
+ $Y2=1.87
r306 67 95 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=1.615
+ $X2=2.25 $Y2=1.53
r307 67 97 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.335 $Y=1.615
+ $X2=2.335 $Y2=1.785
r308 63 94 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.375 $Y=0.725
+ $X2=2.375 $Y2=0.815
r309 63 65 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.375 $Y=0.725
+ $X2=2.375 $Y2=0.39
r310 62 93 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=0.815
+ $X2=1.535 $Y2=0.815
r311 61 94 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0.815
+ $X2=2.375 $Y2=0.815
r312 61 62 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.21 $Y=0.815
+ $X2=1.7 $Y2=0.815
r313 57 93 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.535 $Y=0.725
+ $X2=1.535 $Y2=0.815
r314 57 59 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0.725
+ $X2=1.535 $Y2=0.39
r315 56 92 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=0.815
+ $X2=0.695 $Y2=0.815
r316 55 93 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0.815
+ $X2=1.535 $Y2=0.815
r317 55 56 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.37 $Y=0.815
+ $X2=0.86 $Y2=0.815
r318 51 92 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.695 $Y=0.725
+ $X2=0.695 $Y2=0.815
r319 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.695 $Y=0.725
+ $X2=0.695 $Y2=0.39
r320 49 92 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.53 $Y=0.82
+ $X2=0.695 $Y2=0.815
r321 49 50 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.53 $Y=0.82
+ $X2=0.255 $Y2=0.82
r322 48 91 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.445
+ $X2=0.255 $Y2=1.53
r323 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.255 $Y2=0.82
r324 47 48 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.17 $Y2=1.445
r325 43 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.515 $Y=1.325
+ $X2=9.515 $Y2=1.16
r326 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.515 $Y=1.325
+ $X2=9.515 $Y2=1.985
r327 40 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.515 $Y=0.995
+ $X2=9.515 $Y2=1.16
r328 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.515 $Y=0.995
+ $X2=9.515 $Y2=0.56
r329 36 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.095 $Y=1.325
+ $X2=9.095 $Y2=1.16
r330 36 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.095 $Y=1.325
+ $X2=9.095 $Y2=1.985
r331 33 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.095 $Y=0.995
+ $X2=9.095 $Y2=1.16
r332 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.095 $Y=0.995
+ $X2=9.095 $Y2=0.56
r333 29 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.325
+ $X2=8.675 $Y2=1.16
r334 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.675 $Y=1.325
+ $X2=8.675 $Y2=1.985
r335 26 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=0.995
+ $X2=8.675 $Y2=1.16
r336 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.675 $Y=0.995
+ $X2=8.675 $Y2=0.56
r337 22 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.255 $Y=1.325
+ $X2=8.255 $Y2=1.16
r338 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.255 $Y=1.325
+ $X2=8.255 $Y2=1.985
r339 19 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.255 $Y=0.995
+ $X2=8.255 $Y2=1.16
r340 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.255 $Y=0.995
+ $X2=8.255 $Y2=0.56
r341 6 104 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.215 $Y2=1.96
r342 5 99 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.485 $X2=2.375 $Y2=1.96
r343 4 75 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.235 $X2=3.215 $Y2=0.39
r344 3 65 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.39
r345 2 59 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.4
+ $Y=0.235 $X2=1.535 $Y2=0.39
r346 1 53 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.695 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%A_27_297# 1 2 3 4 5 18 22 24 26 27 28 32 35
+ 37 41
r64 41 43 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.795 $Y=2.3 $X2=2.795
+ $Y2=2.38
r65 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.635 $Y=2.295
+ $X2=3.635 $Y2=1.96
r66 29 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.92 $Y=2.38
+ $X2=2.795 $Y2=2.38
r67 28 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.51 $Y=2.38
+ $X2=3.635 $Y2=2.295
r68 28 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.51 $Y=2.38 $X2=2.92
+ $Y2=2.38
r69 26 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.67 $Y=2.38
+ $X2=2.795 $Y2=2.38
r70 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.67 $Y=2.38 $X2=2.08
+ $Y2=2.38
r71 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.955 $Y=2.295
+ $X2=2.08 $Y2=2.38
r72 24 39 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.955 $Y=2.005
+ $X2=1.955 $Y2=1.895
r73 24 25 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.955 $Y=2.005
+ $X2=1.955 $Y2=2.295
r74 23 37 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.24 $Y=1.895
+ $X2=1.115 $Y2=1.895
r75 22 39 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=1.895
+ $X2=1.955 $Y2=1.895
r76 22 23 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=1.83 $Y=1.895
+ $X2=1.24 $Y2=1.895
r77 19 35 4.18571 $w=2.2e-07 $l=1.58e-07 $layer=LI1_cond $X=0.4 $Y=1.895
+ $X2=0.242 $Y2=1.895
r78 18 37 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.99 $Y=1.895
+ $X2=1.115 $Y2=1.895
r79 18 19 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=0.99 $Y=1.895
+ $X2=0.4 $Y2=1.895
r80 5 32 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.5
+ $Y=1.485 $X2=3.635 $Y2=1.96
r81 4 41 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.485 $X2=2.795 $Y2=2.3
r82 3 39 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.82
+ $Y=1.485 $X2=1.955 $Y2=1.96
r83 2 37 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.115 $Y2=1.96
r84 1 35 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 37 41 45 47
+ 48 49 51 56 65 75 76 79 82 85 88 91
r157 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r158 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r159 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r160 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r161 82 83 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r162 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r163 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r164 73 76 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r165 73 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r166 72 75 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r167 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r168 70 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.22 $Y=2.72
+ $X2=7.095 $Y2=2.72
r169 70 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.22 $Y=2.72
+ $X2=7.59 $Y2=2.72
r170 69 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r171 69 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r172 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r173 66 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.38 $Y=2.72
+ $X2=6.255 $Y2=2.72
r174 66 68 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.38 $Y=2.72
+ $X2=6.67 $Y2=2.72
r175 65 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.97 $Y=2.72
+ $X2=7.095 $Y2=2.72
r176 65 68 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.97 $Y=2.72 $X2=6.67
+ $Y2=2.72
r177 64 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r178 64 83 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=1.61 $Y2=2.72
r179 63 64 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r180 61 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.66 $Y=2.72
+ $X2=1.535 $Y2=2.72
r181 61 63 176.802 $w=1.68e-07 $l=2.71e-06 $layer=LI1_cond $X=1.66 $Y=2.72
+ $X2=4.37 $Y2=2.72
r182 60 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r183 60 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r185 57 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=0.695 $Y2=2.72
r186 57 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=1.15 $Y2=2.72
r187 56 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.535 $Y2=2.72
r188 56 59 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r189 51 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.695 $Y2=2.72
r190 51 53 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.23 $Y2=2.72
r191 49 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r192 49 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r193 47 63 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.45 $Y=2.72 $X2=4.37
+ $Y2=2.72
r194 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.45 $Y=2.72
+ $X2=4.575 $Y2=2.72
r195 43 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=2.635
+ $X2=7.095 $Y2=2.72
r196 43 45 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.095 $Y=2.635
+ $X2=7.095 $Y2=2.34
r197 39 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.635
+ $X2=6.255 $Y2=2.72
r198 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.255 $Y=2.635
+ $X2=6.255 $Y2=2.34
r199 38 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.54 $Y=2.72
+ $X2=5.415 $Y2=2.72
r200 37 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.13 $Y=2.72
+ $X2=6.255 $Y2=2.72
r201 37 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.13 $Y=2.72
+ $X2=5.54 $Y2=2.72
r202 33 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=2.635
+ $X2=5.415 $Y2=2.72
r203 33 35 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.415 $Y=2.635
+ $X2=5.415 $Y2=2.34
r204 32 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.7 $Y=2.72
+ $X2=4.575 $Y2=2.72
r205 31 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=5.415 $Y2=2.72
r206 31 32 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.29 $Y=2.72 $X2=4.7
+ $Y2=2.72
r207 27 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=2.635
+ $X2=4.575 $Y2=2.72
r208 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.575 $Y=2.635
+ $X2=4.575 $Y2=2.34
r209 23 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.635
+ $X2=1.535 $Y2=2.72
r210 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.535 $Y=2.635
+ $X2=1.535 $Y2=2.34
r211 19 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r212 19 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.34
r213 6 45 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.96
+ $Y=1.485 $X2=7.095 $Y2=2.34
r214 5 41 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.12
+ $Y=1.485 $X2=6.255 $Y2=2.34
r215 4 35 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.485 $X2=5.415 $Y2=2.34
r216 3 29 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.485 $X2=4.575 $Y2=2.34
r217 2 25 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=1.485 $X2=1.535 $Y2=2.34
r218 1 21 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.695 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%A_806_297# 1 2 3 4 5 6 7 24 28 32 36 40 42 43
+ 44 45 48 50 54 57 59 61 63 66
c109 4 0 1.28384e-19 $X=6.54 $Y=1.485
r110 52 54 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.305 $Y=2.295
+ $X2=9.305 $Y2=1.96
r111 51 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.59 $Y=2.38
+ $X2=8.465 $Y2=2.38
r112 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.18 $Y=2.38
+ $X2=9.305 $Y2=2.295
r113 50 51 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.18 $Y=2.38
+ $X2=8.59 $Y2=2.38
r114 46 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=2.295
+ $X2=8.465 $Y2=2.38
r115 46 48 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.465 $Y=2.295
+ $X2=8.465 $Y2=2
r116 44 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.34 $Y=2.38
+ $X2=8.465 $Y2=2.38
r117 44 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.34 $Y=2.38 $X2=7.64
+ $Y2=2.38
r118 43 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.515 $Y=2.295
+ $X2=7.64 $Y2=2.38
r119 42 65 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=7.515 $Y=2.005
+ $X2=7.515 $Y2=1.895
r120 42 43 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=7.515 $Y=2.005
+ $X2=7.515 $Y2=2.295
r121 41 63 6.93182 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.8 $Y=1.895
+ $X2=6.675 $Y2=1.895
r122 40 65 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=7.39 $Y=1.895
+ $X2=7.515 $Y2=1.895
r123 40 41 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=7.39 $Y=1.895
+ $X2=6.8 $Y2=1.895
r124 34 63 5.368 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=6.675 $Y=1.785
+ $X2=6.675 $Y2=1.895
r125 34 36 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=1.785
+ $X2=6.675 $Y2=1.62
r126 33 61 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=1.895
+ $X2=5.835 $Y2=1.895
r127 32 63 6.93182 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=1.895
+ $X2=6.675 $Y2=1.895
r128 32 33 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=6.55 $Y=1.895
+ $X2=5.96 $Y2=1.895
r129 29 59 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.12 $Y=1.895
+ $X2=4.995 $Y2=1.895
r130 28 61 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.71 $Y=1.895
+ $X2=5.835 $Y2=1.895
r131 28 29 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=5.71 $Y=1.895
+ $X2=5.12 $Y2=1.895
r132 25 57 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.28 $Y=1.895
+ $X2=4.155 $Y2=1.895
r133 24 59 5.73815 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.87 $Y=1.895
+ $X2=4.995 $Y2=1.895
r134 24 25 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=4.87 $Y=1.895
+ $X2=4.28 $Y2=1.895
r135 7 54 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.17
+ $Y=1.485 $X2=9.305 $Y2=1.96
r136 6 48 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.33
+ $Y=1.485 $X2=8.465 $Y2=2
r137 5 65 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.38
+ $Y=1.485 $X2=7.515 $Y2=1.96
r138 4 63 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.54
+ $Y=1.485 $X2=6.675 $Y2=1.96
r139 4 36 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.485 $X2=6.675 $Y2=1.62
r140 3 61 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.7
+ $Y=1.485 $X2=5.835 $Y2=1.96
r141 2 59 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.86
+ $Y=1.485 $X2=4.995 $Y2=1.96
r142 1 57 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.485 $X2=4.155 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%X 1 2 3 4 5 6 7 26 28 30 34 36 40 44 46 49 52
+ 53 55 56 59 60 62 63 66 69 75
c162 69 0 1.37821e-19 $X=8.05 $Y=0.85
c163 53 0 2.9244e-20 $X=8.3 $Y=0.725
r164 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0.85
+ $X2=8.05 $Y2=0.85
r165 66 75 5.71274 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=5.29 $Y=0.79
+ $X2=5.15 $Y2=0.79
r166 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.85
r167 63 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=0.85
+ $X2=5.29 $Y2=0.85
r168 62 69 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.905 $Y=0.85
+ $X2=8.05 $Y2=0.85
r169 62 63 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=7.905 $Y=0.85
+ $X2=5.435 $Y2=0.85
r170 60 81 11.392 $w=4.33e-07 $l=4.3e-07 $layer=LI1_cond $X=9.817 $Y=1.87
+ $X2=9.817 $Y2=2.3
r171 57 60 6.49077 $w=4.33e-07 $l=2.45e-07 $layer=LI1_cond $X=9.817 $Y=1.625
+ $X2=9.817 $Y2=1.87
r172 57 59 2.75712 $w=3.67e-07 $l=9e-08 $layer=LI1_cond $X=9.817 $Y=1.625
+ $X2=9.817 $Y2=1.535
r173 52 70 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=8.3 $Y=0.83
+ $X2=8.05 $Y2=0.83
r174 52 53 7.95398 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=8.3 $Y=0.83 $X2=8.3
+ $Y2=0.725
r175 49 59 2.75712 $w=3.67e-07 $l=1.19248e-07 $layer=LI1_cond $X=9.885 $Y=1.445
+ $X2=9.817 $Y2=1.535
r176 48 49 20.744 $w=2.98e-07 $l=5.4e-07 $layer=LI1_cond $X=9.885 $Y=0.905
+ $X2=9.885 $Y2=1.445
r177 47 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=0.82
+ $X2=9.305 $Y2=0.82
r178 46 48 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=9.735 $Y=0.82
+ $X2=9.885 $Y2=0.905
r179 46 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.735 $Y=0.82
+ $X2=9.47 $Y2=0.82
r180 42 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=0.735
+ $X2=9.305 $Y2=0.82
r181 42 44 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.305 $Y=0.735
+ $X2=9.305 $Y2=0.39
r182 41 55 6.19399 $w=2e-07 $l=1.34629e-07 $layer=LI1_cond $X=9.01 $Y=1.535
+ $X2=8.885 $Y2=1.555
r183 40 59 4.00159 $w=1.8e-07 $l=2.17e-07 $layer=LI1_cond $X=9.6 $Y=1.535
+ $X2=9.817 $Y2=1.535
r184 40 41 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=9.6 $Y=1.535
+ $X2=9.01 $Y2=1.535
r185 37 53 7.95398 $w=1.9e-07 $l=3.745e-07 $layer=LI1_cond $X=8.63 $Y=0.82
+ $X2=8.3 $Y2=0.725
r186 36 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.14 $Y=0.82
+ $X2=9.305 $Y2=0.82
r187 36 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.14 $Y=0.82
+ $X2=8.63 $Y2=0.82
r188 32 53 0.546715 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.465 $Y=0.725
+ $X2=8.3 $Y2=0.725
r189 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.465 $Y=0.725
+ $X2=8.465 $Y2=0.39
r190 31 51 3.97178 $w=2.2e-07 $l=1.45e-07 $layer=LI1_cond $X=8.17 $Y=1.555
+ $X2=8.025 $Y2=1.555
r191 30 55 6.19399 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.76 $Y=1.555
+ $X2=8.885 $Y2=1.555
r192 30 31 30.9064 $w=2.18e-07 $l=5.9e-07 $layer=LI1_cond $X=8.76 $Y=1.555
+ $X2=8.17 $Y2=1.555
r193 26 51 3.01307 $w=2.9e-07 $l=1.1e-07 $layer=LI1_cond $X=8.025 $Y=1.665
+ $X2=8.025 $Y2=1.555
r194 26 28 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.025 $Y=1.665
+ $X2=8.025 $Y2=1.96
r195 24 75 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=4.575 $Y=0.775
+ $X2=5.15 $Y2=0.775
r196 7 81 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=1.485 $X2=9.725 $Y2=2.3
r197 7 59 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=1.485 $X2=9.725 $Y2=1.62
r198 6 55 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=8.75
+ $Y=1.485 $X2=8.885 $Y2=1.62
r199 5 51 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.9
+ $Y=1.485 $X2=8.045 $Y2=1.61
r200 5 28 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=7.9
+ $Y=1.485 $X2=8.045 $Y2=1.96
r201 4 44 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.17
+ $Y=0.235 $X2=9.305 $Y2=0.39
r202 3 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.33
+ $Y=0.235 $X2=8.465 $Y2=0.39
r203 2 66 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.28
+ $Y=0.235 $X2=5.415 $Y2=0.73
r204 1 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.235 $X2=4.575 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%VGND 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 53 57 61 65 69 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 95 110 128 129
+ 135
r181 135 136 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r182 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r183 126 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r184 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r185 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r186 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r187 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r188 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r189 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r190 117 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r191 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r192 114 135 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.255 $Y2=0
r193 114 116 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=0
+ $X2=6.67 $Y2=0
r194 113 136 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=6.21 $Y2=0
r195 112 113 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r196 110 135 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=6.255 $Y2=0
r197 110 112 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=3.91 $Y2=0
r198 109 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r199 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r200 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r201 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r202 103 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r203 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r204 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r205 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r206 97 132 4.29305 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r207 97 99 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.69
+ $Y2=0
r208 95 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r209 95 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r210 93 125 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.64 $Y=0 $X2=9.43
+ $Y2=0
r211 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.64 $Y=0 $X2=9.725
+ $Y2=0
r212 92 128 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=9.81 $Y=0 $X2=9.89
+ $Y2=0
r213 92 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=0 $X2=9.725
+ $Y2=0
r214 90 122 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.8 $Y=0 $X2=8.51
+ $Y2=0
r215 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.8 $Y=0 $X2=8.885
+ $Y2=0
r216 89 125 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.97 $Y=0 $X2=9.43
+ $Y2=0
r217 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=0 $X2=8.885
+ $Y2=0
r218 87 119 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.96 $Y=0 $X2=7.59
+ $Y2=0
r219 87 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=0 $X2=8.045
+ $Y2=0
r220 86 122 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.13 $Y=0 $X2=8.51
+ $Y2=0
r221 86 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.13 $Y=0 $X2=8.045
+ $Y2=0
r222 84 116 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=0 $X2=6.67
+ $Y2=0
r223 84 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0 $X2=7.095
+ $Y2=0
r224 83 119 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.18 $Y=0 $X2=7.59
+ $Y2=0
r225 83 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0 $X2=7.095
+ $Y2=0
r226 81 108 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.45
+ $Y2=0
r227 81 82 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.685
+ $Y2=0
r228 80 112 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.91
+ $Y2=0
r229 80 82 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.685
+ $Y2=0
r230 78 105 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r231 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.795
+ $Y2=0
r232 77 108 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.45
+ $Y2=0
r233 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.795
+ $Y2=0
r234 75 102 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.61
+ $Y2=0
r235 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.955
+ $Y2=0
r236 74 105 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.53
+ $Y2=0
r237 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.955
+ $Y2=0
r238 72 99 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.69
+ $Y2=0
r239 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.115
+ $Y2=0
r240 71 102 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.61
+ $Y2=0
r241 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.115
+ $Y2=0
r242 67 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.725 $Y=0.085
+ $X2=9.725 $Y2=0
r243 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.725 $Y=0.085
+ $X2=9.725 $Y2=0.39
r244 63 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0.085
+ $X2=8.885 $Y2=0
r245 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.885 $Y=0.085
+ $X2=8.885 $Y2=0.39
r246 59 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=0.085
+ $X2=8.045 $Y2=0
r247 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.045 $Y=0.085
+ $X2=8.045 $Y2=0.39
r248 55 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0
r249 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0.39
r250 51 135 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0
r251 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0.39
r252 47 82 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r253 47 49 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.39
r254 43 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0
r255 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0.39
r256 39 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0
r257 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.955 $Y=0.085
+ $X2=1.955 $Y2=0.39
r258 35 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r259 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.39
r260 31 132 3.02899 $w=2.75e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.18 $Y2=0
r261 31 33 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.222 $Y2=0.39
r262 10 69 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.59
+ $Y=0.235 $X2=9.725 $Y2=0.39
r263 9 65 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.235 $X2=8.885 $Y2=0.39
r264 8 61 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=7.92
+ $Y=0.235 $X2=8.045 $Y2=0.39
r265 7 57 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.96
+ $Y=0.235 $X2=7.095 $Y2=0.39
r266 6 53 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.235 $X2=6.255 $Y2=0.39
r267 5 49 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.235 $X2=3.635 $Y2=0.39
r268 4 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.235 $X2=2.795 $Y2=0.39
r269 3 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.235 $X2=1.955 $Y2=0.39
r270 2 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.115 $Y2=0.39
r271 1 33 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XOR2_4%A_806_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
c85 30 0 1.16143e-19 $X=7.35 $Y=0.815
c86 24 0 1.82209e-19 $X=6.51 $Y=0.815
r87 32 34 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.515 $Y=0.725
+ $X2=7.515 $Y2=0.39
r88 31 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=0.815
+ $X2=6.675 $Y2=0.815
r89 30 32 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=7.35 $Y=0.815
+ $X2=7.515 $Y2=0.725
r90 30 31 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.35 $Y=0.815
+ $X2=6.84 $Y2=0.815
r91 26 40 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.675 $Y=0.725
+ $X2=6.675 $Y2=0.815
r92 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.675 $Y=0.725
+ $X2=6.675 $Y2=0.39
r93 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=6 $Y=0.815 $X2=5.875
+ $Y2=0.815
r94 24 40 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.51 $Y=0.815
+ $X2=6.675 $Y2=0.815
r95 24 25 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.51 $Y=0.815 $X2=6
+ $Y2=0.815
r96 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.875 $Y=0.725
+ $X2=5.875 $Y2=0.815
r97 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=5.875 $Y=0.475
+ $X2=5.875 $Y2=0.365
r98 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.875 $Y=0.475
+ $X2=5.875 $Y2=0.725
r99 18 21 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=4.155 $Y=0.365
+ $X2=4.995 $Y2=0.365
r100 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=5.75 $Y=0.365
+ $X2=5.875 $Y2=0.365
r101 16 21 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=5.75 $Y=0.365
+ $X2=4.995 $Y2=0.365
r102 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.38
+ $Y=0.235 $X2=7.515 $Y2=0.39
r103 4 28 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.54
+ $Y=0.235 $X2=6.675 $Y2=0.39
r104 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.235 $X2=5.835 $Y2=0.73
r105 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.235 $X2=5.835 $Y2=0.39
r106 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.235 $X2=4.995 $Y2=0.39
r107 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.235 $X2=4.155 $Y2=0.39
.ends


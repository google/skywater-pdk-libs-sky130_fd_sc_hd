* File: sky130_fd_sc_hd__maj3_1.pex.spice
* Created: Thu Aug 27 14:27:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MAJ3_1%A 3 7 11 15 17 18 19 20 29 30
c45 11 0 7.04413e-20 $X=1.25 $Y=0.445
r46 28 30 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.04 $Y=1.16
+ $X2=1.25 $Y2=1.16
r47 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.16 $X2=1.04 $Y2=1.16
r48 25 28 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.83 $Y=1.16
+ $X2=1.04 $Y2=1.16
r49 19 20 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=1.87
+ $X2=0.695 $Y2=2.21
r50 18 19 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.87
r51 18 32 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.325
r52 17 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=1.04 $Y2=1.16
r53 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.695 $Y2=1.325
r54 13 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.325
+ $X2=1.25 $Y2=1.16
r55 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.25 $Y=1.325
+ $X2=1.25 $Y2=1.915
r56 9 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=0.995
+ $X2=1.25 $Y2=1.16
r57 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.25 $Y=0.995
+ $X2=1.25 $Y2=0.445
r58 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.83 $Y=1.325
+ $X2=0.83 $Y2=1.16
r59 5 7 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.83 $Y=1.325 $X2=0.83
+ $Y2=1.915
r60 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.83 $Y=0.995
+ $X2=0.83 $Y2=1.16
r61 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.83 $Y=0.995 $X2=0.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%B 3 7 11 15 17 18 25 26
c49 7 0 1.27656e-19 $X=1.61 $Y=1.915
r50 24 26 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=2.03 $Y2=1.16
r51 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.16 $X2=1.82 $Y2=1.16
r52 21 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.61 $Y=1.16
+ $X2=1.82 $Y2=1.16
r53 17 18 9.67483 $w=4.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.702 $Y=1.19
+ $X2=1.702 $Y2=1.53
r54 17 25 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=1.702 $Y=1.19
+ $X2=1.702 $Y2=1.16
r55 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.325
+ $X2=2.03 $Y2=1.16
r56 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.03 $Y=1.325
+ $X2=2.03 $Y2=1.915
r57 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=0.995
+ $X2=2.03 $Y2=1.16
r58 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.03 $Y=0.995
+ $X2=2.03 $Y2=0.445
r59 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.325
+ $X2=1.61 $Y2=1.16
r60 5 7 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.61 $Y=1.325 $X2=1.61
+ $Y2=1.915
r61 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.61 $Y2=1.16
r62 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.61 $Y=0.995 $X2=1.61
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%C 3 6 7 8 11 16 17 18 24
r62 21 24 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.39 $Y=1.16
+ $X2=2.575 $Y2=1.16
r63 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.575
+ $Y=1.16 $X2=2.575 $Y2=1.16
r64 17 18 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=2.585 $Y=0.85
+ $X2=2.585 $Y2=1.16
r65 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.39 $Y=2.465
+ $X2=2.39 $Y2=1.915
r66 13 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=1.325
+ $X2=2.39 $Y2=1.16
r67 13 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.39 $Y=1.325
+ $X2=2.39 $Y2=1.915
r68 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.39 $Y=0.995
+ $X2=2.39 $Y2=1.16
r69 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.39 $Y=0.995
+ $X2=2.39 $Y2=0.445
r70 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=2.54
+ $X2=2.39 $Y2=2.465
r71 7 8 907.596 $w=1.5e-07 $l=1.77e-06 $layer=POLY_cond $X=2.315 $Y=2.54
+ $X2=0.545 $Y2=2.54
r72 3 6 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=1.915
r73 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.47 $Y=2.465
+ $X2=0.545 $Y2=2.54
r74 1 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=2.465 $X2=0.47
+ $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%A_27_47# 1 2 3 4 15 18 22 26 32 34 39 41 42
+ 45 46 48 49 51 55 56 59
c109 55 0 1.84181e-19 $X=3.115 $Y=1.16
c110 49 0 7.04413e-20 $X=2.16 $Y=0.732
c111 45 0 1.33802e-19 $X=3.01 $Y=1.495
c112 39 0 1.27656e-19 $X=2.16 $Y=1.495
r113 56 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.16
+ $X2=3.115 $Y2=1.325
r114 56 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.16
+ $X2=3.115 $Y2=0.995
r115 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.16 $X2=3.115 $Y2=1.16
r116 52 55 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.01 $Y=1.16
+ $X2=3.115 $Y2=1.16
r117 44 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r118 44 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.495
r119 43 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=1.58
+ $X2=2.16 $Y2=1.58
r120 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=3.01 $Y2=1.495
r121 42 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=2.245 $Y2=1.58
r122 40 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.58
r123 40 41 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.815
r124 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=1.495
+ $X2=2.16 $Y2=1.58
r125 38 49 1.22693 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=2.16 $Y=0.825
+ $X2=2.16 $Y2=0.732
r126 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=0.825
+ $X2=2.16 $Y2=1.495
r127 34 41 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.075 $Y=1.947
+ $X2=2.16 $Y2=1.815
r128 34 36 11.0895 $w=2.63e-07 $l=2.55e-07 $layer=LI1_cond $X=2.075 $Y=1.947
+ $X2=1.82 $Y2=1.947
r129 30 49 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.82 $Y=0.732
+ $X2=2.16 $Y2=0.732
r130 30 48 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0.732
+ $X2=1.655 $Y2=0.732
r131 30 32 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.82 $Y=0.64
+ $X2=1.82 $Y2=0.445
r132 29 46 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.395 $Y=0.74
+ $X2=0.265 $Y2=0.74
r133 29 48 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=0.395 $Y=0.74
+ $X2=1.655 $Y2=0.74
r134 24 46 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=0.825
+ $X2=0.265 $Y2=0.74
r135 24 26 48.314 $w=2.58e-07 $l=1.09e-06 $layer=LI1_cond $X=0.265 $Y=0.825
+ $X2=0.265 $Y2=1.915
r136 20 46 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=0.655
+ $X2=0.265 $Y2=0.74
r137 20 22 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.265 $Y=0.655
+ $X2=0.265 $Y2=0.445
r138 18 60 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.105 $Y=1.985
+ $X2=3.105 $Y2=1.325
r139 15 59 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.105 $Y=0.56
+ $X2=3.105 $Y2=0.995
r140 4 36 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.705 $X2=1.82 $Y2=1.915
r141 3 26 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.705 $X2=0.26 $Y2=1.915
r142 2 32 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.235 $X2=1.82 $Y2=0.445
r143 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%VPWR 1 2 9 13 18 19 20 22 32 33 36 39
c44 2 0 1.33802e-19 $X=2.465 $Y=1.705
r45 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r48 30 37 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.205 $Y=2.72
+ $X2=1.08 $Y2=2.72
r51 27 29 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.205 $Y=2.72
+ $X2=2.53 $Y2=2.72
r52 25 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 22 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=1.08 $Y2=2.72
r55 22 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 20 25 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 20 39 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 18 29 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=2.72
+ $X2=2.72 $Y2=2.72
r60 17 32 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.72
+ $X2=2.72 $Y2=2.72
r62 13 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.72 $Y=1.93
+ $X2=2.72 $Y2=2.34
r63 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=2.635
+ $X2=2.72 $Y2=2.72
r64 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.72 $Y=2.635
+ $X2=2.72 $Y2=2.34
r65 7 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2.635
+ $X2=1.08 $Y2=2.72
r66 7 9 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=1.08 $Y=2.635 $X2=1.08
+ $Y2=1.915
r67 2 16 600 $w=1.7e-07 $l=7.51765e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.705 $X2=2.72 $Y2=2.34
r68 2 13 600 $w=1.7e-07 $l=3.49857e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.705 $X2=2.72 $Y2=1.93
r69 1 9 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.705 $X2=1.04 $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%X 1 2 9 12 13 14 15 16 26 33 46
r29 46 47 2.39662 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.43 $Y=1.53
+ $X2=3.43 $Y2=1.495
r30 33 44 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=3.482 $Y=0.85
+ $X2=3.482 $Y2=0.825
r31 16 40 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.43 $Y=1.87
+ $X2=3.43 $Y2=1.66
r32 15 40 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.43 $Y=1.555
+ $X2=3.43 $Y2=1.66
r33 15 46 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.43 $Y=1.555
+ $X2=3.43 $Y2=1.53
r34 15 47 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=3.482 $Y=1.47
+ $X2=3.482 $Y2=1.495
r35 14 15 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=3.482 $Y=1.19
+ $X2=3.482 $Y2=1.47
r36 13 44 2.33681 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=3.425 $Y=0.795
+ $X2=3.425 $Y2=0.825
r37 13 24 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=3.425 $Y=0.795
+ $X2=3.425 $Y2=0.655
r38 13 14 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=3.482 $Y=0.88
+ $X2=3.482 $Y2=1.19
r39 13 33 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=3.482 $Y=0.88
+ $X2=3.482 $Y2=0.85
r40 12 24 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=3.425 $Y=0.51
+ $X2=3.425 $Y2=0.655
r41 12 26 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=3.425 $Y=0.51
+ $X2=3.425 $Y2=0.38
r42 10 16 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.43 $Y=2.16
+ $X2=3.43 $Y2=1.87
r43 9 10 6.10117 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=3.425 $Y=2.34
+ $X2=3.425 $Y2=2.16
r44 2 40 300 $w=1.7e-07 $l=3.15595e-07 $layer=licon1_PDIFF $count=2 $X=3.18
+ $Y=1.485 $X2=3.42 $Y2=1.66
r45 2 9 600 $w=1.7e-07 $l=9.67587e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.42 $Y2=2.34
r46 1 26 91 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=2 $X=3.18
+ $Y=0.235 $X2=3.42 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MAJ3_1%VGND 1 2 9 13 16 17 18 20 30 31 34 37
r53 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r56 28 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.15
+ $Y2=0
r57 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r58 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.04
+ $Y2=0
r59 25 27 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=2.53 $Y2=0
r60 23 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r61 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r62 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.04
+ $Y2=0
r63 20 22 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.69
+ $Y2=0
r64 18 23 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r65 18 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r66 16 27 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r67 16 17 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.712
+ $Y2=0
r68 15 30 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=3.45
+ $Y2=0
r69 15 17 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.88 $Y=0 $X2=2.712
+ $Y2=0
r70 11 17 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.712 $Y=0.085
+ $X2=2.712 $Y2=0
r71 11 13 10.3204 $w=3.33e-07 $l=3e-07 $layer=LI1_cond $X=2.712 $Y=0.085
+ $X2=2.712 $Y2=0.385
r72 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.04 $Y=0.085 $X2=1.04
+ $Y2=0
r73 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.04 $Y=0.085
+ $X2=1.04 $Y2=0.4
r74 2 13 182 $w=1.7e-07 $l=3.11087e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.71 $Y2=0.385
r75 1 9 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.905
+ $Y=0.235 $X2=1.04 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__or2b_4.spice.pex
* Created: Thu Aug 27 14:43:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR2B_4%B_N 3 7 9 10 11 19
c24 9 0 1.76169e-19 $X=0.23 $Y=1.19
r25 16 19 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r26 10 11 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.53
+ $X2=0.257 $Y2=1.87
r27 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.16
+ $X2=0.257 $Y2=1.53
r28 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r29 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r31 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%A_27_53# 1 2 7 9 12 14 15 18 20 21 22 24
c58 14 0 1.76169e-19 $X=1.295 $Y=1.16
r59 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=1.16 $X2=1.005 $Y2=1.16
r60 22 28 9.1679 $w=4.03e-07 $l=2.46037e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.857 $Y2=1.16
r61 22 24 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.68 $Y=1.325
+ $X2=0.68 $Y2=2.2
r62 20 28 10.2928 $w=4.03e-07 $l=4.52416e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.857 $Y2=1.16
r63 20 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.42 $Y2=0.82
r64 16 21 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.42 $Y2=0.82
r65 16 18 10.7809 $w=3.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=0.735
+ $X2=0.265 $Y2=0.445
r66 14 29 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.295 $Y=1.16
+ $X2=1.005 $Y2=1.16
r67 14 15 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.295 $Y=1.16
+ $X2=1.4 $Y2=1.16
r68 10 15 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.4 $Y2=1.16
r69 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.985
r70 7 15 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=1.37 $Y=0.995
+ $X2=1.4 $Y2=1.16
r71 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.37 $Y=0.995 $X2=1.37
+ $Y2=0.56
r72 2 24 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.2
r73 1 18 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%A 3 6 8 11 13
c33 11 0 8.29716e-20 $X=1.85 $Y=1.16
r34 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=1.325
r35 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.16
+ $X2=1.85 $Y2=0.995
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r37 8 12 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=2.07 $Y=1.175 $X2=1.85
+ $Y2=1.175
r38 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.79 $Y=1.985
+ $X2=1.79 $Y2=1.325
r39 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.79 $Y=0.56 $X2=1.79
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%A_219_297# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 42 45 47 49 50 53 56 58 68
c123 49 0 8.29716e-20 $X=2.575 $Y=1.245
r124 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.7 $Y=1.16
+ $X2=3.12 $Y2=1.16
r125 61 65 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.655 $Y=1.16
+ $X2=2.7 $Y2=1.16
r126 61 62 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.655 $Y=1.16
+ $X2=2.28 $Y2=1.16
r127 60 61 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.16 $X2=2.655 $Y2=1.16
r128 57 58 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.517 $Y=0.735
+ $X2=1.517 $Y2=0.905
r129 54 68 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.335 $Y=1.16
+ $X2=3.54 $Y2=1.16
r130 54 66 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.335 $Y=1.16
+ $X2=3.12 $Y2=1.16
r131 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.335
+ $Y=1.16 $X2=3.335 $Y2=1.16
r132 51 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.16
+ $X2=2.575 $Y2=1.16
r133 51 53 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.66 $Y=1.16
+ $X2=3.335 $Y2=1.16
r134 49 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=1.245
+ $X2=2.575 $Y2=1.16
r135 49 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.575 $Y=1.245
+ $X2=2.575 $Y2=1.445
r136 48 56 3.69268 $w=1.7e-07 $l=4.87186e-07 $layer=LI1_cond $X=1.46 $Y=1.53
+ $X2=0.99 $Y2=1.495
r137 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.49 $Y=1.53
+ $X2=2.575 $Y2=1.445
r138 47 48 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.49 $Y=1.53
+ $X2=1.46 $Y2=1.53
r139 45 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.58 $Y=0.4
+ $X2=1.58 $Y2=0.735
r140 42 56 2.96976 $w=3.2e-07 $l=4.09237e-07 $layer=LI1_cond $X=1.375 $Y=1.445
+ $X2=0.99 $Y2=1.495
r141 42 58 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.375 $Y=1.445
+ $X2=1.375 $Y2=0.905
r142 37 39 17.305 $w=4.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.225 $Y=1.63
+ $X2=1.225 $Y2=2.31
r143 35 56 2.96976 $w=3.2e-07 $l=2.88834e-07 $layer=LI1_cond $X=1.225 $Y=1.615
+ $X2=0.99 $Y2=1.495
r144 35 37 0.381727 $w=4.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.225 $Y=1.615
+ $X2=1.225 $Y2=1.63
r145 31 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.325
+ $X2=3.54 $Y2=1.16
r146 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.54 $Y=1.325
+ $X2=3.54 $Y2=1.985
r147 28 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=0.995
+ $X2=3.54 $Y2=1.16
r148 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.54 $Y=0.995
+ $X2=3.54 $Y2=0.56
r149 24 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.16
r150 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=1.325
+ $X2=3.12 $Y2=1.985
r151 21 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=1.16
r152 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.12 $Y=0.995
+ $X2=3.12 $Y2=0.56
r153 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.16
r154 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.325
+ $X2=2.7 $Y2=1.985
r155 14 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=1.16
r156 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=0.995
+ $X2=2.7 $Y2=0.56
r157 10 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.16
r158 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.28 $Y=1.325
+ $X2=2.28 $Y2=1.985
r159 7 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=1.16
r160 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.28 $Y=0.995
+ $X2=2.28 $Y2=0.56
r161 2 39 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.485 $X2=1.22 $Y2=2.31
r162 2 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.485 $X2=1.22 $Y2=1.63
r163 1 45 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 34 46
+ 54 58
r56 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r57 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 49 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r59 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 46 57 3.87298 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=3.625 $Y=2.72
+ $X2=3.882 $Y2=2.72
r61 46 48 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.625 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 45 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 42 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.055 $Y2=2.72
r66 42 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 41 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 37 40 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r72 35 51 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r73 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r74 34 54 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=2.055 $Y2=2.72
r75 34 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.915 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 32 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 30 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.53 $Y2=2.72
r79 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.785 $Y=2.72
+ $X2=2.91 $Y2=2.72
r80 29 48 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.035 $Y=2.72
+ $X2=2.91 $Y2=2.72
r82 25 57 3.27018 $w=2.5e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.882 $Y2=2.72
r83 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.75 $Y=2.635
+ $X2=3.75 $Y2=1.96
r84 21 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=2.635
+ $X2=2.91 $Y2=2.72
r85 21 23 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.91 $Y=2.635
+ $X2=2.91 $Y2=2.3
r86 17 54 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2.72
r87 17 19 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.055 $Y=2.635
+ $X2=2.055 $Y2=2
r88 13 51 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r89 13 15 15.5919 $w=2.53e-07 $l=3.45e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.29
r90 4 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.485 $X2=3.75 $Y2=1.96
r91 3 23 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.485 $X2=2.91 $Y2=2.3
r92 2 19 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=1.485 $X2=2.065 $Y2=2
r93 1 15 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%X 1 2 3 4 15 19 22 23 24 27 31 33 35 39 40 41
+ 43
r73 42 43 12.4275 $w=5.53e-07 $l=5.4e-07 $layer=LI1_cond $X=3.862 $Y=0.905
+ $X2=3.862 $Y2=1.445
r74 38 40 8.64074 $w=5.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.33 $Y=1.7
+ $X2=3.455 $Y2=1.7
r75 38 39 17.4354 $w=5.08e-07 $l=5e-07 $layer=LI1_cond $X=3.33 $Y=1.7 $X2=2.83
+ $Y2=1.7
r76 36 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.82
+ $X2=3.33 $Y2=0.82
r77 35 42 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=3.67 $Y=0.82
+ $X2=3.862 $Y2=0.905
r78 35 36 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=0.82
+ $X2=3.495 $Y2=0.82
r79 33 43 5.71163 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.67 $Y=1.53
+ $X2=3.862 $Y2=1.53
r80 33 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.67 $Y=1.53
+ $X2=3.455 $Y2=1.53
r81 29 38 4.91917 $w=2.5e-07 $l=2.55e-07 $layer=LI1_cond $X=3.33 $Y=1.955
+ $X2=3.33 $Y2=1.7
r82 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.33 $Y=1.955
+ $X2=3.33 $Y2=1.96
r83 25 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.735
+ $X2=3.33 $Y2=0.82
r84 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.33 $Y=0.735
+ $X2=3.33 $Y2=0.4
r85 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=0.82
+ $X2=3.33 $Y2=0.82
r86 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.165 $Y=0.82
+ $X2=2.655 $Y2=0.82
r87 22 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.615 $Y=1.87
+ $X2=2.83 $Y2=1.87
r88 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.49 $Y=1.955
+ $X2=2.615 $Y2=1.87
r89 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.49 $Y=1.955
+ $X2=2.49 $Y2=1.96
r90 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=0.735
+ $X2=2.655 $Y2=0.82
r91 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.49 $Y=0.735
+ $X2=2.49 $Y2=0.4
r92 4 38 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.485 $X2=3.33 $Y2=1.62
r93 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=1.485 $X2=3.33 $Y2=1.96
r94 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.49 $Y2=1.96
r95 2 27 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=3.195
+ $Y=0.235 $X2=3.33 $Y2=0.4
r96 1 15 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.235 $X2=2.49 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_4%VGND 1 2 3 4 15 19 23 26 27 29 30 31 38 51 52
+ 56 65 67
r65 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r66 64 65 9.00983 $w=6.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.24
+ $X2=1.245 $Y2=0.24
r67 61 64 0.184012 $w=6.48e-07 $l=1e-08 $layer=LI1_cond $X=1.15 $Y=0.24 $X2=1.16
+ $Y2=0.24
r68 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 59 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r70 58 61 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r71 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r72 55 58 0.184012 $w=6.48e-07 $l=1e-08 $layer=LI1_cond $X=0.68 $Y=0.24 $X2=0.69
+ $Y2=0.24
r73 55 56 9.10184 $w=6.48e-07 $l=9e-08 $layer=LI1_cond $X=0.68 $Y=0.24 $X2=0.59
+ $Y2=0.24
r74 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r75 49 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r76 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r77 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r78 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r79 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r80 43 67 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.067
+ $Y2=0
r81 43 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.53
+ $Y2=0
r82 42 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r83 42 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r84 41 65 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.245
+ $Y2=0
r85 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r86 38 67 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=1.98 $Y=0 $X2=2.067
+ $Y2=0
r87 38 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=1.61
+ $Y2=0
r88 35 56 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.59
+ $Y2=0
r89 31 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r90 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 29 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.45
+ $Y2=0
r92 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.75
+ $Y2=0
r93 28 51 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.91
+ $Y2=0
r94 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.75
+ $Y2=0
r95 26 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.53
+ $Y2=0
r96 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.91
+ $Y2=0
r97 25 48 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.995 $Y=0 $X2=3.45
+ $Y2=0
r98 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.91
+ $Y2=0
r99 21 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0
r100 21 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0.385
r101 17 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0
r102 17 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0.385
r103 13 67 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.067 $Y=0.085
+ $X2=2.067 $Y2=0
r104 13 15 19.9636 $w=1.73e-07 $l=3.15e-07 $layer=LI1_cond $X=2.067 $Y=0.085
+ $X2=2.067 $Y2=0.4
r105 4 23 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.235 $X2=3.75 $Y2=0.385
r106 3 19 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.235 $X2=2.91 $Y2=0.385
r107 2 15 91 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.235 $X2=2.07 $Y2=0.4
r108 1 64 182 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=1.16 $Y2=0.4
r109 1 55 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.68 $Y2=0.4
.ends


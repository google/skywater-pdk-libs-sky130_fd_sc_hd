* File: sky130_fd_sc_hd__o32a_1.spice
* Created: Thu Aug 27 14:40:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o32a_1.spice.pex"
.subckt sky130_fd_sc_hd__o32a_1  VNB VPB A1 A2 A3 B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_77_199#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_227_47#_M1005_d N_A1_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=5.532 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_227_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.10725 PD=1.04 PS=0.98 NRD=10.152 NRS=3.684 M=1 R=4.33333
+ SA=75001.1 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_A_227_47#_M1001_d N_A3_M1001_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.12675 PD=1.04 PS=1.04 NRD=14.76 NRS=10.152 M=1 R=4.33333
+ SA=75001.6 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1011 N_A_77_199#_M1011_d N_B2_M1011_g N_A_227_47#_M1001_d VNB NSHORT L=0.15
+ W=0.65 AD=0.13325 AS=0.12675 PD=1.06 PS=1.04 NRD=7.38 NRS=5.532 M=1 R=4.33333
+ SA=75002.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1006 N_A_227_47#_M1006_d N_B1_M1006_g N_A_77_199#_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.1885 AS=0.13325 PD=1.88 PS=1.06 NRD=0 NRS=16.608 M=1 R=4.33333
+ SA=75002.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_77_199#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.335 PD=1.27 PS=2.67 NRD=0 NRS=7.8603 M=1 R=6.66667 SA=75000.3
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1010 A_227_297# N_A1_M1010_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=0 M=1 R=6.66667 SA=75000.7 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1003 A_323_297# N_A2_M1003_g A_227_297# VPB PHIGHVT L=0.15 W=1 AD=0.195
+ AS=0.165 PD=1.39 PS=1.33 NRD=27.5603 NRS=21.6503 M=1 R=6.66667 SA=75001.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1000 N_A_77_199#_M1000_d N_A3_M1000_g A_323_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=9.8303 NRS=27.5603 M=1 R=6.66667
+ SA=75001.7 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1007 A_539_297# N_B2_M1007_g N_A_77_199#_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.205 AS=0.195 PD=1.41 PS=1.39 NRD=29.5303 NRS=11.8003 M=1 R=6.66667
+ SA=75002.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g A_539_297# VPB PHIGHVT L=0.15 W=1 AD=0.29
+ AS=0.205 PD=2.58 PS=1.41 NRD=0 NRS=29.5303 M=1 R=6.66667 SA=75002.8 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_61 VPB 0 1.23066e-19 $X=0.14 $Y=2.635
*
.include "sky130_fd_sc_hd__o32a_1.spice.SKY130_FD_SC_HD__O32A_1.pxi"
*
.ends
*
*

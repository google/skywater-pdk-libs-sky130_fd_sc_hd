* File: sky130_fd_sc_hd__a21bo_1.spice.SKY130_FD_SC_HD__A21BO_1.pxi
* Created: Thu Aug 27 14:00:02 2020
* 
x_PM_SKY130_FD_SC_HD__A21BO_1%B1_N N_B1_N_c_66_n N_B1_N_c_67_n N_B1_N_c_71_n
+ N_B1_N_M1002_g N_B1_N_c_68_n N_B1_N_M1005_g N_B1_N_c_72_n B1_N B1_N B1_N B1_N
+ N_B1_N_c_70_n PM_SKY130_FD_SC_HD__A21BO_1%B1_N
x_PM_SKY130_FD_SC_HD__A21BO_1%A_27_413# N_A_27_413#_M1005_s N_A_27_413#_M1002_s
+ N_A_27_413#_c_104_n N_A_27_413#_M1009_g N_A_27_413#_c_111_n
+ N_A_27_413#_M1000_g N_A_27_413#_c_106_n N_A_27_413#_c_113_n
+ N_A_27_413#_c_107_n N_A_27_413#_c_108_n N_A_27_413#_c_114_n
+ N_A_27_413#_c_115_n N_A_27_413#_c_109_n PM_SKY130_FD_SC_HD__A21BO_1%A_27_413#
x_PM_SKY130_FD_SC_HD__A21BO_1%A1 N_A1_M1008_g N_A1_M1006_g A1 A1 N_A1_c_169_n
+ N_A1_c_170_n N_A1_c_171_n PM_SKY130_FD_SC_HD__A21BO_1%A1
x_PM_SKY130_FD_SC_HD__A21BO_1%A2 N_A2_c_206_n N_A2_M1004_g N_A2_M1003_g A2 A2
+ N_A2_c_208_n PM_SKY130_FD_SC_HD__A21BO_1%A2
x_PM_SKY130_FD_SC_HD__A21BO_1%A_215_297# N_A_215_297#_M1009_d
+ N_A_215_297#_M1000_s N_A_215_297#_c_241_n N_A_215_297#_M1007_g
+ N_A_215_297#_M1001_g N_A_215_297#_c_247_n N_A_215_297#_c_242_n
+ N_A_215_297#_c_273_n N_A_215_297#_c_243_n N_A_215_297#_c_244_n
+ N_A_215_297#_c_253_n N_A_215_297#_c_245_n
+ PM_SKY130_FD_SC_HD__A21BO_1%A_215_297#
x_PM_SKY130_FD_SC_HD__A21BO_1%VPWR N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_M1001_s
+ N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n VPWR N_VPWR_c_321_n
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_317_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n PM_SKY130_FD_SC_HD__A21BO_1%VPWR
x_PM_SKY130_FD_SC_HD__A21BO_1%A_298_297# N_A_298_297#_M1000_d
+ N_A_298_297#_M1003_d N_A_298_297#_c_376_n N_A_298_297#_c_382_n
+ N_A_298_297#_c_380_n PM_SKY130_FD_SC_HD__A21BO_1%A_298_297#
x_PM_SKY130_FD_SC_HD__A21BO_1%X N_X_M1007_d N_X_M1001_d X X X X X X
+ PM_SKY130_FD_SC_HD__A21BO_1%X
x_PM_SKY130_FD_SC_HD__A21BO_1%VGND N_VGND_M1005_d N_VGND_M1004_d N_VGND_c_406_n
+ VGND N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n PM_SKY130_FD_SC_HD__A21BO_1%VGND
cc_1 VNB N_B1_N_c_66_n 0.0362948f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.83
cc_2 VNB N_B1_N_c_67_n 0.0206114f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=0.83
cc_3 VNB N_B1_N_c_68_n 0.0208821f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=0.755
cc_4 VNB B1_N 0.0223168f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_5 VNB N_B1_N_c_70_n 0.0398605f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_6 VNB N_A_27_413#_c_104_n 0.0208294f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=0.445
cc_7 VNB N_A_27_413#_M1009_g 0.0283255f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_8 VNB N_A_27_413#_c_106_n 0.00318682f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_9 VNB N_A_27_413#_c_107_n 0.00531009f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_10 VNB N_A_27_413#_c_108_n 0.00233044f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_11 VNB N_A_27_413#_c_109_n 0.00824026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_169_n 0.0205063f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.89
cc_13 VNB N_A1_c_170_n 0.00466283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_171_n 0.0165619f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_15 VNB N_A2_c_206_n 0.0202629f $X=-0.19 $Y=-0.24 $X2=0.74 $Y2=0.83
cc_16 VNB A2 0.00454214f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=0.445
cc_17 VNB N_A2_c_208_n 0.0304111f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_18 VNB N_A_215_297#_c_241_n 0.022309f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=0.445
cc_19 VNB N_A_215_297#_c_242_n 0.00164823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_297#_c_243_n 0.00421745f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=0.51
cc_21 VNB N_A_215_297#_c_244_n 0.0101121f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.16
cc_22 VNB N_A_215_297#_c_245_n 0.0331829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_317_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB X 0.0458952f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=0.445
cc_25 VNB N_VGND_c_406_n 0.00709f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=0.905
cc_26 VNB N_VGND_c_407_n 0.0282268f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_27 VNB N_VGND_c_408_n 0.0180353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_409_n 0.204974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_410_n 0.00471252f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=1.16
cc_30 VNB N_VGND_c_411_n 0.0309008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_412_n 0.0219033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_B1_N_c_71_n 0.0221206f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.965
cc_33 VPB N_B1_N_c_72_n 0.0329977f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.89
cc_34 VPB N_B1_N_c_70_n 0.0498291f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_35 VPB N_A_27_413#_c_104_n 0.0146384f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.445
cc_36 VPB N_A_27_413#_c_111_n 0.0186745f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.89
cc_37 VPB N_A_27_413#_c_106_n 0.0025294f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_38 VPB N_A_27_413#_c_113_n 0.0151368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_413#_c_114_n 0.0151053f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=0.51
cc_40 VPB N_A_27_413#_c_115_n 0.00647464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_413#_c_109_n 0.0246292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A1_M1006_g 0.0171313f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.755
cc_43 VPB N_A1_c_169_n 0.0045919f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.89
cc_44 VPB N_A1_c_170_n 0.00249245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A2_M1003_g 0.0220104f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.755
cc_46 VPB A2 0.0051489f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.445
cc_47 VPB N_A2_c_208_n 0.00922834f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_48 VPB N_A_215_297#_M1001_g 0.0263573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_215_297#_c_247_n 0.0104272f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_50 VPB N_A_215_297#_c_243_n 0.00255235f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=0.51
cc_51 VPB N_A_215_297#_c_244_n 0.002514f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_52 VPB N_A_215_297#_c_245_n 0.00971524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_318_n 0.00629611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_319_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_55 VPB N_VPWR_c_320_n 0.0165295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_321_n 0.014663f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=0.51
cc_57 VPB N_VPWR_c_322_n 0.0260519f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_58 VPB N_VPWR_c_323_n 0.016105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_324_n 0.0177171f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_317_n 0.0612292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_326_n 0.00545784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_327_n 0.00436716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_328_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB X 0.0469694f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.445
cc_65 N_B1_N_c_68_n N_A_27_413#_M1009_g 0.015982f $X=0.815 $Y=0.755 $X2=0 $Y2=0
cc_66 N_B1_N_c_71_n N_A_27_413#_c_113_n 9.84418e-19 $X=0.47 $Y=1.965 $X2=0 $Y2=0
cc_67 N_B1_N_c_72_n N_A_27_413#_c_113_n 0.00171886f $X=0.47 $Y=1.89 $X2=0 $Y2=0
cc_68 N_B1_N_c_66_n N_A_27_413#_c_107_n 0.0155659f $X=0.74 $Y=0.83 $X2=0 $Y2=0
cc_69 N_B1_N_c_68_n N_A_27_413#_c_107_n 0.00680553f $X=0.815 $Y=0.755 $X2=0
+ $Y2=0
cc_70 B1_N N_A_27_413#_c_107_n 0.097832f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_71 N_B1_N_c_70_n N_A_27_413#_c_107_n 0.0163227f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B1_N_c_66_n N_A_27_413#_c_108_n 0.00280248f $X=0.74 $Y=0.83 $X2=0 $Y2=0
cc_73 N_B1_N_c_71_n N_A_27_413#_c_114_n 0.00753037f $X=0.47 $Y=1.965 $X2=0 $Y2=0
cc_74 N_B1_N_c_72_n N_A_27_413#_c_114_n 0.024097f $X=0.47 $Y=1.89 $X2=0 $Y2=0
cc_75 B1_N N_A_27_413#_c_114_n 0.016773f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_76 N_B1_N_c_72_n N_A_27_413#_c_115_n 0.00284219f $X=0.47 $Y=1.89 $X2=0 $Y2=0
cc_77 N_B1_N_c_66_n N_A_27_413#_c_109_n 0.014593f $X=0.74 $Y=0.83 $X2=0 $Y2=0
cc_78 B1_N N_A_27_413#_c_109_n 4.32293e-19 $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_79 N_B1_N_c_70_n N_A_27_413#_c_109_n 0.0258101f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B1_N_c_71_n N_A_215_297#_c_247_n 0.00383273f $X=0.47 $Y=1.965 $X2=0
+ $Y2=0
cc_81 N_B1_N_c_72_n N_A_215_297#_c_247_n 8.66108e-19 $X=0.47 $Y=1.89 $X2=0 $Y2=0
cc_82 N_B1_N_c_66_n N_A_215_297#_c_253_n 3.41491e-19 $X=0.74 $Y=0.83 $X2=0 $Y2=0
cc_83 N_B1_N_c_71_n N_VPWR_c_318_n 0.0108265f $X=0.47 $Y=1.965 $X2=0 $Y2=0
cc_84 N_B1_N_c_71_n N_VPWR_c_321_n 0.00343969f $X=0.47 $Y=1.965 $X2=0 $Y2=0
cc_85 N_B1_N_c_72_n N_VPWR_c_321_n 3.04006e-19 $X=0.47 $Y=1.89 $X2=0 $Y2=0
cc_86 N_B1_N_c_71_n N_VPWR_c_317_n 0.00505663f $X=0.47 $Y=1.965 $X2=0 $Y2=0
cc_87 N_B1_N_c_68_n N_VGND_c_406_n 0.00800034f $X=0.815 $Y=0.755 $X2=0 $Y2=0
cc_88 N_B1_N_c_66_n N_VGND_c_407_n 5.08484e-19 $X=0.74 $Y=0.83 $X2=0 $Y2=0
cc_89 N_B1_N_c_67_n N_VGND_c_407_n 0.00357448f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_90 N_B1_N_c_68_n N_VGND_c_407_n 0.00579368f $X=0.815 $Y=0.755 $X2=0 $Y2=0
cc_91 B1_N N_VGND_c_407_n 0.0113151f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_92 N_B1_N_c_67_n N_VGND_c_409_n 0.00411268f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_93 N_B1_N_c_68_n N_VGND_c_409_n 0.0123166f $X=0.815 $Y=0.755 $X2=0 $Y2=0
cc_94 B1_N N_VGND_c_409_n 0.00846606f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_95 N_A_27_413#_c_106_n N_A1_M1006_g 0.026262f $X=1.415 $Y=1.285 $X2=0 $Y2=0
cc_96 N_A_27_413#_M1009_g N_A1_c_169_n 0.0190178f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_97 N_A_27_413#_M1009_g N_A1_c_170_n 3.23241e-19 $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_98 N_A_27_413#_c_106_n N_A1_c_170_n 0.00151655f $X=1.415 $Y=1.285 $X2=0 $Y2=0
cc_99 N_A_27_413#_M1009_g N_A1_c_171_n 0.011482f $X=1.415 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A_27_413#_c_104_n N_A_215_297#_c_247_n 0.00785716f $X=1.34 $Y=1.285
+ $X2=0 $Y2=0
cc_101 N_A_27_413#_c_111_n N_A_215_297#_c_247_n 0.0148281f $X=1.415 $Y=1.385
+ $X2=0 $Y2=0
cc_102 N_A_27_413#_c_106_n N_A_215_297#_c_247_n 6.70457e-19 $X=1.415 $Y=1.285
+ $X2=0 $Y2=0
cc_103 N_A_27_413#_c_114_n N_A_215_297#_c_247_n 0.0168192f $X=0.685 $Y=1.845
+ $X2=0 $Y2=0
cc_104 N_A_27_413#_c_115_n N_A_215_297#_c_247_n 0.0388279f $X=0.72 $Y=1.44 $X2=0
+ $Y2=0
cc_105 N_A_27_413#_c_109_n N_A_215_297#_c_247_n 0.00190392f $X=0.72 $Y=1.285
+ $X2=0 $Y2=0
cc_106 N_A_27_413#_M1009_g N_A_215_297#_c_242_n 0.00710966f $X=1.415 $Y=0.56
+ $X2=0 $Y2=0
cc_107 N_A_27_413#_c_107_n N_A_215_297#_c_242_n 0.00492807f $X=0.6 $Y=0.45 $X2=0
+ $Y2=0
cc_108 N_A_27_413#_c_104_n N_A_215_297#_c_244_n 0.0130017f $X=1.34 $Y=1.285
+ $X2=0 $Y2=0
cc_109 N_A_27_413#_M1009_g N_A_215_297#_c_244_n 0.00673267f $X=1.415 $Y=0.56
+ $X2=0 $Y2=0
cc_110 N_A_27_413#_c_106_n N_A_215_297#_c_244_n 0.00898417f $X=1.415 $Y=1.285
+ $X2=0 $Y2=0
cc_111 N_A_27_413#_c_107_n N_A_215_297#_c_244_n 0.00691896f $X=0.6 $Y=0.45 $X2=0
+ $Y2=0
cc_112 N_A_27_413#_c_108_n N_A_215_297#_c_244_n 0.0135717f $X=0.685 $Y=1.335
+ $X2=0 $Y2=0
cc_113 N_A_27_413#_M1009_g N_A_215_297#_c_253_n 0.0106194f $X=1.415 $Y=0.56
+ $X2=0 $Y2=0
cc_114 N_A_27_413#_c_111_n N_VPWR_c_318_n 0.00257049f $X=1.415 $Y=1.385 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_114_n N_VPWR_c_318_n 0.0230597f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_116 N_A_27_413#_c_111_n N_VPWR_c_319_n 0.00120409f $X=1.415 $Y=1.385 $X2=0
+ $Y2=0
cc_117 N_A_27_413#_c_113_n N_VPWR_c_321_n 0.0133604f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_118 N_A_27_413#_c_114_n N_VPWR_c_321_n 0.00268735f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_119 N_A_27_413#_c_111_n N_VPWR_c_322_n 0.00549284f $X=1.415 $Y=1.385 $X2=0
+ $Y2=0
cc_120 N_A_27_413#_M1002_s N_VPWR_c_317_n 0.00232867f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_121 N_A_27_413#_c_111_n N_VPWR_c_317_n 0.0111628f $X=1.415 $Y=1.385 $X2=0
+ $Y2=0
cc_122 N_A_27_413#_c_113_n N_VPWR_c_317_n 0.0088929f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_123 N_A_27_413#_c_114_n N_VPWR_c_317_n 0.005636f $X=0.685 $Y=1.845 $X2=0
+ $Y2=0
cc_124 N_A_27_413#_c_104_n N_VGND_c_406_n 0.00408228f $X=1.34 $Y=1.285 $X2=0
+ $Y2=0
cc_125 N_A_27_413#_M1009_g N_VGND_c_406_n 0.00780909f $X=1.415 $Y=0.56 $X2=0
+ $Y2=0
cc_126 N_A_27_413#_c_107_n N_VGND_c_406_n 0.0260855f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_127 N_A_27_413#_c_107_n N_VGND_c_407_n 0.0131702f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_128 N_A_27_413#_M1005_s N_VGND_c_409_n 0.00262373f $X=0.475 $Y=0.235 $X2=0
+ $Y2=0
cc_129 N_A_27_413#_M1009_g N_VGND_c_409_n 0.00645325f $X=1.415 $Y=0.56 $X2=0
+ $Y2=0
cc_130 N_A_27_413#_c_107_n N_VGND_c_409_n 0.00871059f $X=0.6 $Y=0.45 $X2=0 $Y2=0
cc_131 N_A_27_413#_M1009_g N_VGND_c_411_n 0.00391345f $X=1.415 $Y=0.56 $X2=0
+ $Y2=0
cc_132 N_A1_c_171_n N_A2_c_206_n 0.0405088f $X=1.845 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A1_M1006_g N_A2_M1003_g 0.0397966f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A1_c_169_n A2 2.29085e-19 $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A1_c_170_n A2 0.0356787f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_c_169_n N_A2_c_208_n 0.020677f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_c_170_n N_A2_c_208_n 0.00487013f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A1_M1006_g N_A_215_297#_c_247_n 0.00105527f $X=1.835 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A1_c_170_n N_A_215_297#_c_247_n 0.00863938f $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A1_c_169_n N_A_215_297#_c_242_n 2.92424e-19 $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A1_c_170_n N_A_215_297#_c_242_n 0.00390684f $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A1_c_171_n N_A_215_297#_c_242_n 0.00360403f $X=1.845 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A1_c_169_n N_A_215_297#_c_273_n 3.59559e-19 $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A1_c_170_n N_A_215_297#_c_273_n 0.0259761f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_c_171_n N_A_215_297#_c_273_n 0.00927988f $X=1.845 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_A1_c_169_n N_A_215_297#_c_244_n 0.00179433f $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A1_c_170_n N_A_215_297#_c_244_n 0.0251992f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A1_c_170_n N_A_215_297#_c_253_n 0.00260947f $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A1_c_171_n N_A_215_297#_c_253_n 0.00853354f $X=1.845 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A1_c_170_n N_VPWR_M1006_d 0.00207672f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A1_M1006_g N_VPWR_c_319_n 0.00926151f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A1_M1006_g N_VPWR_c_322_n 0.00365202f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A1_M1006_g N_VPWR_c_317_n 0.00431919f $X=1.835 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_M1006_g N_A_298_297#_c_376_n 0.0106382f $X=1.835 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A1_c_170_n N_A_298_297#_c_376_n 0.024986f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_c_171_n N_VGND_c_409_n 0.00576843f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A1_c_171_n N_VGND_c_411_n 0.00412344f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_158 A2 N_A_215_297#_M1001_g 0.00282072f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A2_c_206_n N_A_215_297#_c_273_n 0.0194864f $X=2.265 $Y=0.995 $X2=0
+ $Y2=0
cc_160 A2 N_A_215_297#_c_273_n 0.0185637f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A2_c_208_n N_A_215_297#_c_273_n 0.00161783f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A2_c_206_n N_A_215_297#_c_243_n 0.00456157f $X=2.265 $Y=0.995 $X2=0
+ $Y2=0
cc_163 A2 N_A_215_297#_c_243_n 0.0228466f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A2_c_208_n N_A_215_297#_c_243_n 0.00109545f $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A2_c_206_n N_A_215_297#_c_253_n 0.00150262f $X=2.265 $Y=0.995 $X2=0
+ $Y2=0
cc_166 A2 N_A_215_297#_c_245_n 0.00107098f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A2_c_208_n N_A_215_297#_c_245_n 0.0164764f $X=2.475 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VPWR_c_319_n 0.00856494f $X=2.265 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_VPWR_c_320_n 0.00671408f $X=2.265 $Y=1.985 $X2=0 $Y2=0
cc_170 A2 N_VPWR_c_320_n 0.00881347f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A2_M1003_g N_VPWR_c_323_n 0.00365202f $X=2.265 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A2_M1003_g N_VPWR_c_317_n 0.00561806f $X=2.265 $Y=1.985 $X2=0 $Y2=0
cc_173 A2 N_A_298_297#_M1003_d 0.005012f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_M1003_g N_A_298_297#_c_376_n 0.0153058f $X=2.265 $Y=1.985 $X2=0
+ $Y2=0
cc_175 A2 N_A_298_297#_c_380_n 0.0145803f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A2_c_208_n N_A_298_297#_c_380_n 6.99907e-19 $X=2.475 $Y=1.16 $X2=0
+ $Y2=0
cc_177 A2 X 0.00503432f $X=2.435 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A2_c_206_n N_VGND_c_409_n 0.00710803f $X=2.265 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A2_c_206_n N_VGND_c_411_n 0.0042361f $X=2.265 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_206_n N_VGND_c_412_n 0.00930856f $X=2.265 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_215_297#_c_247_n N_VPWR_c_318_n 0.0192373f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_182 N_A_215_297#_M1001_g N_VPWR_c_320_n 0.00473775f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_215_297#_c_243_n N_VPWR_c_320_n 0.0218437f $X=3.005 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_215_297#_c_245_n N_VPWR_c_320_n 0.00174884f $X=3.21 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_215_297#_c_247_n N_VPWR_c_322_n 0.0197891f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_186 N_A_215_297#_M1001_g N_VPWR_c_324_n 0.00585385f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_215_297#_M1000_s N_VPWR_c_317_n 0.00213747f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_188 N_A_215_297#_M1001_g N_VPWR_c_317_n 0.0128672f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_215_297#_c_247_n N_VPWR_c_317_n 0.0123896f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_190 N_A_215_297#_c_244_n N_A_298_297#_c_382_n 0.00168982f $X=1.47 $Y=1.195
+ $X2=0 $Y2=0
cc_191 N_A_215_297#_c_241_n X 0.0265335f $X=3.21 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_215_297#_c_243_n X 0.0302729f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_215_297#_c_273_n N_VGND_M1004_d 0.0230455f $X=2.84 $Y=0.72 $X2=0
+ $Y2=0
cc_194 N_A_215_297#_c_243_n N_VGND_M1004_d 0.00111895f $X=3.005 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_215_297#_c_244_n N_VGND_c_406_n 0.0127167f $X=1.47 $Y=1.195 $X2=0
+ $Y2=0
cc_196 N_A_215_297#_c_253_n N_VGND_c_406_n 0.0462329f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_197 N_A_215_297#_c_241_n N_VGND_c_408_n 0.00585385f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_215_297#_M1009_d N_VGND_c_409_n 0.00215535f $X=1.49 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_215_297#_c_241_n N_VGND_c_409_n 0.0130165f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_215_297#_c_273_n N_VGND_c_409_n 0.0187482f $X=2.84 $Y=0.72 $X2=0
+ $Y2=0
cc_201 N_A_215_297#_c_253_n N_VGND_c_409_n 0.0154886f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_202 N_A_215_297#_c_273_n N_VGND_c_411_n 0.00898324f $X=2.84 $Y=0.72 $X2=0
+ $Y2=0
cc_203 N_A_215_297#_c_253_n N_VGND_c_411_n 0.0240234f $X=1.625 $Y=0.38 $X2=0
+ $Y2=0
cc_204 N_A_215_297#_c_241_n N_VGND_c_412_n 0.00924068f $X=3.21 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_215_297#_c_273_n N_VGND_c_412_n 0.053646f $X=2.84 $Y=0.72 $X2=0 $Y2=0
cc_206 N_A_215_297#_c_245_n N_VGND_c_412_n 7.87819e-19 $X=3.21 $Y=1.16 $X2=0
+ $Y2=0
cc_207 N_A_215_297#_c_273_n A_382_47# 0.00465604f $X=2.84 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_208 N_VPWR_c_317_n N_A_298_297#_M1000_d 0.00393371f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_209 N_VPWR_c_317_n N_A_298_297#_M1003_d 0.00397607f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_M1006_d N_A_298_297#_c_376_n 0.00348901f $X=1.91 $Y=1.485 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_319_n N_A_298_297#_c_376_n 0.0166462f $X=2.05 $Y=2.24 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_322_n N_A_298_297#_c_376_n 0.00198277f $X=1.885 $Y=2.72 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_323_n N_A_298_297#_c_376_n 0.00202057f $X=2.825 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_317_n N_A_298_297#_c_376_n 0.00904154f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_322_n N_A_298_297#_c_382_n 0.0110342f $X=1.885 $Y=2.72 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_317_n N_A_298_297#_c_382_n 0.00681992f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_320_n N_A_298_297#_c_380_n 0.0387966f $X=3 $Y=1.66 $X2=0 $Y2=0
cc_218 N_VPWR_c_323_n N_A_298_297#_c_380_n 0.0108942f $X=2.825 $Y=2.72 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_317_n N_A_298_297#_c_380_n 0.00643678f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_317_n N_X_M1001_d 0.00265971f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_221 N_VPWR_c_324_n X 0.0170805f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_317_n X 0.0106557f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_223 X N_VGND_c_408_n 0.0170805f $X=3.365 $Y=0.425 $X2=0 $Y2=0
cc_224 N_X_M1007_d N_VGND_c_409_n 0.00265971f $X=3.285 $Y=0.235 $X2=0 $Y2=0
cc_225 X N_VGND_c_409_n 0.0106557f $X=3.365 $Y=0.425 $X2=0 $Y2=0
cc_226 N_VGND_c_409_n A_382_47# 0.00322965f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o211a_1.spice
* Created: Tue Sep  1 19:20:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211a_1.pex.spice"
.subckt sky130_fd_sc_hd__o211a_1  VNB VPB A1 A2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_79_21#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_215_47#_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.169 PD=0.975 PS=1.82 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1005 N_A_215_47#_M1005_d N_A2_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.105625 PD=1.09 PS=0.975 NRD=0 NRS=3.684 M=1 R=4.33333 SA=75000.7
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1006 A_510_47# N_B1_M1006_g N_A_215_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.143 PD=1 PS=1.09 NRD=22.152 NRS=30.456 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_A_79_21#_M1004_d N_C1_M1004_g A_510_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.195 AS=0.11375 PD=1.9 PS=1 NRD=6.456 NRS=22.152 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_79_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 A_297_297# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.1625
+ AS=0.26 PD=1.325 PS=2.52 NRD=21.1578 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.8
+ A=0.15 P=2.3 MULT=1
MM1008 N_A_79_21#_M1008_d N_A2_M1008_g A_297_297# VPB PHIGHVT L=0.15 W=1 AD=0.22
+ AS=0.1625 PD=1.44 PS=1.325 NRD=0 NRS=21.1578 M=1 R=6.66667 SA=75000.7
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_79_21#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.22 PD=1.35 PS=1.44 NRD=6.8753 NRS=32.4853 M=1 R=6.66667
+ SA=75001.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1003 N_A_79_21#_M1003_d N_C1_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3 AS=0.175 PD=2.6 PS=1.35 NRD=6.8753 NRS=6.8753 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__o211a_1.pxi.spice"
*
.ends
*
*

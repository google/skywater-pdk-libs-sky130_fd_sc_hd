* File: sky130_fd_sc_hd__xnor2_2.spice.pex
* Created: Thu Aug 27 14:49:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__XNOR2_2%B 1 3 6 8 10 13 15 17 20 22 24 27 29 35 37
+ 38 40 43 44 45 50 55
r119 44 45 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=2.93 $Y=1.53
+ $X2=1.15 $Y2=1.53
r120 43 45 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=1.53
+ $X2=1.15 $Y2=1.53
r121 41 55 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.755 $Y=1.16
+ $X2=4.02 $Y2=1.16
r122 41 52 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.755 $Y=1.16
+ $X2=3.565 $Y2=1.16
r123 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=1.16 $X2=3.755 $Y2=1.16
r124 38 40 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=3.1 $Y=1.18
+ $X2=3.755 $Y2=1.18
r125 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.445
+ $X2=2.93 $Y2=1.53
r126 36 38 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.015 $Y=1.285
+ $X2=3.1 $Y2=1.18
r127 36 37 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.015 $Y=1.285
+ $X2=3.015 $Y2=1.445
r128 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.875 $Y=1.445
+ $X2=0.96 $Y2=1.53
r129 34 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.875 $Y=1.285
+ $X2=0.875 $Y2=1.445
r130 32 50 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.65 $Y=1.16
+ $X2=0.905 $Y2=1.16
r131 32 47 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.16
+ $X2=0.485 $Y2=1.16
r132 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=1.16 $X2=0.65 $Y2=1.16
r133 29 34 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.79 $Y=1.18
+ $X2=0.875 $Y2=1.285
r134 29 31 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.79 $Y=1.18
+ $X2=0.65 $Y2=1.18
r135 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.325
+ $X2=4.02 $Y2=1.16
r136 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.02 $Y=1.325
+ $X2=4.02 $Y2=1.985
r137 22 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=0.995
+ $X2=4.02 $Y2=1.16
r138 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.02 $Y=0.995
+ $X2=4.02 $Y2=0.56
r139 18 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.16
r140 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=1.985
r141 15 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=1.16
r142 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.565 $Y=0.995
+ $X2=3.565 $Y2=0.56
r143 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.16
r144 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.325
+ $X2=0.905 $Y2=1.985
r145 8 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r146 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r147 4 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.16
r148 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.985
r149 1 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.16
r150 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 33
+ 35 38
c95 27 0 1.39696e-19 $X=3.145 $Y=1.985
c96 1 0 7.533e-20 $X=1.325 $Y=0.995
r97 42 44 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.42 $Y=1.16
+ $X2=1.745 $Y2=1.16
r98 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.42
+ $Y=1.16 $X2=1.42 $Y2=1.16
r99 39 42 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.325 $Y=1.16
+ $X2=1.42 $Y2=1.16
r100 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r101 35 44 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=1.745 $Y2=1.16
r102 35 37 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=2.46 $Y2=1.16
r103 33 38 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=2.46 $Y2=1.175
r104 33 43 36.0455 $w=1.98e-07 $l=6.5e-07 $layer=LI1_cond $X=2.07 $Y=1.175
+ $X2=1.42 $Y2=1.175
r105 30 31 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.725 $Y=1.16
+ $X2=3.145 $Y2=1.16
r106 29 37 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.65 $Y=1.16
+ $X2=2.46 $Y2=1.16
r107 29 30 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.16
+ $X2=2.725 $Y2=1.16
r108 25 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.16
r109 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=1.985
r110 22 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=1.16
r111 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=0.56
r112 18 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.325
+ $X2=2.725 $Y2=1.16
r113 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.725 $Y=1.325
+ $X2=2.725 $Y2=1.985
r114 15 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=0.995
+ $X2=2.725 $Y2=1.16
r115 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.725 $Y=0.995
+ $X2=2.725 $Y2=0.56
r116 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.16
r117 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.745 $Y=1.325
+ $X2=1.745 $Y2=1.985
r118 8 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=1.16
r119 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.745 $Y=0.995
+ $X2=1.745 $Y2=0.56
r120 4 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.16
r121 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.325 $Y=1.325
+ $X2=1.325 $Y2=1.985
r122 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=1.16
r123 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.325 $Y=0.995
+ $X2=1.325 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%A_27_297# 1 2 3 4 13 15 18 20 22 25 28 31 33
+ 35 39 43 46 47 48 50 51 53 57 59 61 65
c137 33 0 7.533e-20 $X=0.695 $Y=0.73
r138 54 65 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.13 $Y=1.16
+ $X2=5.38 $Y2=1.16
r139 54 62 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=5.13 $Y=1.16
+ $X2=4.96 $Y2=1.16
r140 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.16 $X2=5.13 $Y2=1.16
r141 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.805 $Y=1.16
+ $X2=5.13 $Y2=1.16
r142 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.72 $Y=1.245
+ $X2=4.805 $Y2=1.16
r143 49 50 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.72 $Y=1.245
+ $X2=4.72 $Y2=1.455
r144 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=1.54
+ $X2=4.72 $Y2=1.455
r145 47 48 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=4.635 $Y=1.54
+ $X2=3.48 $Y2=1.54
r146 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.395 $Y=1.625
+ $X2=3.48 $Y2=1.54
r147 45 46 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.395 $Y=1.625
+ $X2=3.395 $Y2=1.785
r148 44 61 6.87424 $w=1.75e-07 $l=1.27475e-07 $layer=LI1_cond $X=2.08 $Y=1.87
+ $X2=1.955 $Y2=1.875
r149 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.31 $Y=1.87
+ $X2=3.395 $Y2=1.785
r150 43 44 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.31 $Y=1.87
+ $X2=2.08 $Y2=1.87
r151 40 59 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.24 $Y=1.875
+ $X2=1.115 $Y2=1.875
r152 39 61 6.87424 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=1.875
+ $X2=1.955 $Y2=1.875
r153 39 40 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.83 $Y=1.875
+ $X2=1.24 $Y2=1.875
r154 36 57 2.8704 $w=1.8e-07 $l=1.58e-07 $layer=LI1_cond $X=0.4 $Y=1.875
+ $X2=0.242 $Y2=1.875
r155 35 59 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=0.99 $Y=1.875
+ $X2=1.115 $Y2=1.875
r156 35 36 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.99 $Y=1.875
+ $X2=0.4 $Y2=1.875
r157 31 33 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=0.315 $Y=0.77
+ $X2=0.695 $Y2=0.77
r158 28 57 3.61314 $w=2.72e-07 $l=1.08995e-07 $layer=LI1_cond $X=0.2 $Y=1.785
+ $X2=0.242 $Y2=1.875
r159 27 31 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.2 $Y=0.895
+ $X2=0.315 $Y2=0.77
r160 27 28 44.5945 $w=2.28e-07 $l=8.9e-07 $layer=LI1_cond $X=0.2 $Y=0.895
+ $X2=0.2 $Y2=1.785
r161 23 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.325
+ $X2=5.38 $Y2=1.16
r162 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.38 $Y=1.325
+ $X2=5.38 $Y2=1.985
r163 20 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=0.995
+ $X2=5.38 $Y2=1.16
r164 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.38 $Y=0.995
+ $X2=5.38 $Y2=0.56
r165 16 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=1.325
+ $X2=4.96 $Y2=1.16
r166 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.96 $Y=1.325
+ $X2=4.96 $Y2=1.985
r167 13 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=0.995
+ $X2=4.96 $Y2=1.16
r168 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.96 $Y=0.995
+ $X2=4.96 $Y2=0.56
r169 4 61 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.82
+ $Y=1.485 $X2=1.955 $Y2=1.96
r170 3 59 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.115 $Y2=1.96
r171 2 57 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
r172 1 33 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.695 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%VPWR 1 2 3 4 5 18 22 26 30 32 34 37 38 39 41
+ 46 51 60 65 68 71 75
c106 37 0 1.96631e-19 $X=4.625 $Y=2.72
r107 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r108 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 63 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r113 60 74 5.77705 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.722 $Y2=2.72
r114 60 62 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.29 $Y2=2.72
r115 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 59 72 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=2.99 $Y2=2.72
r117 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 56 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=2.935 $Y2=2.72
r119 56 58 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 55 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 55 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r123 52 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.66 $Y=2.72
+ $X2=1.535 $Y2=2.72
r124 52 54 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.66 $Y=2.72
+ $X2=2.53 $Y2=2.72
r125 51 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.935 $Y2=2.72
r126 51 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.53 $Y2=2.72
r127 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r128 50 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r129 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r130 47 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=0.695 $Y2=2.72
r131 47 49 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.82 $Y=2.72
+ $X2=1.15 $Y2=2.72
r132 46 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.535 $Y2=2.72
r133 46 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r134 41 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.695 $Y2=2.72
r135 41 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=2.72
+ $X2=0.23 $Y2=2.72
r136 39 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r138 37 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.37 $Y2=2.72
r139 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.75 $Y2=2.72
r140 36 62 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=5.29 $Y2=2.72
r141 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.75 $Y2=2.72
r142 32 74 2.85481 $w=4.3e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.68 $Y=2.635
+ $X2=5.722 $Y2=2.72
r143 32 34 18.0907 $w=4.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.68 $Y=2.635
+ $X2=5.68 $Y2=1.96
r144 28 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=2.635
+ $X2=4.75 $Y2=2.72
r145 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.75 $Y=2.635
+ $X2=4.75 $Y2=2.3
r146 24 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=2.635
+ $X2=2.935 $Y2=2.72
r147 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.935 $Y=2.635
+ $X2=2.935 $Y2=2.3
r148 20 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.635
+ $X2=1.535 $Y2=2.72
r149 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=2.635
+ $X2=1.535 $Y2=2.3
r150 16 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r151 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.3
r152 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.455
+ $Y=1.485 $X2=5.59 $Y2=1.96
r153 4 30 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.75 $Y2=2.3
r154 3 26 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.485 $X2=2.935 $Y2=2.3
r155 2 22 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=1.485 $X2=1.535 $Y2=2.3
r156 1 18 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.485 $X2=0.695 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%A_474_297# 1 2 3 10 13 17 18 21 24 25
c56 24 0 1.96631e-19 $X=3.47 $Y=2.21
c57 18 0 1.39696e-19 $X=2.695 $Y=2.21
r58 25 34 6.02816 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.392 $Y=2.21
+ $X2=3.392 $Y2=2.38
r59 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.47 $Y=2.21
+ $X2=3.47 $Y2=2.21
r60 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.55 $Y=2.21
+ $X2=2.55 $Y2=2.21
r61 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.21
+ $X2=2.55 $Y2=2.21
r62 17 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.325 $Y=2.21
+ $X2=3.47 $Y2=2.21
r63 17 18 0.779701 $w=1.4e-07 $l=6.3e-07 $layer=MET1_cond $X=3.325 $Y=2.21
+ $X2=2.695 $Y2=2.21
r64 13 15 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.23 $Y=2.3 $X2=4.23
+ $Y2=2.38
r65 11 34 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.555 $Y=2.38
+ $X2=3.392 $Y2=2.38
r66 10 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.105 $Y=2.38
+ $X2=4.23 $Y2=2.38
r67 10 11 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.105 $Y=2.38
+ $X2=3.555 $Y2=2.38
r68 3 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=1.485 $X2=4.23 $Y2=2.3
r69 2 25 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.485 $X2=3.355 $Y2=2.3
r70 1 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.485 $X2=2.515 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%Y 1 2 3 4 13 15 20 21 24 25 34
r52 25 28 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=3.83 $Y=1.88 $X2=3.83
+ $Y2=1.96
r53 22 34 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=5.7 $Y=1.52 $X2=5.79
+ $Y2=1.52
r54 22 37 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=5.7 $Y=1.52 $X2=5.17
+ $Y2=1.52
r55 22 24 20.2416 $w=3.88e-07 $l=6.85e-07 $layer=LI1_cond $X=5.7 $Y=1.415
+ $X2=5.7 $Y2=0.73
r56 21 33 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.7 $Y=0.475 $X2=5.7
+ $Y2=0.39
r57 21 24 7.5352 $w=3.88e-07 $l=2.55e-07 $layer=LI1_cond $X=5.7 $Y=0.475 $X2=5.7
+ $Y2=0.73
r58 20 31 3.18546 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=1.795
+ $X2=5.17 $Y2=1.96
r59 20 37 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.17 $Y=1.795
+ $X2=5.17 $Y2=1.625
r60 15 33 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.505 $Y=0.39
+ $X2=5.7 $Y2=0.39
r61 15 17 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.505 $Y=0.39
+ $X2=4.75 $Y2=0.39
r62 14 25 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.935 $Y=1.88
+ $X2=3.83 $Y2=1.88
r63 13 31 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=5.045 $Y=1.88
+ $X2=5.17 $Y2=1.96
r64 13 14 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.045 $Y=1.88
+ $X2=3.935 $Y2=1.88
r65 4 37 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=1.485 $X2=5.17 $Y2=1.62
r66 4 31 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=1.485 $X2=5.17 $Y2=1.96
r67 3 28 600 $w=1.7e-07 $l=5.53512e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=1.485 $X2=3.81 $Y2=1.96
r68 2 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.235 $X2=5.59 $Y2=0.39
r69 2 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.235 $X2=5.59 $Y2=0.73
r70 1 17 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%A_27_47# 1 2 3 10 14 15 16 20
r42 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.955 $Y=0.725
+ $X2=1.955 $Y2=0.39
r43 17 25 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0.815
+ $X2=1.155 $Y2=0.815
r44 16 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.79 $Y=0.815
+ $X2=1.955 $Y2=0.725
r45 16 17 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.79 $Y=0.815
+ $X2=1.28 $Y2=0.815
r46 15 25 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=0.725
+ $X2=1.155 $Y2=0.815
r47 14 23 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.155 $Y=0.475
+ $X2=1.155 $Y2=0.365
r48 14 15 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.155 $Y=0.475
+ $X2=1.155 $Y2=0.725
r49 10 23 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0.365
+ $X2=1.155 $Y2=0.365
r50 10 12 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=1.03 $Y=0.365
+ $X2=0.275 $Y2=0.365
r51 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.82
+ $Y=0.235 $X2=1.955 $Y2=0.39
r52 2 25 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.115 $Y2=0.73
r53 2 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.115 $Y2=0.39
r54 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 39 40 41 63 64
r88 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r89 61 64 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r90 60 63 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r91 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r92 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r93 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r94 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r95 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r96 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r97 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r98 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r99 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r100 44 48 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r101 41 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r102 41 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r103 39 57 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=3.91 $Y2=0
r104 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.23
+ $Y2=0
r105 38 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r106 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.23
+ $Y2=0
r107 36 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=2.99
+ $Y2=0
r108 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.355
+ $Y2=0
r109 35 57 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.91
+ $Y2=0
r110 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.355
+ $Y2=0
r111 33 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.07
+ $Y2=0
r112 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.515
+ $Y2=0
r113 32 54 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.99
+ $Y2=0
r114 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.515
+ $Y2=0
r115 30 48 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.15
+ $Y2=0
r116 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.535
+ $Y2=0
r117 29 51 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=2.07
+ $Y2=0
r118 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.535
+ $Y2=0
r119 25 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0
r120 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0.39
r121 21 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0
r122 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0.39
r123 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r124 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.39
r125 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0
r126 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.535 $Y=0.085
+ $X2=1.535 $Y2=0.39
r127 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.23 $Y2=0.39
r128 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.235 $X2=3.355 $Y2=0.39
r129 2 19 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.37
+ $Y=0.235 $X2=2.515 $Y2=0.39
r130 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.235 $X2=1.535 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__XNOR2_2%A_560_47# 1 2 3 12 14 15 18 22 24 25
r56 24 25 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=0.775
+ $X2=5.005 $Y2=0.775
r57 21 22 8.8761 $w=1.8e-07 $l=1.83e-07 $layer=LI1_cond $X=3.975 $Y=0.815
+ $X2=3.792 $Y2=0.815
r58 21 25 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=3.975 $Y=0.815
+ $X2=5.005 $Y2=0.815
r59 16 22 1.0296 $w=3.65e-07 $l=9e-08 $layer=LI1_cond $X=3.792 $Y=0.725
+ $X2=3.792 $Y2=0.815
r60 16 18 10.5772 $w=3.63e-07 $l=3.35e-07 $layer=LI1_cond $X=3.792 $Y=0.725
+ $X2=3.792 $Y2=0.39
r61 14 22 8.8761 $w=1.8e-07 $l=1.82e-07 $layer=LI1_cond $X=3.61 $Y=0.815
+ $X2=3.792 $Y2=0.815
r62 14 15 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.61 $Y=0.815
+ $X2=3.1 $Y2=0.815
r63 10 15 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.935 $Y=0.725
+ $X2=3.1 $Y2=0.815
r64 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.935 $Y=0.725
+ $X2=2.935 $Y2=0.39
r65 3 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.035
+ $Y=0.235 $X2=5.17 $Y2=0.73
r66 2 18 91 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_NDIFF $count=2 $X=3.64
+ $Y=0.235 $X2=3.81 $Y2=0.39
r67 1 12 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.39
.ends


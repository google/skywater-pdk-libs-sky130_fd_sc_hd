* File: sky130_fd_sc_hd__a21oi_2.pxi.spice
* Created: Thu Aug 27 14:01:22 2020
* 
x_PM_SKY130_FD_SC_HD__A21OI_2%A2 N_A2_c_56_n N_A2_M1002_g N_A2_M1001_g
+ N_A2_M1003_g N_A2_M1005_g N_A2_c_71_p N_A2_c_58_n N_A2_c_59_n N_A2_c_60_n A2
+ N_A2_c_61_n N_A2_c_62_n PM_SKY130_FD_SC_HD__A21OI_2%A2
x_PM_SKY130_FD_SC_HD__A21OI_2%A1 N_A1_c_136_n N_A1_M1000_g N_A1_M1006_g
+ N_A1_c_137_n N_A1_M1009_g N_A1_M1008_g A1 N_A1_c_138_n N_A1_c_139_n
+ PM_SKY130_FD_SC_HD__A21OI_2%A1
x_PM_SKY130_FD_SC_HD__A21OI_2%B1 N_B1_M1004_g N_B1_M1010_g N_B1_M1007_g
+ N_B1_M1011_g N_B1_c_189_n B1 B1 N_B1_c_191_n PM_SKY130_FD_SC_HD__A21OI_2%B1
x_PM_SKY130_FD_SC_HD__A21OI_2%A_27_297# N_A_27_297#_M1002_d N_A_27_297#_M1006_s
+ N_A_27_297#_M1005_d N_A_27_297#_M1011_d N_A_27_297#_c_234_n
+ N_A_27_297#_c_235_n N_A_27_297#_c_243_n N_A_27_297#_c_273_p
+ N_A_27_297#_c_246_n N_A_27_297#_c_248_n N_A_27_297#_c_250_n
+ N_A_27_297#_c_236_n N_A_27_297#_c_251_n N_A_27_297#_c_237_n
+ N_A_27_297#_c_252_n PM_SKY130_FD_SC_HD__A21OI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__A21OI_2%VPWR N_VPWR_M1002_s N_VPWR_M1008_d N_VPWR_c_292_n
+ N_VPWR_c_293_n VPWR N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n
+ N_VPWR_c_291_n N_VPWR_c_298_n N_VPWR_c_299_n PM_SKY130_FD_SC_HD__A21OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A21OI_2%Y N_Y_M1000_d N_Y_M1004_d N_Y_M1010_s N_Y_c_345_n
+ N_Y_c_347_n N_Y_c_350_n N_Y_c_343_n N_Y_c_369_n Y N_Y_c_370_n
+ PM_SKY130_FD_SC_HD__A21OI_2%Y
x_PM_SKY130_FD_SC_HD__A21OI_2%VGND N_VGND_M1001_s N_VGND_M1003_s N_VGND_M1007_s
+ N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n VGND N_VGND_c_398_n N_VGND_c_399_n
+ PM_SKY130_FD_SC_HD__A21OI_2%VGND
cc_1 VNB N_A2_c_56_n 0.027828f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.305
cc_2 VNB N_A2_M1001_g 0.0238696f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_3 VNB N_A2_c_58_n 8.46397e-19 $X=-0.19 $Y=-0.24 $X2=1.767 $Y2=1.495
cc_4 VNB N_A2_c_59_n 0.00305053f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_5 VNB N_A2_c_60_n 0.0192728f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_6 VNB N_A2_c_61_n 0.0160618f $X=-0.19 $Y=-0.24 $X2=0.4 $Y2=1.16
cc_7 VNB N_A2_c_62_n 0.0161891f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=0.995
cc_8 VNB N_A1_c_136_n 0.0163968f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.305
cc_9 VNB N_A1_c_137_n 0.0157491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A1_c_138_n 0.00455563f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_11 VNB N_A1_c_139_n 0.030863f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_12 VNB N_B1_M1004_g 0.0177296f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_13 VNB N_B1_M1007_g 0.0225381f $X=-0.19 $Y=-0.24 $X2=1.71 $Y2=0.56
cc_14 VNB N_B1_c_189_n 0.0250418f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.585
cc_15 VNB B1 0.00340572f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_16 VNB N_B1_c_191_n 0.0436892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_291_n 0.136896f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_18 VNB N_Y_c_343_n 0.00125468f $X=-0.19 $Y=-0.24 $X2=1.767 $Y2=1.245
cc_19 VNB N_VGND_c_391_n 0.0110651f $X=-0.19 $Y=-0.24 $X2=1.71 $Y2=0.56
cc_20 VNB N_VGND_c_392_n 0.030637f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.325
cc_21 VNB N_VGND_c_393_n 0.0028319f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=1.585
cc_22 VNB N_VGND_c_394_n 0.0115788f $X=-0.19 $Y=-0.24 $X2=1.767 $Y2=1.245
cc_23 VNB N_VGND_c_395_n 0.0290736f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_24 VNB N_VGND_c_396_n 0.0367309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_397_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.245
cc_26 VNB N_VGND_c_398_n 0.0182775f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.53
cc_27 VNB N_VGND_c_399_n 0.180115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_A2_c_56_n 0.00514747f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.305
cc_29 VPB N_A2_M1002_g 0.023393f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_30 VPB N_A2_M1005_g 0.0172688f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_31 VPB N_A2_c_58_n 0.00325856f $X=-0.19 $Y=1.305 $X2=1.767 $Y2=1.495
cc_32 VPB N_A2_c_60_n 0.00439782f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_33 VPB N_A2_c_61_n 0.00896505f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.16
cc_34 VPB N_A1_M1006_g 0.0187884f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.56
cc_35 VPB N_A1_M1008_g 0.0189179f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_36 VPB N_A1_c_138_n 2.41965e-19 $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_37 VPB N_A1_c_139_n 0.00485795f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_38 VPB N_B1_M1010_g 0.0197171f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.56
cc_39 VPB N_B1_M1011_g 0.0222682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_B1_c_189_n 0.00257374f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.585
cc_41 VPB B1 0.0131786f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_42 VPB N_B1_c_191_n 0.0150524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_297#_c_234_n 0.0113777f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_44 VPB N_A_27_297#_c_235_n 0.0134872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_236_n 0.00795084f $X=-0.19 $Y=1.305 $X2=0.402 $Y2=1.16
cc_46 VPB N_A_27_297#_c_237_n 0.0192814f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=0.995
cc_47 VPB N_VPWR_c_292_n 4.11703e-19 $X=-0.19 $Y=1.305 $X2=1.71 $Y2=0.995
cc_48 VPB N_VPWR_c_293_n 0.00407289f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.985
cc_49 VPB N_VPWR_c_294_n 0.0150591f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.585
cc_50 VPB N_VPWR_c_295_n 0.0147069f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_51 VPB N_VPWR_c_296_n 0.0392278f $X=-0.19 $Y=1.305 $X2=0.4 $Y2=1.16
cc_52 VPB N_VPWR_c_291_n 0.0462919f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_53 VPB N_VPWR_c_298_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_299_n 0.00323844f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.585
cc_55 VPB N_Y_c_343_n 0.00138898f $X=-0.19 $Y=1.305 $X2=1.767 $Y2=1.245
cc_56 N_A2_M1001_g N_A1_c_136_n 0.0401357f $X=0.495 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_57 N_A2_M1002_g N_A1_M1006_g 0.0437939f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A2_c_71_p N_A1_M1006_g 0.0103426f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_59 N_A2_c_61_n N_A1_M1006_g 0.00437137f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A2_c_62_n N_A1_c_137_n 0.0387062f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A2_M1005_g N_A1_M1008_g 0.045988f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A2_c_71_p N_A1_M1008_g 0.0107822f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_63 N_A2_c_56_n N_A1_c_138_n 3.15434e-19 $X=0.49 $Y=1.305 $X2=0 $Y2=0
cc_64 N_A2_M1001_g N_A1_c_138_n 2.57604e-19 $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_65 N_A2_c_71_p N_A1_c_138_n 0.0392259f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_66 N_A2_c_59_n N_A1_c_138_n 0.0197969f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A2_c_60_n N_A1_c_138_n 8.4532e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A2_c_61_n N_A1_c_138_n 0.0248345f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A2_c_56_n N_A1_c_139_n 0.00155214f $X=0.49 $Y=1.305 $X2=0 $Y2=0
cc_70 N_A2_M1001_g N_A1_c_139_n 0.0160113f $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_71 N_A2_c_71_p N_A1_c_139_n 0.00224497f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_72 N_A2_c_58_n N_A1_c_139_n 0.00392425f $X=1.767 $Y=1.495 $X2=0 $Y2=0
cc_73 N_A2_c_59_n N_A1_c_139_n 8.25011e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A2_c_60_n N_A1_c_139_n 0.0387062f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A2_c_61_n N_A1_c_139_n 0.0010512f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A2_c_60_n N_B1_M1004_g 0.0219204f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A2_c_62_n N_B1_M1004_g 0.0218321f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A2_M1005_g N_B1_M1010_g 0.0289349f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A2_c_71_p N_B1_M1010_g 0.0016751f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_80 N_A2_c_58_n N_B1_c_189_n 0.00206837f $X=1.767 $Y=1.495 $X2=0 $Y2=0
cc_81 N_A2_c_59_n N_B1_c_189_n 0.00148742f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A2_c_61_n N_A_27_297#_M1002_d 0.0115922f $X=0.4 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A2_c_71_p N_A_27_297#_M1006_s 0.0033536f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_84 N_A2_c_71_p N_A_27_297#_M1005_d 0.00252765f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_85 N_A2_c_56_n N_A_27_297#_c_234_n 4.73008e-19 $X=0.49 $Y=1.305 $X2=0 $Y2=0
cc_86 N_A2_c_61_n N_A_27_297#_c_234_n 0.0180812f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A2_M1002_g N_A_27_297#_c_243_n 0.0115953f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A2_c_71_p N_A_27_297#_c_243_n 0.0203099f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_89 N_A2_c_61_n N_A_27_297#_c_243_n 0.0128715f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A2_M1005_g N_A_27_297#_c_246_n 0.00837828f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A2_c_71_p N_A_27_297#_c_246_n 0.0293958f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_92 N_A2_M1005_g N_A_27_297#_c_248_n 8.93985e-19 $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A2_c_71_p N_A_27_297#_c_248_n 0.00467621f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_94 N_A2_M1005_g N_A_27_297#_c_250_n 0.00409646f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A2_M1005_g N_A_27_297#_c_251_n 0.00213389f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A2_c_71_p N_A_27_297#_c_252_n 0.0128761f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_97 N_A2_c_71_p N_VPWR_M1002_s 0.0074785f $X=1.605 $Y=1.585 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A2_c_61_n N_VPWR_M1002_s 8.3234e-19 $X=0.4 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_99 N_A2_c_71_p N_VPWR_M1008_d 0.00638346f $X=1.605 $Y=1.585 $X2=0 $Y2=0
cc_100 N_A2_M1002_g N_VPWR_c_292_n 0.00785369f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A2_M1005_g N_VPWR_c_293_n 0.00268723f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A2_M1002_g N_VPWR_c_294_n 0.00351072f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_VPWR_c_296_n 0.00418507f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A2_M1002_g N_VPWR_c_291_n 0.00501961f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A2_M1005_g N_VPWR_c_291_n 0.00572068f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A2_M1001_g N_Y_c_345_n 0.00110268f $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A2_c_62_n N_Y_c_345_n 0.0013659f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A2_c_59_n N_Y_c_347_n 0.0146866f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A2_c_60_n N_Y_c_347_n 0.00275815f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A2_c_62_n N_Y_c_347_n 0.0119595f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A2_M1001_g N_Y_c_350_n 5.19255e-19 $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A2_c_58_n N_Y_c_343_n 0.0111251f $X=1.767 $Y=1.495 $X2=0 $Y2=0
cc_113 N_A2_c_59_n N_Y_c_343_n 0.00733837f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A2_c_60_n N_Y_c_343_n 4.88086e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A2_c_56_n N_VGND_c_392_n 0.00359819f $X=0.49 $Y=1.305 $X2=0 $Y2=0
cc_116 N_A2_M1001_g N_VGND_c_392_n 0.00474835f $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A2_c_61_n N_VGND_c_392_n 0.0205819f $X=0.4 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A2_c_62_n N_VGND_c_393_n 0.0084534f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A2_M1001_g N_VGND_c_396_n 0.00585385f $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_120 N_A2_c_62_n N_VGND_c_396_n 0.00351072f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A2_M1001_g N_VGND_c_399_n 0.0115687f $X=0.495 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A2_c_62_n N_VGND_c_399_n 0.00395482f $X=1.77 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A1_M1006_g N_A_27_297#_c_243_n 0.0116015f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A1_M1008_g N_A_27_297#_c_246_n 0.0100175f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A1_M1008_g N_A_27_297#_c_250_n 4.78112e-19 $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A1_M1006_g N_VPWR_c_292_n 0.00643202f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A1_M1008_g N_VPWR_c_292_n 5.31014e-19 $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A1_M1008_g N_VPWR_c_293_n 0.00139158f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A1_M1006_g N_VPWR_c_295_n 0.00351072f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A1_M1008_g N_VPWR_c_295_n 0.00433717f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A1_M1006_g N_VPWR_c_291_n 0.0040731f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A1_M1008_g N_VPWR_c_291_n 0.00586678f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A1_c_136_n N_Y_c_345_n 0.00711674f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A1_c_137_n N_Y_c_345_n 0.00615696f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A1_c_137_n N_Y_c_347_n 0.00812647f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A1_c_138_n N_Y_c_347_n 0.00750973f $X=1.29 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_c_136_n N_Y_c_350_n 0.00383391f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A1_c_137_n N_Y_c_350_n 7.52978e-19 $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_138_n N_Y_c_350_n 0.0192671f $X=1.29 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A1_c_139_n N_Y_c_350_n 0.0022587f $X=1.35 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A1_c_137_n N_VGND_c_393_n 0.00173186f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_136_n N_VGND_c_396_n 0.00526178f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_137_n N_VGND_c_396_n 0.0041289f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_136_n N_VGND_c_399_n 0.00939774f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_c_137_n N_VGND_c_399_n 0.00557866f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_146 B1 N_A_27_297#_M1011_d 0.00579253f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_147 N_B1_M1010_g N_A_27_297#_c_248_n 0.00326762f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B1_M1010_g N_A_27_297#_c_250_n 0.00420773f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B1_M1011_g N_A_27_297#_c_250_n 4.612e-19 $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B1_M1010_g N_A_27_297#_c_236_n 0.0103776f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B1_M1011_g N_A_27_297#_c_236_n 0.0139439f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B1_M1010_g N_A_27_297#_c_251_n 7.39973e-19 $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B1_M1011_g N_A_27_297#_c_237_n 0.0113733f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_154 B1 N_A_27_297#_c_237_n 0.0245501f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_155 N_B1_c_191_n N_A_27_297#_c_237_n 0.00201808f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B1_M1010_g N_VPWR_c_296_n 0.00357835f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B1_M1011_g N_VPWR_c_296_n 0.00357877f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B1_M1010_g N_VPWR_c_291_n 0.00525234f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B1_M1011_g N_VPWR_c_291_n 0.00636899f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B1_M1004_g N_Y_c_347_n 0.014506f $X=2.19 $Y=0.56 $X2=0 $Y2=0
cc_161 N_B1_M1004_g N_Y_c_343_n 0.00343708f $X=2.19 $Y=0.56 $X2=0 $Y2=0
cc_162 N_B1_M1010_g N_Y_c_343_n 0.00191308f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_163 N_B1_M1007_g N_Y_c_343_n 0.0100221f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_164 N_B1_M1011_g N_Y_c_343_n 0.0200094f $X=2.61 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B1_c_189_n N_Y_c_343_n 0.0210389f $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_166 B1 N_Y_c_343_n 0.044347f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_167 N_B1_M1007_g N_Y_c_369_n 0.00248656f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_168 N_B1_M1007_g N_Y_c_370_n 0.0059052f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_169 N_B1_M1004_g N_VGND_c_393_n 0.00311401f $X=2.19 $Y=0.56 $X2=0 $Y2=0
cc_170 N_B1_M1007_g N_VGND_c_395_n 0.0168464f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_171 B1 N_VGND_c_395_n 0.0249504f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_172 N_B1_c_191_n N_VGND_c_395_n 0.00402147f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_173 N_B1_M1004_g N_VGND_c_398_n 0.00422112f $X=2.19 $Y=0.56 $X2=0 $Y2=0
cc_174 N_B1_M1007_g N_VGND_c_398_n 0.00465454f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_175 N_B1_M1004_g N_VGND_c_399_n 0.00572598f $X=2.19 $Y=0.56 $X2=0 $Y2=0
cc_176 N_B1_M1007_g N_VGND_c_399_n 0.00895587f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_27_297#_c_243_n N_VPWR_M1002_s 0.00353311f $X=1.05 $Y=1.98 $X2=-0.19
+ $Y2=1.305
cc_178 N_A_27_297#_c_246_n N_VPWR_M1008_d 0.00326959f $X=1.815 $Y=1.94 $X2=0
+ $Y2=0
cc_179 N_A_27_297#_c_243_n N_VPWR_c_292_n 0.0163189f $X=1.05 $Y=1.98 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_246_n N_VPWR_c_293_n 0.012114f $X=1.815 $Y=1.94 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_235_n N_VPWR_c_294_n 0.0176542f $X=0.275 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_243_n N_VPWR_c_294_n 0.00264265f $X=1.05 $Y=1.98 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_243_n N_VPWR_c_295_n 0.0027458f $X=1.05 $Y=1.98 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_273_p N_VPWR_c_295_n 0.0116518f $X=1.135 $Y=2.3 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_246_n N_VPWR_c_295_n 0.00300834f $X=1.815 $Y=1.94 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_246_n N_VPWR_c_296_n 0.00211912f $X=1.815 $Y=1.94 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_c_236_n N_VPWR_c_296_n 0.0567977f $X=2.785 $Y=2.375 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_c_251_n N_VPWR_c_296_n 0.0189223f $X=2.145 $Y=2.375 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_M1002_d N_VPWR_c_291_n 0.00239704f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_M1006_s N_VPWR_c_291_n 0.00264218f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_M1005_d N_VPWR_c_291_n 0.00215201f $X=1.845 $Y=1.485 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_M1011_d N_VPWR_c_291_n 0.00292111f $X=2.685 $Y=1.485 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_235_n N_VPWR_c_291_n 0.00990784f $X=0.275 $Y=2.3 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_243_n N_VPWR_c_291_n 0.0104634f $X=1.05 $Y=1.98 $X2=0 $Y2=0
cc_195 N_A_27_297#_c_273_p N_VPWR_c_291_n 0.00644138f $X=1.135 $Y=2.3 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_246_n N_VPWR_c_291_n 0.0106736f $X=1.815 $Y=1.94 $X2=0
+ $Y2=0
cc_197 N_A_27_297#_c_236_n N_VPWR_c_291_n 0.0343717f $X=2.785 $Y=2.375 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_251_n N_VPWR_c_291_n 0.012254f $X=2.145 $Y=2.375 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_236_n N_Y_M1010_s 0.00312899f $X=2.785 $Y=2.375 $X2=0 $Y2=0
cc_200 N_A_27_297#_c_236_n N_Y_c_343_n 0.0175943f $X=2.785 $Y=2.375 $X2=0 $Y2=0
cc_201 N_A_27_297#_c_237_n N_Y_c_343_n 0.024516f $X=2.92 $Y=1.96 $X2=0 $Y2=0
cc_202 N_VPWR_c_291_n N_Y_M1010_s 0.00216833f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_203 N_Y_c_347_n N_VGND_M1003_s 0.00798906f $X=2.295 $Y=0.7 $X2=0 $Y2=0
cc_204 N_Y_c_345_n N_VGND_c_393_n 0.0063786f $X=1.135 $Y=0.36 $X2=0 $Y2=0
cc_205 N_Y_c_347_n N_VGND_c_393_n 0.0180367f $X=2.295 $Y=0.7 $X2=0 $Y2=0
cc_206 N_Y_c_343_n N_VGND_c_395_n 0.0029149f $X=2.4 $Y=1.61 $X2=0 $Y2=0
cc_207 N_Y_c_369_n N_VGND_c_395_n 0.0133992f $X=2.4 $Y=0.76 $X2=0 $Y2=0
cc_208 N_Y_c_370_n N_VGND_c_395_n 0.0266427f $X=2.4 $Y=0.42 $X2=0 $Y2=0
cc_209 N_Y_c_345_n N_VGND_c_396_n 0.0196639f $X=1.135 $Y=0.36 $X2=0 $Y2=0
cc_210 N_Y_c_347_n N_VGND_c_396_n 0.00720366f $X=2.295 $Y=0.7 $X2=0 $Y2=0
cc_211 N_Y_c_347_n N_VGND_c_398_n 0.00312282f $X=2.295 $Y=0.7 $X2=0 $Y2=0
cc_212 N_Y_c_370_n N_VGND_c_398_n 0.0192685f $X=2.4 $Y=0.42 $X2=0 $Y2=0
cc_213 N_Y_M1000_d N_VGND_c_399_n 0.00223231f $X=0.995 $Y=0.235 $X2=0 $Y2=0
cc_214 N_Y_M1004_d N_VGND_c_399_n 0.00224147f $X=2.265 $Y=0.235 $X2=0 $Y2=0
cc_215 N_Y_c_345_n N_VGND_c_399_n 0.0126929f $X=1.135 $Y=0.36 $X2=0 $Y2=0
cc_216 N_Y_c_347_n N_VGND_c_399_n 0.0185643f $X=2.295 $Y=0.7 $X2=0 $Y2=0
cc_217 N_Y_c_370_n N_VGND_c_399_n 0.0118083f $X=2.4 $Y=0.42 $X2=0 $Y2=0
cc_218 N_Y_c_347_n A_114_47# 0.00529826f $X=2.295 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_219 N_VGND_c_399_n A_285_47# 0.011755f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_220 N_VGND_c_399_n A_114_47# 0.00239227f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a31o_4.spice
* Created: Thu Aug 27 14:04:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a31o_4.spice.pex"
.subckt sky130_fd_sc_hd__a31o_4  VNB VPB A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A3_M1021_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.2 SB=75005.4
+ A=0.0975 P=1.6 MULT=1
MM1008 A_109_47# N_A2_M1008_g A_193_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=14.76 M=1 R=4.33333 SA=75000.6
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1011 A_193_47# N_A1_M1011_g N_A_277_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75004.6 A=0.0975 P=1.6 MULT=1
MM1010 A_361_47# N_A1_M1010_g N_A_277_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1018 A_445_47# N_A2_M1018_g A_361_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75001.9
+ SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A3_M1023_g A_445_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.10725 PD=0.98 PS=0.98 NRD=6.456 NRS=20.304 M=1 R=4.33333 SA=75002.3
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1004 N_A_277_47#_M1004_d N_B1_M1004_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75002.8
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1022 N_A_277_47#_M1004_d N_B1_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75003.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1022_s N_A_277_47#_M1013_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75004.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A_277_47#_M1015_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1015_d N_A_277_47#_M1016_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1017_d N_A_277_47#_M1017_g N_X_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_297#_M1005_d N_A3_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_297#_M1003_d N_A2_M1003_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_27_297#_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1020 N_VPWR_M1002_d N_A1_M1020_g N_A_27_297#_M1020_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1014 N_A_27_297#_M1020_s N_A2_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.165 PD=1.27 PS=1.33 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_27_297#_M1012_d N_A3_M1012_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.165 PD=1.33 PS=1.33 NRD=10.8153 NRS=10.8153 M=1 R=6.66667
+ SA=75002.3 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1000 N_A_277_47#_M1000_d N_B1_M1000_g N_A_27_297#_M1012_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.165 PD=1.27 PS=1.33 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1006 N_A_277_47#_M1000_d N_B1_M1006_g N_A_27_297#_M1006_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_277_47#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1001_d N_A_277_47#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1009 N_X_M1009_d N_A_277_47#_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1019 N_X_M1009_d N_A_277_47#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.5 PD=1.27 PS=3 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.4
+ A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_53 VNB 0 1.75522e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__a31o_4.spice.SKY130_FD_SC_HD__A31O_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__o211a_1.spice.pex
* Created: Thu Aug 27 14:34:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211A_1%A_79_21# 1 2 3 12 16 18 21 24 25 26 29 31 34
+ 37 40 42 46
c88 24 0 1.31813e-19 $X=1.04 $Y=1.495
c89 18 0 1.55223e-20 $X=0.955 $Y=1.16
r90 42 44 17.172 $w=4.98e-07 $l=4.85e-07 $layer=LI1_cond $X=3.14 $Y=0.38
+ $X2=3.14 $Y2=0.865
r91 35 46 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=1.665
+ $X2=3.14 $Y2=1.58
r92 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.225 $Y=1.665
+ $X2=3.225 $Y2=2.34
r93 34 46 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.975 $Y=1.495
+ $X2=3.14 $Y2=1.58
r94 34 44 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.975 $Y=1.495
+ $X2=2.975 $Y2=0.865
r95 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=1.58
+ $X2=2.095 $Y2=1.58
r96 31 46 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=1.58 $X2=3.14
+ $Y2=1.58
r97 31 32 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.89 $Y=1.58
+ $X2=2.26 $Y2=1.58
r98 27 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=1.665
+ $X2=2.095 $Y2=1.58
r99 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.095 $Y=1.665
+ $X2=2.095 $Y2=2.34
r100 25 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=1.58
+ $X2=2.095 $Y2=1.58
r101 25 26 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.93 $Y=1.58
+ $X2=1.125 $Y2=1.58
r102 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.04 $Y=1.495
+ $X2=1.125 $Y2=1.58
r103 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.04 $Y=1.245
+ $X2=1.04 $Y2=1.495
r104 21 47 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.47 $Y2=1.16
r105 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r106 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.955 $Y=1.16
+ $X2=1.04 $Y2=1.245
r107 18 20 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.955 $Y=1.16
+ $X2=0.595 $Y2=1.16
r108 14 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.16
r109 14 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.47 $Y=1.295
+ $X2=0.47 $Y2=1.985
r110 10 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.16
r111 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
r112 3 46 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.485 $X2=3.225 $Y2=1.66
r113 3 37 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.485 $X2=3.225 $Y2=2.34
r114 2 40 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.485 $X2=2.095 $Y2=1.66
r115 2 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.485 $X2=2.095 $Y2=2.34
r116 1 42 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=3.05
+ $Y=0.235 $X2=3.225 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%A1 3 6 8 11 13
c36 11 0 3.01083e-19 $X=1.465 $Y=1.16
r37 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=1.325
r38 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.16
+ $X2=1.465 $Y2=0.995
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.16 $X2=1.465 $Y2=1.16
r40 8 12 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.635 $Y=1.175
+ $X2=1.465 $Y2=1.175
r41 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.985
+ $X2=1.41 $Y2=1.325
r42 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.56 $X2=1.41
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%A2 3 6 8 11 13
c32 11 0 1.55223e-20 $X=2.055 $Y=1.16
c33 8 0 1.73117e-19 $X=2.095 $Y=1.19
r34 11 14 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.16 $X2=2
+ $Y2=1.325
r35 11 13 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.16 $X2=2
+ $Y2=0.995
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.16 $X2=2.055 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.885 $Y=1.985
+ $X2=1.885 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.885 $Y=0.56
+ $X2=1.885 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%B1 3 6 8 11 13
r30 11 14 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.16
+ $X2=2.545 $Y2=1.325
r31 11 13 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.16
+ $X2=2.545 $Y2=0.995
r32 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.555
+ $Y=1.16 $X2=2.555 $Y2=1.16
r33 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.475 $Y=1.985
+ $X2=2.475 $Y2=1.325
r34 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.475 $Y=0.56
+ $X2=2.475 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%C1 1 3 6 9 10 13
r28 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.16 $X2=3.41 $Y2=1.16
r29 8 13 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.05 $Y=1.16 $X2=3.41
+ $Y2=1.16
r30 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.05 $Y=1.16 $X2=2.975
+ $Y2=1.16
r31 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.325
+ $X2=2.975 $Y2=1.16
r32 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.975 $Y=1.325
+ $X2=2.975 $Y2=1.985
r33 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=0.995
+ $X2=2.975 $Y2=1.16
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.975 $Y=0.995
+ $X2=2.975 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%X 1 2 10 13 14 15 16 17 22
r18 17 31 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=2.21
+ $X2=0.255 $Y2=2.34
r19 16 17 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.255 $Y=1.87
+ $X2=0.255 $Y2=2.21
r20 15 22 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.51
+ $X2=0.255 $Y2=0.38
r21 13 14 8.29786 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=1.495
r22 11 16 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.87
r23 11 13 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.66
r24 10 14 38.6597 $w=1.73e-07 $l=6.1e-07 $layer=LI1_cond $X=0.172 $Y=0.885
+ $X2=0.172 $Y2=1.495
r25 9 15 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.51
r26 9 10 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.885
r27 2 31 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r28 2 13 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r29 1 22 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%VPWR 1 2 3 12 16 20 24 27 28 29 31 44 45 48
+ 51
c46 2 0 1.31813e-19 $X=1.075 $Y=1.485
r47 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 49 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r53 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r55 38 41 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 36 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.16 $Y2=2.72
r58 36 38 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 31 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r60 31 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r61 29 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 27 41 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.56 $Y=2.72 $X2=2.53
+ $Y2=2.72
r64 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=2.72
+ $X2=2.725 $Y2=2.72
r65 26 44 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=2.72
+ $X2=2.725 $Y2=2.72
r67 22 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=2.635
+ $X2=2.725 $Y2=2.72
r68 22 24 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.725 $Y=2.635
+ $X2=2.725 $Y2=2
r69 18 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=2.635
+ $X2=1.16 $Y2=2.72
r70 18 20 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.16 $Y=2.635
+ $X2=1.16 $Y2=2
r71 17 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r72 16 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.16 $Y2=2.72
r73 16 17 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.765 $Y2=2.72
r74 12 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.66
+ $X2=0.68 $Y2=2.34
r75 10 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r76 10 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r77 3 24 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.485 $X2=2.725 $Y2=2
r78 2 20 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2
r79 1 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r80 1 12 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%VGND 1 2 9 11 15 17 19 29 30 33 36
r44 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r45 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r46 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r49 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r50 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r51 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r52 24 36 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.76 $Y=0 $X2=1.647
+ $Y2=0
r53 24 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.76 $Y=0 $X2=2.07
+ $Y2=0
r54 19 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.72
+ $Y2=0
r55 19 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r56 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 13 36 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.647 $Y=0.085
+ $X2=1.647 $Y2=0
r59 13 15 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.647 $Y=0.085
+ $X2=1.647 $Y2=0.38
r60 12 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.72
+ $Y2=0
r61 11 36 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.647
+ $Y2=0
r62 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=0.845
+ $Y2=0
r63 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r64 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r65 2 15 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.65 $Y2=0.38
r66 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_1%A_215_47# 1 2 9 11 12 15
c36 12 0 1.27966e-19 $X=1.365 $Y=0.82
r37 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.095 $Y=0.735
+ $X2=2.095 $Y2=0.38
r38 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.93 $Y=0.82
+ $X2=2.095 $Y2=0.735
r39 11 12 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.93 $Y=0.82
+ $X2=1.365 $Y2=0.82
r40 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.365 $Y2=0.82
r41 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.2 $Y=0.735 $X2=1.2
+ $Y2=0.38
r42 2 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=0.235 $X2=2.095 $Y2=0.38
r43 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends


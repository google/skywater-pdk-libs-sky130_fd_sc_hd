# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 0.620000 1.305000 0.995000 ;
        RECT 0.970000 0.995000 1.430000 1.325000 ;
        RECT 0.970000 1.325000 1.305000 1.695000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 9.575000 1.725000 ;
        RECT 6.275000 0.615000 9.575000 0.855000 ;
        RECT 9.325000 0.855000 9.575000 1.445000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.660000 0.085000 ;
        RECT 0.085000  0.085000 0.445000 0.825000 ;
        RECT 0.970000  0.085000 1.305000 0.445000 ;
        RECT 2.655000  0.085000 2.985000 0.485000 ;
        RECT 3.495000  0.085000 3.825000 0.485000 ;
        RECT 4.335000  0.085000 4.665000 0.485000 ;
        RECT 5.175000  0.085000 5.505000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.660000 2.805000 ;
        RECT 0.085000 1.785000 0.445000 2.635000 ;
        RECT 0.970000 1.865000 1.305000 2.635000 ;
        RECT 2.415000 2.235000 2.745000 2.635000 ;
        RECT 3.255000 2.235000 3.585000 2.635000 ;
        RECT 4.095000 2.235000 4.425000 2.635000 ;
        RECT 4.935000 2.235000 5.265000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.600000 0.995000 0.800000 1.615000 ;
      RECT 0.615000 0.280000 0.800000 0.995000 ;
      RECT 0.615000 1.615000 0.800000 2.465000 ;
      RECT 1.475000 0.255000 1.985000 0.825000 ;
      RECT 1.475000 1.495000 1.825000 2.465000 ;
      RECT 1.600000 0.825000 1.985000 1.025000 ;
      RECT 1.600000 1.025000 5.925000 1.275000 ;
      RECT 1.600000 1.275000 1.825000 1.495000 ;
      RECT 1.995000 1.895000 9.575000 2.065000 ;
      RECT 1.995000 2.065000 2.245000 2.465000 ;
      RECT 2.155000 0.255000 2.485000 0.655000 ;
      RECT 2.155000 0.655000 6.105000 0.855000 ;
      RECT 2.915000 2.065000 3.085000 2.465000 ;
      RECT 3.155000 0.275000 3.325000 0.655000 ;
      RECT 3.755000 2.065000 3.925000 2.465000 ;
      RECT 3.995000 0.255000 4.165000 0.655000 ;
      RECT 4.595000 2.065000 4.765000 2.465000 ;
      RECT 4.835000 0.275000 5.005000 0.655000 ;
      RECT 5.435000 2.065000 9.575000 2.465000 ;
      RECT 5.675000 0.255000 9.575000 0.445000 ;
      RECT 5.675000 0.445000 6.105000 0.655000 ;
      RECT 6.175000 1.025000 9.155000 1.275000 ;
    LAYER mcon ;
      RECT 0.605000 1.105000 0.775000 1.275000 ;
      RECT 6.580000 1.105000 6.750000 1.275000 ;
    LAYER met1 ;
      RECT 0.545000 1.075000 0.835000 1.120000 ;
      RECT 0.545000 1.120000 6.810000 1.260000 ;
      RECT 0.545000 1.260000 0.835000 1.305000 ;
      RECT 6.520000 1.075000 6.810000 1.120000 ;
      RECT 6.520000 1.260000 6.810000 1.305000 ;
  END
END sky130_fd_sc_hd__ebufn_8
END LIBRARY

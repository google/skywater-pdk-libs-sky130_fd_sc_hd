* File: sky130_fd_sc_hd__nor4b_2.pxi.spice
* Created: Thu Aug 27 14:33:09 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4B_2%A N_A_c_92_n N_A_M1009_g N_A_M1007_g N_A_c_93_n
+ N_A_M1016_g N_A_M1013_g A A A N_A_c_95_n PM_SKY130_FD_SC_HD__NOR4B_2%A
x_PM_SKY130_FD_SC_HD__NOR4B_2%B N_B_c_136_n N_B_M1011_g N_B_M1003_g N_B_c_137_n
+ N_B_M1012_g N_B_M1015_g B B B N_B_c_139_n PM_SKY130_FD_SC_HD__NOR4B_2%B
x_PM_SKY130_FD_SC_HD__NOR4B_2%C N_C_c_179_n N_C_M1004_g N_C_M1010_g N_C_c_180_n
+ N_C_M1005_g N_C_M1014_g C C N_C_c_182_n PM_SKY130_FD_SC_HD__NOR4B_2%C
x_PM_SKY130_FD_SC_HD__NOR4B_2%A_694_21# N_A_694_21#_M1017_s N_A_694_21#_M1008_s
+ N_A_694_21#_c_224_n N_A_694_21#_M1001_g N_A_694_21#_M1000_g
+ N_A_694_21#_c_225_n N_A_694_21#_M1006_g N_A_694_21#_M1002_g
+ N_A_694_21#_c_226_n N_A_694_21#_c_227_n N_A_694_21#_c_228_n
+ N_A_694_21#_c_229_n N_A_694_21#_c_230_n N_A_694_21#_c_236_n
+ N_A_694_21#_c_231_n PM_SKY130_FD_SC_HD__NOR4B_2%A_694_21#
x_PM_SKY130_FD_SC_HD__NOR4B_2%D_N N_D_N_M1017_g N_D_N_M1008_g N_D_N_c_295_n
+ N_D_N_c_296_n D_N D_N D_N N_D_N_c_298_n N_D_N_c_299_n
+ PM_SKY130_FD_SC_HD__NOR4B_2%D_N
x_PM_SKY130_FD_SC_HD__NOR4B_2%A_27_297# N_A_27_297#_M1007_d N_A_27_297#_M1013_d
+ N_A_27_297#_M1015_s N_A_27_297#_c_326_n N_A_27_297#_c_327_n
+ N_A_27_297#_c_328_n N_A_27_297#_c_351_p N_A_27_297#_c_329_n
+ N_A_27_297#_c_330_n N_A_27_297#_c_331_n PM_SKY130_FD_SC_HD__NOR4B_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR4B_2%VPWR N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_c_369_n
+ N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n VPWR
+ N_VPWR_c_374_n N_VPWR_c_368_n N_VPWR_c_376_n PM_SKY130_FD_SC_HD__NOR4B_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR4B_2%A_277_297# N_A_277_297#_M1003_d
+ N_A_277_297#_M1010_s N_A_277_297#_c_430_n N_A_277_297#_c_426_n
+ N_A_277_297#_c_438_n N_A_277_297#_c_444_p
+ PM_SKY130_FD_SC_HD__NOR4B_2%A_277_297#
x_PM_SKY130_FD_SC_HD__NOR4B_2%A_474_297# N_A_474_297#_M1010_d
+ N_A_474_297#_M1014_d N_A_474_297#_M1002_d N_A_474_297#_c_445_n
+ N_A_474_297#_c_446_n N_A_474_297#_c_447_n N_A_474_297#_c_448_n
+ N_A_474_297#_c_470_n N_A_474_297#_c_460_n N_A_474_297#_c_463_n
+ PM_SKY130_FD_SC_HD__NOR4B_2%A_474_297#
x_PM_SKY130_FD_SC_HD__NOR4B_2%Y N_Y_M1009_s N_Y_M1011_s N_Y_M1004_s N_Y_M1001_d
+ N_Y_M1000_s N_Y_c_496_n N_Y_c_486_n N_Y_c_487_n N_Y_c_504_n N_Y_c_488_n
+ N_Y_c_516_n N_Y_c_489_n N_Y_c_520_n N_Y_c_490_n N_Y_c_491_n N_Y_c_492_n Y Y
+ N_Y_c_493_n Y N_Y_c_554_n PM_SKY130_FD_SC_HD__NOR4B_2%Y
x_PM_SKY130_FD_SC_HD__NOR4B_2%VGND N_VGND_M1009_d N_VGND_M1016_d N_VGND_M1012_d
+ N_VGND_M1004_d N_VGND_M1005_d N_VGND_M1006_s N_VGND_M1017_d N_VGND_c_585_n
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n
+ N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n
+ N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n VGND
+ N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n PM_SKY130_FD_SC_HD__NOR4B_2%VGND
cc_1 VNB N_A_c_92_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_93_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB A 0.0210886f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.105
cc_4 VNB N_A_c_95_n 0.0369647f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B_c_136_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_6 VNB N_B_c_137_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_7 VNB B 0.0232054f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.105
cc_8 VNB N_B_c_139_n 0.0369647f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_9 VNB N_C_c_179_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_C_c_180_n 0.015991f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_11 VNB C 0.00523478f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.105
cc_12 VNB N_C_c_182_n 0.0369611f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_13 VNB N_A_694_21#_c_224_n 0.0159884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_694_21#_c_225_n 0.0192233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_694_21#_c_226_n 0.0259551f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_16 VNB N_A_694_21#_c_227_n 0.00263734f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_17 VNB N_A_694_21#_c_228_n 0.00110808f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.18
cc_18 VNB N_A_694_21#_c_229_n 0.0426408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_694_21#_c_230_n 0.0168523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_694_21#_c_231_n 4.62534e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D_N_c_295_n 0.00629781f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_22 VNB N_D_N_c_296_n 0.0265991f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_23 VNB D_N 9.59049e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D_N_c_298_n 0.0213565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_D_N_c_299_n 0.0181249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_368_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_486_n 0.00248283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_487_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_29 VNB N_Y_c_488_n 0.0123035f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_30 VNB N_Y_c_489_n 0.00248283f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.18
cc_31 VNB N_Y_c_490_n 0.00244444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_491_n 0.00244444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_492_n 0.0015406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_493_n 8.38427e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_585_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_586_n 0.0327449f $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=1.16
cc_37 VNB N_VGND_c_587_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.18
cc_38 VNB N_VGND_c_588_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.18
cc_39 VNB N_VGND_c_589_n 0.00677439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_590_n 0.0198702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_591_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_592_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_593_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_594_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_595_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_596_n 0.0039398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_597_n 0.0110534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_598_n 0.0194526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_599_n 0.00480869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_600_n 0.295612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_601_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_602_n 0.0270624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A_M1007_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_A_M1013_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_55 VPB N_A_c_95_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_56 VPB N_B_M1003_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_57 VPB N_B_M1015_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_58 VPB N_B_c_139_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_59 VPB N_C_M1010_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_60 VPB N_C_M1014_g 0.0184813f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_61 VPB N_C_c_182_n 0.00480901f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_62 VPB N_A_694_21#_M1000_g 0.0187825f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_63 VPB N_A_694_21#_M1002_g 0.0220422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_694_21#_c_226_n 0.00412255f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_65 VPB N_A_694_21#_c_229_n 0.0223977f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_694_21#_c_236_n 0.0128805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_694_21#_c_231_n 0.0165053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_D_N_M1008_g 0.0639063f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_69 VPB N_D_N_c_296_n 0.0077491f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_70 VPB D_N 0.0391179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_297#_c_326_n 0.0332602f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_72 VPB N_A_27_297#_c_327_n 0.00226814f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.105
cc_73 VPB N_A_27_297#_c_328_n 0.0103161f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.105
cc_74 VPB N_A_27_297#_c_329_n 0.00688307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_297#_c_330_n 0.0047044f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_76 VPB N_A_27_297#_c_331_n 0.00234762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_369_n 0.00489695f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_78 VPB N_VPWR_c_370_n 0.00517963f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_79 VPB N_VPWR_c_371_n 0.0110534f $X=-0.19 $Y=1.305 $X2=0.13 $Y2=1.105
cc_80 VPB N_VPWR_c_372_n 0.101328f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.105
cc_81 VPB N_VPWR_c_373_n 0.00478242f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.105
cc_82 VPB N_VPWR_c_374_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_368_n 0.0565492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_376_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_277_297#_c_426_n 0.0111956f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_86 VPB N_A_474_297#_c_445_n 0.00608777f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_87 VPB N_A_474_297#_c_446_n 0.00247808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_474_297#_c_447_n 0.00523353f $X=-0.19 $Y=1.305 $X2=0.13 $Y2=1.105
cc_89 VPB N_A_474_297#_c_448_n 0.00257883f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.105
cc_90 VPB Y 0.0012835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB Y 0.00125905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 N_A_c_93_n N_B_c_136_n 0.0195487f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_A_M1013_g N_B_M1003_g 0.0195487f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 A B 0.0168093f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_95 A N_B_c_139_n 0.00573515f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_95_n N_B_c_139_n 0.0195487f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_M1007_g N_A_27_297#_c_326_n 0.0102794f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_M1013_g N_A_27_297#_c_326_n 6.39698e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_M1007_g N_A_27_297#_c_327_n 0.0107189f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_M1013_g N_A_27_297#_c_327_n 0.0132641f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 A N_A_27_297#_c_327_n 0.0389132f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_c_95_n N_A_27_297#_c_327_n 0.00211509f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_M1007_g N_A_27_297#_c_328_n 0.00149004f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_104 A N_A_27_297#_c_328_n 0.0275988f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_105 A N_A_27_297#_c_329_n 0.00107215f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_106 A N_A_27_297#_c_331_n 0.0214236f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VPWR_c_369_n 0.00274642f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1013_g N_VPWR_c_369_n 0.00296718f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_M1013_g N_VPWR_c_372_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_M1007_g N_VPWR_c_374_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1007_g N_VPWR_c_368_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1013_g N_VPWR_c_368_n 0.010464f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_c_92_n N_Y_c_496_n 0.00539651f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_c_93_n N_Y_c_496_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_93_n N_Y_c_486_n 0.00865686f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_116 A N_Y_c_486_n 0.0293675f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A_c_92_n N_Y_c_487_n 0.00262807f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_93_n N_Y_c_487_n 0.00113286f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_119 A N_Y_c_487_n 0.0266272f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A_c_95_n N_Y_c_487_n 0.00230339f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_c_93_n N_Y_c_504_n 5.22228e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_92_n N_VGND_c_586_n 0.00366155f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_123 A N_VGND_c_586_n 0.0209094f $X=1.05 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_c_93_n N_VGND_c_587_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_92_n N_VGND_c_591_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_93_n N_VGND_c_591_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_92_n N_VGND_c_600_n 0.0104557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_93_n N_VGND_c_600_n 0.0057435f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_129 B C 0.0168827f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_130 B N_C_c_182_n 0.00852834f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B_M1003_g N_A_27_297#_c_329_n 0.0150585f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B_M1015_g N_A_27_297#_c_329_n 0.010363f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_133 B N_A_27_297#_c_329_n 0.0533009f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_134 N_B_c_139_n N_A_27_297#_c_329_n 0.00211509f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B_M1003_g N_A_27_297#_c_330_n 5.39745e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B_M1015_g N_A_27_297#_c_330_n 0.00689323f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B_M1003_g N_VPWR_c_372_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B_M1015_g N_VPWR_c_372_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B_M1003_g N_VPWR_c_368_n 0.0106871f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B_M1015_g N_VPWR_c_368_n 0.00660224f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_M1015_g N_A_277_297#_c_426_n 0.0115198f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1015_g N_A_474_297#_c_447_n 3.68548e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_143 B N_A_474_297#_c_447_n 0.0307707f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_144 N_B_c_136_n N_Y_c_496_n 5.22228e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B_c_136_n N_Y_c_486_n 0.0100722f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B_c_136_n N_Y_c_504_n 0.00630972f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_137_n N_Y_c_504_n 0.0109565f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_148 N_B_c_137_n N_Y_c_488_n 0.0109318f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_149 B N_Y_c_488_n 0.0720239f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_150 N_B_c_136_n N_Y_c_490_n 0.00151671f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_137_n N_Y_c_490_n 0.00113286f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_152 B N_Y_c_490_n 0.0214636f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_153 N_B_c_139_n N_Y_c_490_n 0.00230339f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B_c_136_n N_VGND_c_587_n 0.00146339f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B_c_136_n N_VGND_c_600_n 0.0057435f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B_c_137_n N_VGND_c_600_n 0.0070399f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B_c_136_n N_VGND_c_601_n 0.00423334f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B_c_137_n N_VGND_c_601_n 0.00423334f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B_c_137_n N_VGND_c_602_n 0.00336547f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_160 N_C_c_180_n N_A_694_21#_c_224_n 0.0190517f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_161 N_C_M1014_g N_A_694_21#_M1000_g 0.0190517f $X=3.125 $Y=1.985 $X2=0 $Y2=0
cc_162 C N_A_694_21#_c_226_n 0.0106418f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_163 N_C_c_182_n N_A_694_21#_c_226_n 0.0190517f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_164 N_C_M1010_g N_A_27_297#_c_329_n 3.35158e-19 $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_165 N_C_M1010_g N_VPWR_c_372_n 0.00357877f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_166 N_C_M1014_g N_VPWR_c_372_n 0.00585385f $X=3.125 $Y=1.985 $X2=0 $Y2=0
cc_167 N_C_M1010_g N_VPWR_c_368_n 0.00660224f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_168 N_C_M1014_g N_VPWR_c_368_n 0.0106871f $X=3.125 $Y=1.985 $X2=0 $Y2=0
cc_169 N_C_M1010_g N_A_277_297#_c_426_n 0.0115198f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_170 N_C_M1010_g N_A_474_297#_c_445_n 0.00689323f $X=2.705 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_C_M1014_g N_A_474_297#_c_445_n 5.38818e-19 $X=3.125 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_C_M1010_g N_A_474_297#_c_446_n 0.0103205f $X=2.705 $Y=1.985 $X2=0 $Y2=0
cc_173 N_C_M1014_g N_A_474_297#_c_446_n 0.0132131f $X=3.125 $Y=1.985 $X2=0 $Y2=0
cc_174 C N_A_474_297#_c_446_n 0.028136f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_175 N_C_c_182_n N_A_474_297#_c_446_n 0.00211509f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_176 N_C_M1010_g N_A_474_297#_c_447_n 0.00181203f $X=2.705 $Y=1.985 $X2=0
+ $Y2=0
cc_177 C N_A_474_297#_c_448_n 0.0214236f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_178 N_C_c_179_n N_Y_c_488_n 0.0123466f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_179 N_C_c_179_n N_Y_c_516_n 0.0109565f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C_c_180_n N_Y_c_516_n 0.00630972f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_181 N_C_c_180_n N_Y_c_489_n 0.00865686f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_182 C N_Y_c_489_n 0.0335195f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_183 N_C_c_180_n N_Y_c_520_n 5.22228e-19 $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_184 N_C_c_179_n N_Y_c_491_n 0.00151671f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C_c_180_n N_Y_c_491_n 0.00113286f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_186 C N_Y_c_491_n 0.0214636f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_187 N_C_c_182_n N_Y_c_491_n 0.00230339f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_188 C Y 0.0158574f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_189 N_C_c_182_n N_Y_c_493_n 3.69674e-19 $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_190 N_C_c_180_n N_VGND_c_588_n 0.00146339f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_191 N_C_c_179_n N_VGND_c_593_n 0.00423334f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_192 N_C_c_180_n N_VGND_c_593_n 0.00423334f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_193 N_C_c_179_n N_VGND_c_600_n 0.0070399f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_194 N_C_c_180_n N_VGND_c_600_n 0.0057435f $X=3.125 $Y=0.995 $X2=0 $Y2=0
cc_195 N_C_c_179_n N_VGND_c_602_n 0.00336547f $X=2.705 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_694_21#_c_236_n N_D_N_M1008_g 0.00181686f $X=4.695 $Y=2.285 $X2=0
+ $Y2=0
cc_197 N_A_694_21#_c_228_n N_D_N_c_295_n 0.0147859f $X=4.485 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_694_21#_c_229_n N_D_N_c_295_n 7.33016e-19 $X=4.485 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_694_21#_c_230_n N_D_N_c_295_n 0.0011748f $X=4.695 $Y=0.66 $X2=0 $Y2=0
cc_200 N_A_694_21#_c_231_n N_D_N_c_295_n 0.00327196f $X=4.642 $Y=2.035 $X2=0
+ $Y2=0
cc_201 N_A_694_21#_c_228_n N_D_N_c_296_n 5.14425e-19 $X=4.485 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_694_21#_c_229_n N_D_N_c_296_n 0.0211508f $X=4.485 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_694_21#_c_231_n N_D_N_c_296_n 0.0171405f $X=4.642 $Y=2.035 $X2=0
+ $Y2=0
cc_204 N_A_694_21#_c_231_n D_N 0.022806f $X=4.642 $Y=2.035 $X2=0 $Y2=0
cc_205 N_A_694_21#_c_227_n N_D_N_c_298_n 0.00454127f $X=4.55 $Y=1.075 $X2=0
+ $Y2=0
cc_206 N_A_694_21#_c_230_n N_D_N_c_298_n 0.00348716f $X=4.695 $Y=0.66 $X2=0
+ $Y2=0
cc_207 N_A_694_21#_M1000_g N_VPWR_c_372_n 0.00357877f $X=3.545 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_694_21#_M1002_g N_VPWR_c_372_n 0.00357877f $X=3.965 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_694_21#_c_236_n N_VPWR_c_372_n 0.0210237f $X=4.695 $Y=2.285 $X2=0
+ $Y2=0
cc_210 N_A_694_21#_M1008_s N_VPWR_c_368_n 0.00244558f $X=4.57 $Y=2.065 $X2=0
+ $Y2=0
cc_211 N_A_694_21#_M1000_g N_VPWR_c_368_n 0.00525237f $X=3.545 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_694_21#_M1002_g N_VPWR_c_368_n 0.00655123f $X=3.965 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_694_21#_c_236_n N_VPWR_c_368_n 0.0134053f $X=4.695 $Y=2.285 $X2=0
+ $Y2=0
cc_214 N_A_694_21#_M1000_g N_A_474_297#_c_448_n 2.5798e-19 $X=3.545 $Y=1.985
+ $X2=0 $Y2=0
cc_215 N_A_694_21#_M1000_g N_A_474_297#_c_460_n 0.0121306f $X=3.545 $Y=1.985
+ $X2=0 $Y2=0
cc_216 N_A_694_21#_M1002_g N_A_474_297#_c_460_n 0.00991691f $X=3.965 $Y=1.985
+ $X2=0 $Y2=0
cc_217 N_A_694_21#_c_236_n N_A_474_297#_c_460_n 0.0135088f $X=4.695 $Y=2.285
+ $X2=0 $Y2=0
cc_218 N_A_694_21#_c_229_n N_A_474_297#_c_463_n 0.00700853f $X=4.485 $Y=1.16
+ $X2=0 $Y2=0
cc_219 N_A_694_21#_c_231_n N_A_474_297#_c_463_n 0.0390847f $X=4.642 $Y=2.035
+ $X2=0 $Y2=0
cc_220 N_A_694_21#_c_224_n N_Y_c_516_n 5.22228e-19 $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_694_21#_c_224_n N_Y_c_489_n 0.0103201f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_694_21#_c_224_n N_Y_c_520_n 0.00630972f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_694_21#_c_225_n N_Y_c_520_n 0.00539651f $X=3.965 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A_694_21#_c_224_n N_Y_c_492_n 0.00221107f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_694_21#_c_225_n N_Y_c_492_n 0.00230016f $X=3.965 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_694_21#_c_230_n N_Y_c_492_n 3.49029e-19 $X=4.695 $Y=0.66 $X2=0 $Y2=0
cc_227 N_A_694_21#_M1000_g Y 0.00329139f $X=3.545 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_694_21#_M1002_g Y 0.0042161f $X=3.965 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A_694_21#_c_226_n Y 0.0238815f $X=4.04 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_694_21#_c_228_n Y 0.00829564f $X=4.485 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_694_21#_c_231_n Y 0.014002f $X=4.642 $Y=2.035 $X2=0 $Y2=0
cc_232 N_A_694_21#_c_224_n N_Y_c_493_n 0.00208232f $X=3.545 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_694_21#_c_225_n N_Y_c_493_n 0.0024642f $X=3.965 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_694_21#_c_226_n N_Y_c_493_n 0.00701755f $X=4.04 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_694_21#_c_227_n N_Y_c_493_n 0.00477319f $X=4.55 $Y=1.075 $X2=0 $Y2=0
cc_236 N_A_694_21#_M1000_g Y 2.42171e-19 $X=3.545 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_694_21#_M1002_g Y 0.00891195f $X=3.965 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A_694_21#_c_224_n N_VGND_c_588_n 0.00146448f $X=3.545 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A_694_21#_c_225_n N_VGND_c_589_n 0.00340598f $X=3.965 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A_694_21#_c_229_n N_VGND_c_589_n 0.00973477f $X=4.485 $Y=1.16 $X2=0
+ $Y2=0
cc_241 N_A_694_21#_c_230_n N_VGND_c_589_n 0.0409286f $X=4.695 $Y=0.66 $X2=0
+ $Y2=0
cc_242 N_A_694_21#_c_230_n N_VGND_c_590_n 0.00688443f $X=4.695 $Y=0.66 $X2=0
+ $Y2=0
cc_243 N_A_694_21#_c_224_n N_VGND_c_595_n 0.00423334f $X=3.545 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_694_21#_c_225_n N_VGND_c_595_n 0.00541359f $X=3.965 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_694_21#_c_230_n N_VGND_c_598_n 0.0139512f $X=4.695 $Y=0.66 $X2=0
+ $Y2=0
cc_246 N_A_694_21#_c_224_n N_VGND_c_600_n 0.0057435f $X=3.545 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_694_21#_c_225_n N_VGND_c_600_n 0.0108276f $X=3.965 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_694_21#_c_230_n N_VGND_c_600_n 0.0126265f $X=4.695 $Y=0.66 $X2=0
+ $Y2=0
cc_249 N_D_N_M1008_g N_VPWR_c_370_n 0.00482366f $X=4.905 $Y=2.275 $X2=0 $Y2=0
cc_250 D_N N_VPWR_c_370_n 0.00449283f $X=5.205 $Y=1.445 $X2=0 $Y2=0
cc_251 N_D_N_M1008_g N_VPWR_c_372_n 0.00585385f $X=4.905 $Y=2.275 $X2=0 $Y2=0
cc_252 N_D_N_M1008_g N_VPWR_c_368_n 0.0129108f $X=4.905 $Y=2.275 $X2=0 $Y2=0
cc_253 D_N N_VPWR_c_368_n 0.00836565f $X=5.205 $Y=1.445 $X2=0 $Y2=0
cc_254 N_D_N_c_298_n N_VGND_c_589_n 0.00167989f $X=4.967 $Y=0.995 $X2=0 $Y2=0
cc_255 N_D_N_c_295_n N_VGND_c_590_n 0.0102878f $X=5.185 $Y=1.18 $X2=0 $Y2=0
cc_256 N_D_N_c_296_n N_VGND_c_590_n 0.0026033f $X=4.97 $Y=1.16 $X2=0 $Y2=0
cc_257 N_D_N_c_298_n N_VGND_c_590_n 0.00391398f $X=4.967 $Y=0.995 $X2=0 $Y2=0
cc_258 N_D_N_c_299_n N_VGND_c_590_n 0.00375502f $X=5.31 $Y=1.285 $X2=0 $Y2=0
cc_259 N_D_N_c_298_n N_VGND_c_598_n 0.00510437f $X=4.967 $Y=0.995 $X2=0 $Y2=0
cc_260 N_D_N_c_298_n N_VGND_c_600_n 0.00512902f $X=4.967 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_327_n N_VPWR_M1007_s 0.00165831f $X=0.975 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_262 N_A_27_297#_c_327_n N_VPWR_c_369_n 0.0126919f $X=0.975 $Y=1.54 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_c_351_p N_VPWR_c_372_n 0.0142343f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_264 N_A_27_297#_c_326_n N_VPWR_c_374_n 0.0217551f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_265 N_A_27_297#_M1007_d N_VPWR_c_368_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_266 N_A_27_297#_M1013_d N_VPWR_c_368_n 0.00284632f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_267 N_A_27_297#_M1015_s N_VPWR_c_368_n 0.00210147f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_c_326_n N_VPWR_c_368_n 0.0128119f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_269 N_A_27_297#_c_351_p N_VPWR_c_368_n 0.00955092f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_270 N_A_27_297#_c_329_n N_A_277_297#_M1003_d 0.00165831f $X=1.775 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_271 N_A_27_297#_c_329_n N_A_277_297#_c_430_n 0.0126766f $X=1.775 $Y=1.54
+ $X2=0 $Y2=0
cc_272 N_A_27_297#_M1015_s N_A_277_297#_c_426_n 0.00480843f $X=1.805 $Y=1.485
+ $X2=0 $Y2=0
cc_273 N_A_27_297#_c_329_n N_A_277_297#_c_426_n 0.00256303f $X=1.775 $Y=1.54
+ $X2=0 $Y2=0
cc_274 N_A_27_297#_c_330_n N_A_277_297#_c_426_n 0.02056f $X=1.94 $Y=1.63 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_330_n N_A_474_297#_c_445_n 0.0420409f $X=1.94 $Y=1.63 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_329_n N_A_474_297#_c_447_n 0.0159283f $X=1.775 $Y=1.54
+ $X2=0 $Y2=0
cc_277 N_A_27_297#_c_329_n N_Y_c_486_n 0.00297279f $X=1.775 $Y=1.54 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_329_n N_Y_c_490_n 0.0021668f $X=1.775 $Y=1.54 $X2=0 $Y2=0
cc_279 N_A_27_297#_c_328_n N_VGND_c_586_n 5.77871e-19 $X=0.425 $Y=1.54 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_368_n N_A_277_297#_M1003_d 0.0024645f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_281 N_VPWR_c_368_n N_A_277_297#_M1010_s 0.0024645f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_372_n N_A_277_297#_c_426_n 0.0842112f $X=4.99 $Y=2.72 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_368_n N_A_277_297#_c_426_n 0.0521979f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_372_n N_A_277_297#_c_438_n 0.0128741f $X=4.99 $Y=2.72 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_368_n N_A_277_297#_c_438_n 0.00808434f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_368_n N_A_474_297#_M1010_d 0.00210147f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_287 N_VPWR_c_368_n N_A_474_297#_M1014_d 0.00246446f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_368_n N_A_474_297#_M1002_d 0.00226678f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_372_n N_A_474_297#_c_470_n 0.0143053f $X=4.99 $Y=2.72 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_368_n N_A_474_297#_c_470_n 0.00962794f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_372_n N_A_474_297#_c_460_n 0.0485934f $X=4.99 $Y=2.72 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_368_n N_A_474_297#_c_460_n 0.0298944f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_368_n N_Y_M1000_s 0.00216833f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_A_277_297#_c_426_n N_A_474_297#_M1010_d 0.00480843f $X=2.83 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_295 N_A_277_297#_c_426_n N_A_474_297#_c_445_n 0.0249051f $X=2.83 $Y=2.38
+ $X2=0 $Y2=0
cc_296 N_A_277_297#_M1010_s N_A_474_297#_c_446_n 0.00165831f $X=2.78 $Y=1.485
+ $X2=0 $Y2=0
cc_297 N_A_277_297#_c_426_n N_A_474_297#_c_446_n 0.00256303f $X=2.83 $Y=2.38
+ $X2=0 $Y2=0
cc_298 N_A_277_297#_c_444_p N_A_474_297#_c_446_n 0.0126766f $X=2.915 $Y=1.96
+ $X2=0 $Y2=0
cc_299 N_A_474_297#_c_460_n N_Y_M1000_s 0.00312348f $X=4.05 $Y=2.38 $X2=0 $Y2=0
cc_300 N_A_474_297#_c_446_n N_Y_c_488_n 0.00231077f $X=3.21 $Y=1.54 $X2=0 $Y2=0
cc_301 N_A_474_297#_c_447_n N_Y_c_488_n 7.2602e-19 $X=2.66 $Y=1.54 $X2=0 $Y2=0
cc_302 N_A_474_297#_c_446_n N_Y_c_491_n 0.0021668f $X=3.21 $Y=1.54 $X2=0 $Y2=0
cc_303 N_A_474_297#_c_448_n Y 0.0026016f $X=3.335 $Y=1.625 $X2=0 $Y2=0
cc_304 N_A_474_297#_c_460_n Y 0.00341243f $X=4.05 $Y=2.38 $X2=0 $Y2=0
cc_305 N_A_474_297#_c_460_n N_Y_c_554_n 0.0118832f $X=4.05 $Y=2.38 $X2=0 $Y2=0
cc_306 N_Y_c_486_n N_VGND_M1016_d 0.00162089f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_307 N_Y_c_488_n N_VGND_M1012_d 0.00281828f $X=2.75 $Y=0.815 $X2=0 $Y2=0
cc_308 N_Y_c_488_n N_VGND_M1004_d 0.00281828f $X=2.75 $Y=0.815 $X2=0 $Y2=0
cc_309 N_Y_c_489_n N_VGND_M1005_d 0.00162089f $X=3.59 $Y=0.815 $X2=0 $Y2=0
cc_310 N_Y_c_487_n N_VGND_c_586_n 0.00834802f $X=0.845 $Y=0.815 $X2=0 $Y2=0
cc_311 N_Y_c_486_n N_VGND_c_587_n 0.0122559f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_312 N_Y_c_489_n N_VGND_c_588_n 0.0122559f $X=3.59 $Y=0.815 $X2=0 $Y2=0
cc_313 N_Y_c_492_n N_VGND_c_589_n 0.00751095f $X=3.755 $Y=0.815 $X2=0 $Y2=0
cc_314 N_Y_c_496_n N_VGND_c_591_n 0.0188551f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_315 N_Y_c_486_n N_VGND_c_591_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_316 N_Y_c_488_n N_VGND_c_593_n 0.00198695f $X=2.75 $Y=0.815 $X2=0 $Y2=0
cc_317 N_Y_c_516_n N_VGND_c_593_n 0.0188551f $X=2.915 $Y=0.39 $X2=0 $Y2=0
cc_318 N_Y_c_489_n N_VGND_c_593_n 0.00198695f $X=3.59 $Y=0.815 $X2=0 $Y2=0
cc_319 N_Y_c_489_n N_VGND_c_595_n 0.00198695f $X=3.59 $Y=0.815 $X2=0 $Y2=0
cc_320 N_Y_c_520_n N_VGND_c_595_n 0.0188888f $X=3.755 $Y=0.39 $X2=0 $Y2=0
cc_321 N_Y_M1009_s N_VGND_c_600_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_322 N_Y_M1011_s N_VGND_c_600_n 0.00215201f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_323 N_Y_M1004_s N_VGND_c_600_n 0.00215201f $X=2.78 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_M1001_d N_VGND_c_600_n 0.00215201f $X=3.62 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_496_n N_VGND_c_600_n 0.0122069f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_326 N_Y_c_486_n N_VGND_c_600_n 0.00835832f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_327 N_Y_c_504_n N_VGND_c_600_n 0.0122069f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_328 N_Y_c_488_n N_VGND_c_600_n 0.0104597f $X=2.75 $Y=0.815 $X2=0 $Y2=0
cc_329 N_Y_c_516_n N_VGND_c_600_n 0.0122069f $X=2.915 $Y=0.39 $X2=0 $Y2=0
cc_330 N_Y_c_489_n N_VGND_c_600_n 0.00835832f $X=3.59 $Y=0.815 $X2=0 $Y2=0
cc_331 N_Y_c_520_n N_VGND_c_600_n 0.0122162f $X=3.755 $Y=0.39 $X2=0 $Y2=0
cc_332 N_Y_c_486_n N_VGND_c_601_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_333 N_Y_c_504_n N_VGND_c_601_n 0.0188551f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_334 N_Y_c_488_n N_VGND_c_601_n 0.00198695f $X=2.75 $Y=0.815 $X2=0 $Y2=0
cc_335 N_Y_c_488_n N_VGND_c_602_n 0.0564849f $X=2.75 $Y=0.815 $X2=0 $Y2=0

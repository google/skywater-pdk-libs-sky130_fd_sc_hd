* File: sky130_fd_sc_hd__nor4b_4.spice.pex
* Created: Thu Aug 27 14:33:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4B_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r76 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.58 $Y=1.16
+ $X2=1.73 $Y2=1.16
r77 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r78 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.58 $Y2=1.16
r79 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r80 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=0.56 $Y=1.16
+ $X2=0.89 $Y2=1.16
r81 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=1.16 $X2=0.56 $Y2=1.16
r82 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.47 $Y=1.16 $X2=0.56
+ $Y2=1.16
r83 29 40 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=1.135 $Y=1.18
+ $X2=1.58 $Y2=1.18
r84 29 35 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=1.135 $Y=1.18
+ $X2=0.56 $Y2=1.18
r85 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r86 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r87 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r89 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r90 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r91 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r92 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r93 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r94 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r95 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r96 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r97 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r98 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r99 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r79 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.26 $Y=1.16
+ $X2=3.41 $Y2=1.16
r80 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.26
+ $Y=1.16 $X2=3.26 $Y2=1.16
r81 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.26 $Y2=1.16
r82 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r83 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.24 $Y=1.16
+ $X2=2.57 $Y2=1.16
r84 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r85 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.15 $Y=1.16 $X2=2.24
+ $Y2=1.16
r86 29 40 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=2.975 $Y=1.18
+ $X2=3.26 $Y2=1.18
r87 29 35 38.8182 $w=2.08e-07 $l=7.35e-07 $layer=LI1_cond $X=2.975 $Y=1.18
+ $X2=2.24 $Y2=1.18
r88 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r89 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r90 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r92 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r93 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r94 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r95 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r96 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r98 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r100 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r102 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r79 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.46 $Y=1.16
+ $X2=5.61 $Y2=1.16
r80 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.46
+ $Y=1.16 $X2=5.46 $Y2=1.16
r81 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.19 $Y=1.16
+ $X2=5.46 $Y2=1.16
r82 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16
+ $X2=5.19 $Y2=1.16
r83 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.77 $Y2=1.16
r84 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.44
+ $Y=1.16 $X2=4.44 $Y2=1.16
r85 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.35 $Y=1.16 $X2=4.44
+ $Y2=1.16
r86 29 40 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=4.835 $Y=1.18
+ $X2=5.46 $Y2=1.18
r87 29 35 20.8615 $w=2.08e-07 $l=3.95e-07 $layer=LI1_cond $X=4.835 $Y=1.18
+ $X2=4.44 $Y2=1.18
r88 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r89 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r90 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r92 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r93 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r94 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r95 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r96 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r97 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r98 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r99 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r100 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r101 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.985
r102 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r103 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%A_1191_21# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 35 41 43 44 45 46 48 52 61 62 63
c118 61 0 1.47166e-19 $X=7.555 $Y=1.16
r119 68 69 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.87 $Y2=1.16
r120 66 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.45 $Y2=1.16
r121 63 71 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.365 $Y=1.16
+ $X2=7.29 $Y2=1.16
r122 62 63 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=7.555 $Y=1.16
+ $X2=7.365 $Y2=1.16
r123 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.555
+ $Y=1.16 $X2=7.555 $Y2=1.16
r124 52 54 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=8.017 $Y=1.63
+ $X2=8.017 $Y2=2.31
r125 50 52 0.172006 $w=3.33e-07 $l=5e-09 $layer=LI1_cond $X=8.017 $Y=1.625
+ $X2=8.017 $Y2=1.63
r126 46 56 28.8364 $w=1.68e-07 $l=4.42e-07 $layer=LI1_cond $X=7.997 $Y=0.82
+ $X2=7.555 $Y2=0.82
r127 46 48 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=7.997 $Y=0.735
+ $X2=7.997 $Y2=0.39
r128 44 50 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=7.85 $Y=1.54
+ $X2=8.017 $Y2=1.625
r129 44 45 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.85 $Y=1.54
+ $X2=7.64 $Y2=1.54
r130 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=1.455
+ $X2=7.64 $Y2=1.54
r131 42 61 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.555 $Y=1.285
+ $X2=7.555 $Y2=1.18
r132 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.555 $Y=1.285
+ $X2=7.555 $Y2=1.455
r133 41 61 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.555 $Y=1.075
+ $X2=7.555 $Y2=1.18
r134 40 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.905
+ $X2=7.555 $Y2=0.82
r135 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.555 $Y=0.905
+ $X2=7.555 $Y2=1.075
r136 38 71 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.14 $Y=1.16
+ $X2=7.29 $Y2=1.16
r137 38 69 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.14 $Y=1.16
+ $X2=6.87 $Y2=1.16
r138 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.14
+ $Y=1.16 $X2=7.14 $Y2=1.16
r139 35 61 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=1.18
+ $X2=7.555 $Y2=1.18
r140 35 37 17.4286 $w=2.08e-07 $l=3.3e-07 $layer=LI1_cond $X=7.47 $Y=1.18
+ $X2=7.14 $Y2=1.18
r141 31 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.16
r142 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.985
r143 28 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.16
r144 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=0.56
r145 24 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r146 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r147 21 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r148 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r149 17 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r150 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r151 14 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r152 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r153 10 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r154 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r155 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r156 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
r157 2 54 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=7.895
+ $Y=1.485 $X2=8.02 $Y2=2.31
r158 2 52 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.895
+ $Y=1.485 $X2=8.02 $Y2=1.63
r159 1 48 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=7.895
+ $Y=0.235 $X2=8.02 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%D_N 3 6 8 11 13 18
c29 11 0 1.47166e-19 $X=8.395 $Y=1.16
r30 12 18 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=8.395 $Y=1.18
+ $X2=8.51 $Y2=1.18
r31 11 14 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=8.357 $Y=1.16
+ $X2=8.357 $Y2=1.325
r32 11 13 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=8.357 $Y=1.16
+ $X2=8.357 $Y2=0.995
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.395
+ $Y=1.16 $X2=8.395 $Y2=1.16
r34 8 18 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=8.515 $Y=1.18 $X2=8.51
+ $Y2=1.18
r35 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.23 $Y=1.985
+ $X2=8.23 $Y2=1.325
r36 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.23 $Y=0.56 $X2=8.23
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%A_27_297# 1 2 3 4 5 18 22 23 26 28 30 31 32
+ 36 38 42 45 50
r64 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=2.295
+ $X2=3.62 $Y2=1.96
r65 39 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.905 $Y=2.38
+ $X2=2.78 $Y2=2.38
r66 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.495 $Y=2.38
+ $X2=3.62 $Y2=2.295
r67 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.495 $Y=2.38
+ $X2=2.905 $Y2=2.38
r68 34 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.295
+ $X2=2.78 $Y2=2.38
r69 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.78 $Y=2.295
+ $X2=2.78 $Y2=1.96
r70 33 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=2.38
+ $X2=1.94 $Y2=2.38
r71 32 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.78 $Y2=2.38
r72 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.065 $Y2=2.38
r73 31 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=2.38
r74 30 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.625
+ $X2=1.94 $Y2=1.54
r75 30 31 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.94 $Y=1.625
+ $X2=1.94 $Y2=2.295
r76 29 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.54
+ $X2=1.1 $Y2=1.54
r77 28 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=1.54
+ $X2=1.94 $Y2=1.54
r78 28 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.815 $Y=1.54
+ $X2=1.225 $Y2=1.54
r79 24 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.625
+ $X2=1.1 $Y2=1.54
r80 24 26 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.1 $Y=1.625 $X2=1.1
+ $Y2=2.3
r81 22 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=1.1 $Y2=1.54
r82 22 23 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=0.425 $Y2=1.54
r83 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r84 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.425 $Y2=1.54
r85 16 18 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.63
r86 5 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.96
r87 4 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r88 3 49 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2.3
r89 3 47 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.62
r90 2 45 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.62
r91 2 26 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.3
r92 1 20 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r93 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%VPWR 1 2 3 12 16 18 20 24 26 31 36 42 45 49
r104 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r105 45 46 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r106 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 40 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r108 40 46 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 39 40 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r110 37 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.52 $Y2=2.72
r111 37 39 417.866 $w=1.68e-07 $l=6.405e-06 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=8.05 $Y2=2.72
r112 36 48 3.80631 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.547 $Y2=2.72
r113 36 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.05 $Y2=2.72
r114 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r115 35 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 32 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=0.7 $Y2=2.72
r118 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=1.15 $Y2=2.72
r119 31 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.52 $Y2=2.72
r120 31 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.15 $Y2=2.72
r121 26 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.7 $Y2=2.72
r122 26 28 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r123 24 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r125 20 23 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.47 $Y=1.63
+ $X2=8.47 $Y2=2.31
r126 18 48 3.21157 $w=2.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=8.47 $Y=2.635
+ $X2=8.547 $Y2=2.72
r127 18 23 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.47 $Y=2.635
+ $X2=8.47 $Y2=2.31
r128 14 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r129 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=1.96
r130 10 42 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r131 10 12 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=1.96
r132 3 23 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=2.31
r133 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=1.63
r134 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r135 1 12 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%A_445_297# 1 2 3 4 15 19 23 28 30 32 34
r58 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=1.54
+ $X2=4.56 $Y2=1.54
r59 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.275 $Y=1.54
+ $X2=5.4 $Y2=1.54
r60 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.275 $Y=1.54
+ $X2=4.685 $Y2=1.54
r61 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=1.54
+ $X2=3.2 $Y2=1.54
r62 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=1.54
+ $X2=4.56 $Y2=1.54
r63 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.435 $Y=1.54
+ $X2=3.325 $Y2=1.54
r64 16 28 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.485 $Y=1.54
+ $X2=2.36 $Y2=1.54
r65 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=1.54
+ $X2=3.2 $Y2=1.54
r66 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.075 $Y=1.54
+ $X2=2.485 $Y2=1.54
r67 4 34 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.62
r68 3 32 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.62
r69 2 30 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.62
r70 1 28 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%A_803_297# 1 2 3 4 5 18 20 21 24 26 30 32 36
+ 38 42 44 46 47
r65 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.5 $Y=2.295
+ $X2=7.5 $Y2=1.96
r66 39 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.38
+ $X2=6.66 $Y2=2.38
r67 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.375 $Y=2.38
+ $X2=7.5 $Y2=2.295
r68 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.375 $Y=2.38
+ $X2=6.785 $Y2=2.38
r69 34 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.295
+ $X2=6.66 $Y2=2.38
r70 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.66 $Y=2.295
+ $X2=6.66 $Y2=1.96
r71 33 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=2.38
+ $X2=5.82 $Y2=2.38
r72 32 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=2.38
+ $X2=6.66 $Y2=2.38
r73 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.535 $Y=2.38
+ $X2=5.945 $Y2=2.38
r74 28 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.295
+ $X2=5.82 $Y2=2.38
r75 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.82 $Y=2.295
+ $X2=5.82 $Y2=1.62
r76 27 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.38
+ $X2=4.98 $Y2=2.38
r77 26 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=2.38
+ $X2=5.82 $Y2=2.38
r78 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.695 $Y=2.38
+ $X2=5.105 $Y2=2.38
r79 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=2.38
r80 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.98 $Y=2.295
+ $X2=4.98 $Y2=1.96
r81 20 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.98 $Y2=2.38
r82 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.855 $Y=2.38
+ $X2=4.265 $Y2=2.38
r83 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.14 $Y=2.295
+ $X2=4.265 $Y2=2.38
r84 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=2.295
+ $X2=4.14 $Y2=1.96
r85 5 42 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=1.96
r86 4 36 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.96
r87 3 46 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.3
r88 3 30 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=1.62
r89 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=1.96
r90 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.485 $X2=4.14 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45 47
+ 51 53 57 59 63 65 69 72 73 75 79 83 84 85 86 87 88 91 93 94
c201 91 0 1.70807e-19 $X=6.24 $Y=1.62
r202 89 94 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.24 $Y=1.625
+ $X2=6.24 $Y2=1.87
r203 89 91 3.14896 $w=3e-07 $l=1.07121e-07 $layer=LI1_cond $X=6.24 $Y=1.625
+ $X2=6.29 $Y2=1.54
r204 77 79 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.08 $Y=0.725
+ $X2=7.08 $Y2=0.39
r205 76 91 3.44808 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.465 $Y=1.54
+ $X2=6.29 $Y2=1.54
r206 75 93 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=1.54
+ $X2=7.08 $Y2=1.54
r207 75 76 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.955 $Y=1.54
+ $X2=6.465 $Y2=1.54
r208 74 88 5.1752 $w=1.8e-07 $l=1.95e-07 $layer=LI1_cond $X=6.465 $Y=0.815
+ $X2=6.27 $Y2=0.815
r209 73 77 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.915 $Y=0.815
+ $X2=7.08 $Y2=0.725
r210 73 74 27.7273 $w=1.78e-07 $l=4.5e-07 $layer=LI1_cond $X=6.915 $Y=0.815
+ $X2=6.465 $Y2=0.815
r211 72 91 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.29 $Y=1.455 $X2=6.29
+ $Y2=1.54
r212 71 88 1.36226 $w=3.5e-07 $l=9.94987e-08 $layer=LI1_cond $X=6.29 $Y=0.905
+ $X2=6.27 $Y2=0.815
r213 71 72 18.1098 $w=3.48e-07 $l=5.5e-07 $layer=LI1_cond $X=6.29 $Y=0.905
+ $X2=6.29 $Y2=1.455
r214 67 88 1.36226 $w=3.3e-07 $l=1.03923e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.27 $Y2=0.815
r215 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.39
r216 66 87 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0.815
+ $X2=5.4 $Y2=0.815
r217 65 88 5.1752 $w=1.8e-07 $l=1.95e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=6.27 $Y2=0.815
r218 65 66 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=5.565 $Y2=0.815
r219 61 87 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.4 $Y=0.725 $X2=5.4
+ $Y2=0.815
r220 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.4 $Y=0.725
+ $X2=5.4 $Y2=0.39
r221 60 86 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=0.815
+ $X2=4.56 $Y2=0.815
r222 59 87 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=5.4 $Y2=0.815
r223 59 60 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.235 $Y=0.815
+ $X2=4.725 $Y2=0.815
r224 55 86 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.56 $Y=0.725
+ $X2=4.56 $Y2=0.815
r225 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.725
+ $X2=4.56 $Y2=0.39
r226 54 85 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=0.815
+ $X2=3.2 $Y2=0.815
r227 53 86 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=4.56 $Y2=0.815
r228 53 54 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=3.365 $Y2=0.815
r229 49 85 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.2 $Y=0.725 $X2=3.2
+ $Y2=0.815
r230 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.2 $Y=0.725
+ $X2=3.2 $Y2=0.39
r231 48 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0.815
+ $X2=2.36 $Y2=0.815
r232 47 85 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=3.2 $Y2=0.815
r233 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.035 $Y=0.815
+ $X2=2.525 $Y2=0.815
r234 43 84 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.36 $Y=0.725
+ $X2=2.36 $Y2=0.815
r235 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.36 $Y=0.725
+ $X2=2.36 $Y2=0.39
r236 42 83 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=0.815
+ $X2=1.52 $Y2=0.815
r237 41 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0.815
+ $X2=2.36 $Y2=0.815
r238 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.195 $Y=0.815
+ $X2=1.685 $Y2=0.815
r239 37 83 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.52 $Y=0.725
+ $X2=1.52 $Y2=0.815
r240 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=0.725
+ $X2=1.52 $Y2=0.39
r241 35 83 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=1.52 $Y2=0.815
r242 35 36 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=0.845 $Y2=0.815
r243 31 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.845 $Y2=0.815
r244 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.68 $Y2=0.39
r245 10 93 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=1.62
r246 9 91 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.62
r247 8 79 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.39
r248 7 69 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
r249 6 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.39
r250 5 57 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.39
r251 4 51 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.39
r252 3 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.39
r253 2 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r254 1 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4B_4%VGND 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 51 55 59 63 65 67 70 71 73 74 76 77 78 79 81 82 84 85 86 113 123 126 128 132
r157 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r158 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r159 125 126 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.235
+ $X2=4.225 $Y2=0.235
r160 121 125 4.29841 $w=6.38e-07 $l=2.3e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=4.14 $Y2=0.235
r161 121 123 14.3415 $w=6.38e-07 $l=3.75e-07 $layer=LI1_cond $X=3.91 $Y=0.235
+ $X2=3.535 $Y2=0.235
r162 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r163 116 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r164 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r165 113 131 3.80631 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=8.355 $Y=0
+ $X2=8.547 $Y2=0
r166 113 115 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=0
+ $X2=8.05 $Y2=0
r167 112 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r168 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r169 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r170 109 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r171 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r172 106 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.82 $Y2=0
r173 106 108 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r174 105 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r175 105 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=3.91 $Y2=0
r176 104 126 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.225 $Y2=0
r177 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r178 101 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r179 100 123 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=3.535 $Y2=0
r180 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r181 97 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r182 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r183 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r184 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r185 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r186 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r187 88 118 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r188 88 90 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r189 86 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r190 86 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r191 84 111 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.415 $Y=0
+ $X2=7.13 $Y2=0
r192 84 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=0 $X2=7.5
+ $Y2=0
r193 83 115 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.585 $Y=0
+ $X2=8.05 $Y2=0
r194 83 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.5
+ $Y2=0
r195 81 108 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r196 81 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0 $X2=6.66
+ $Y2=0
r197 80 111 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.13 $Y2=0
r198 80 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.66
+ $Y2=0
r199 78 104 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.83 $Y2=0
r200 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r201 76 96 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=2.53 $Y2=0
r202 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.78
+ $Y2=0
r203 75 100 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=3.45 $Y2=0
r204 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.78
+ $Y2=0
r205 73 93 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r206 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r207 72 96 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.53 $Y2=0
r208 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r209 70 90 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r210 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r211 69 93 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=1.61 $Y2=0
r212 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r213 65 131 3.21157 $w=2.3e-07 $l=1.17346e-07 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.547 $Y2=0
r214 65 67 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.47 $Y2=0.39
r215 61 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r216 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.39
r217 57 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0
r218 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0.39
r219 53 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r220 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.39
r221 52 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r222 51 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r223 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r224 47 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r225 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r226 43 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r227 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.39
r228 39 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r229 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.39
r230 35 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r231 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.39
r232 31 118 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r233 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r234 10 67 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.39
r235 9 63 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.39
r236 8 59 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r237 7 55 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.39
r238 6 49 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r239 5 125 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.235 $X2=4.14 $Y2=0.39
r240 4 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.39
r241 3 41 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r242 2 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r243 1 33 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends


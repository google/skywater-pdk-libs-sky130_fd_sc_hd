# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.570000 1.700000 ;
    END
  END A
  PIN X
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.660000 0.255000 3.105000 0.825000 ;
        RECT 2.660000 1.495000 3.565000 1.675000 ;
        RECT 2.660000 1.675000 3.105000 2.465000 ;
        RECT 2.735000 0.825000 3.105000 0.995000 ;
        RECT 2.735000 0.995000 3.565000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.690000  0.085000 1.075000 0.485000 ;
        RECT 2.105000  0.085000 2.490000 0.485000 ;
        RECT 3.700000  0.085000 4.085000 0.485000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.690000 2.210000 1.075000 2.635000 ;
        RECT 2.105000 2.210000 2.490000 2.635000 ;
        RECT 3.700000 2.210000 4.085000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.520000 0.655000 ;
      RECT 0.085000 0.655000 1.075000 0.825000 ;
      RECT 0.085000 1.870000 1.075000 2.040000 ;
      RECT 0.085000 2.040000 0.520000 2.465000 ;
      RECT 0.740000 0.825000 1.075000 0.995000 ;
      RECT 0.740000 0.995000 1.150000 1.325000 ;
      RECT 0.740000 1.325000 1.075000 1.870000 ;
      RECT 1.245000 0.255000 1.515000 0.825000 ;
      RECT 1.245000 1.495000 1.970000 1.675000 ;
      RECT 1.245000 1.675000 1.515000 2.465000 ;
      RECT 1.320000 0.825000 1.515000 0.995000 ;
      RECT 1.320000 0.995000 1.970000 1.495000 ;
      RECT 1.685000 0.255000 1.935000 0.655000 ;
      RECT 1.685000 0.655000 2.490000 0.825000 ;
      RECT 1.685000 1.845000 2.490000 2.040000 ;
      RECT 1.685000 2.040000 1.935000 2.465000 ;
      RECT 2.140000 0.825000 2.490000 0.995000 ;
      RECT 2.140000 0.995000 2.565000 1.325000 ;
      RECT 2.140000 1.325000 2.490000 1.845000 ;
      RECT 3.275000 0.255000 3.530000 0.655000 ;
      RECT 3.275000 0.655000 4.085000 0.825000 ;
      RECT 3.275000 1.845000 4.085000 2.040000 ;
      RECT 3.275000 2.040000 3.530000 2.465000 ;
      RECT 3.735000 0.825000 4.085000 0.995000 ;
      RECT 3.735000 0.995000 4.160000 1.325000 ;
      RECT 3.735000 1.325000 4.085000 1.845000 ;
      RECT 4.255000 0.255000 4.515000 0.825000 ;
      RECT 4.255000 1.495000 4.515000 2.465000 ;
      RECT 4.330000 0.825000 4.515000 1.495000 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1

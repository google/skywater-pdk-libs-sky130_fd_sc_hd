* File: sky130_fd_sc_hd__lpflow_inputisolatch_1.pxi.spice
* Created: Tue Sep  1 19:12:27 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%SLEEP_B N_SLEEP_B_c_116_n
+ N_SLEEP_B_c_111_n N_SLEEP_B_M1015_g N_SLEEP_B_c_117_n N_SLEEP_B_M1012_g
+ N_SLEEP_B_c_112_n N_SLEEP_B_c_118_n SLEEP_B N_SLEEP_B_c_113_n
+ N_SLEEP_B_c_114_n SLEEP_B PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%SLEEP_B
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_27_47# N_A_27_47#_M1015_s
+ N_A_27_47#_M1012_s N_A_27_47#_M1010_g N_A_27_47#_M1002_g N_A_27_47#_M1009_g
+ N_A_27_47#_c_152_n N_A_27_47#_c_153_n N_A_27_47#_M1001_g N_A_27_47#_c_166_n
+ N_A_27_47#_c_280_p N_A_27_47#_c_167_n N_A_27_47#_c_155_n N_A_27_47#_c_156_n
+ N_A_27_47#_c_168_n N_A_27_47#_c_169_n N_A_27_47#_c_170_n N_A_27_47#_c_157_n
+ N_A_27_47#_c_158_n N_A_27_47#_c_172_n N_A_27_47#_c_159_n N_A_27_47#_c_160_n
+ N_A_27_47#_c_174_n N_A_27_47#_c_175_n N_A_27_47#_c_176_n N_A_27_47#_c_161_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_27_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%D N_D_M1004_g N_D_M1013_g D
+ N_D_c_290_n N_D_c_291_n D PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%D
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_193_47# N_A_193_47#_M1010_d
+ N_A_193_47#_M1002_d N_A_193_47#_M1014_g N_A_193_47#_M1003_g
+ N_A_193_47#_c_332_n N_A_193_47#_c_333_n N_A_193_47#_c_341_n
+ N_A_193_47#_c_342_n N_A_193_47#_c_334_n N_A_193_47#_c_335_n
+ N_A_193_47#_c_336_n N_A_193_47#_c_343_n N_A_193_47#_c_344_n
+ N_A_193_47#_c_337_n N_A_193_47#_c_338_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_193_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_629_21# N_A_629_21#_M1008_s
+ N_A_629_21#_M1007_s N_A_629_21#_M1005_g N_A_629_21#_M1011_g
+ N_A_629_21#_c_455_n N_A_629_21#_c_456_n N_A_629_21#_c_452_n
+ N_A_629_21#_c_465_p N_A_629_21#_c_468_p
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_629_21#
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_476_47# N_A_476_47#_M1014_d
+ N_A_476_47#_M1009_d N_A_476_47#_c_509_n N_A_476_47#_M1008_g
+ N_A_476_47#_M1007_g N_A_476_47#_c_510_n N_A_476_47#_M1006_g
+ N_A_476_47#_M1000_g N_A_476_47#_c_511_n N_A_476_47#_c_512_n
+ N_A_476_47#_c_522_n N_A_476_47#_c_523_n N_A_476_47#_c_513_n
+ N_A_476_47#_c_514_n N_A_476_47#_c_520_n N_A_476_47#_c_515_n
+ PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%A_476_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VPWR N_VPWR_M1012_d N_VPWR_M1013_s
+ N_VPWR_M1011_d N_VPWR_M1007_d N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n
+ N_VPWR_c_613_n VPWR N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n
+ N_VPWR_c_617_n N_VPWR_c_609_n N_VPWR_c_619_n N_VPWR_c_620_n N_VPWR_c_621_n
+ N_VPWR_c_622_n PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%Q N_Q_M1006_d N_Q_M1000_d Q Q Q Q
+ N_Q_c_691_n PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%Q
x_PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VGND N_VGND_M1015_d N_VGND_M1004_s
+ N_VGND_M1005_d N_VGND_M1008_d N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ N_VGND_c_705_n N_VGND_c_706_n VGND N_VGND_c_707_n N_VGND_c_708_n
+ N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n
+ N_VGND_c_714_n N_VGND_c_715_n PM_SKY130_FD_SC_HD__LPFLOW_INPUTISOLATCH_1%VGND
cc_1 VNB N_SLEEP_B_c_111_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_SLEEP_B_c_112_n 0.0269894f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB N_SLEEP_B_c_113_n 0.0212418f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_4 VNB N_SLEEP_B_c_114_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.07
cc_5 VNB SLEEP_B 0.0153903f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.275
cc_6 VNB N_A_27_47#_M1010_g 0.0406707f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.18
cc_7 VNB N_A_27_47#_c_152_n 0.0132134f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.22
cc_8 VNB N_A_27_47#_c_153_n 0.00482312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1001_g 0.0422907f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_10 VNB N_A_27_47#_c_155_n 0.00300884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_156_n 0.00637392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_157_n 0.00668532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_158_n 0.0251933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_159_n 4.92268e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_160_n 0.00502604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_161_n 0.0190638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_D_M1013_g 0.0145876f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_290_n 0.0345228f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_19 VNB N_D_c_291_n 0.0176004f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_20 VNB D 0.00677853f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_193_47#_c_332_n 0.00725367f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.75
cc_22 VNB N_A_193_47#_c_333_n 0.00219325f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_193_47#_c_334_n 0.00523587f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.275
cc_24 VNB N_A_193_47#_c_335_n 0.0275313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_193_47#_c_336_n 0.00368432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_193_47#_c_337_n 0.00449519f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_338_n 0.0176559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_629_21#_M1005_g 0.0514221f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.18
cc_29 VNB N_A_629_21#_c_452_n 0.00161624f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_30 VNB N_A_476_47#_c_509_n 0.0199362f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_31 VNB N_A_476_47#_c_510_n 0.0192326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_476_47#_c_511_n 0.0437903f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_33 VNB N_A_476_47#_c_512_n 0.0290757f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_34 VNB N_A_476_47#_c_513_n 0.00368943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_476_47#_c_514_n 0.00973996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_476_47#_c_515_n 0.00318788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_609_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB Q 0.0131477f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.18
cc_39 VNB N_Q_c_691_n 0.0263331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_702_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.75
cc_41 VNB N_VGND_c_703_n 0.00623966f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.22
cc_42 VNB N_VGND_c_704_n 0.00708664f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_43 VNB N_VGND_c_705_n 0.0202314f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.4
cc_44 VNB N_VGND_c_706_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.277
cc_45 VNB N_VGND_c_707_n 0.0153958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_708_n 0.0168401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_709_n 0.0396117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_710_n 0.0191314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_711_n 0.277704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_712_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_713_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_714_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_715_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VPB N_SLEEP_B_c_116_n 0.0191615f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.675
cc_55 VPB N_SLEEP_B_c_117_n 0.0175976f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.825
cc_56 VPB N_SLEEP_B_c_118_n 0.028256f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.75
cc_57 VPB N_SLEEP_B_c_113_n 0.0104393f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_58 VPB SLEEP_B 0.0153801f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.275
cc_59 VPB N_A_27_47#_M1002_g 0.0313098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_60 VPB N_A_27_47#_M1009_g 0.0297117f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.75
cc_61 VPB N_A_27_47#_c_152_n 0.0165043f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.22
cc_62 VPB N_A_27_47#_c_153_n 0.00915765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_166_n 0.0112459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_167_n 0.00167773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_168_n 0.00265225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_169_n 0.00479024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_170_n 0.00511037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_158_n 0.0374771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_172_n 0.00249827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_159_n 4.9608e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_174_n 0.00390582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_175_n 0.00947367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_176_n 0.0119477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_161_n 0.0200724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_D_M1013_g 0.0416231f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_76 VPB N_A_193_47#_M1003_g 0.0194322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_193_47#_c_332_n 0.00453726f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.75
cc_78 VPB N_A_193_47#_c_341_n 0.00402821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_193_47#_c_342_n 0.00965908f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_80 VPB N_A_193_47#_c_343_n 0.00654274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_193_47#_c_344_n 0.0263514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_193_47#_c_337_n 0.00266526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_629_21#_M1005_g 0.0162878f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.18
cc_84 VPB N_A_629_21#_M1011_g 0.0257045f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_85 VPB N_A_629_21#_c_455_n 0.00536583f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.75
cc_86 VPB N_A_629_21#_c_456_n 0.0471252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_629_21#_c_452_n 0.00235089f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_88 VPB N_A_476_47#_M1007_g 0.0230156f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_476_47#_M1000_g 0.0219746f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.22
cc_90 VPB N_A_476_47#_c_511_n 0.0151805f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_91 VPB N_A_476_47#_c_512_n 0.00400545f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_92 VPB N_A_476_47#_c_520_n 0.00524045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_476_47#_c_515_n 0.00200173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_610_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.75
cc_95 VPB N_VPWR_c_611_n 0.00470153f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.22
cc_96 VPB N_VPWR_c_612_n 0.0218842f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_97 VPB N_VPWR_c_613_n 0.00467718f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.4
cc_98 VPB N_VPWR_c_614_n 0.0154981f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.277
cc_99 VPB N_VPWR_c_615_n 0.015602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_616_n 0.0371591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_617_n 0.0184665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_609_n 0.0581437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_619_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_620_n 0.0108022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_621_n 0.00324376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_622_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB Q 0.00545527f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.18
cc_108 VPB Q 0.0250272f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.22
cc_109 VPB N_Q_c_691_n 0.0159642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 N_SLEEP_B_c_111_n N_A_27_47#_M1010_g 0.018783f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_111 N_SLEEP_B_c_114_n N_A_27_47#_M1010_g 0.00469172f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_112 N_SLEEP_B_c_118_n N_A_27_47#_M1002_g 0.0224183f $X=0.47 $Y=1.75 $X2=0
+ $Y2=0
cc_113 N_SLEEP_B_c_117_n N_A_27_47#_c_167_n 0.00214396f $X=0.47 $Y=1.825 $X2=0
+ $Y2=0
cc_114 N_SLEEP_B_c_111_n N_A_27_47#_c_155_n 0.00663556f $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_115 N_SLEEP_B_c_112_n N_A_27_47#_c_155_n 0.0105293f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_116 N_SLEEP_B_c_112_n N_A_27_47#_c_156_n 0.00657185f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_117 N_SLEEP_B_c_113_n N_A_27_47#_c_156_n 3.35813e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_118 SLEEP_B N_A_27_47#_c_156_n 0.0125186f $X=0.21 $Y=1.275 $X2=0 $Y2=0
cc_119 N_SLEEP_B_c_117_n N_A_27_47#_c_168_n 0.00928899f $X=0.47 $Y=1.825 $X2=0
+ $Y2=0
cc_120 N_SLEEP_B_c_118_n N_A_27_47#_c_168_n 0.00942493f $X=0.47 $Y=1.75 $X2=0
+ $Y2=0
cc_121 N_SLEEP_B_c_118_n N_A_27_47#_c_169_n 0.0056661f $X=0.47 $Y=1.75 $X2=0
+ $Y2=0
cc_122 N_SLEEP_B_c_113_n N_A_27_47#_c_169_n 2.59784e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_123 SLEEP_B N_A_27_47#_c_169_n 0.0134567f $X=0.21 $Y=1.275 $X2=0 $Y2=0
cc_124 N_SLEEP_B_c_116_n N_A_27_47#_c_170_n 0.00225292f $X=0.305 $Y=1.675 $X2=0
+ $Y2=0
cc_125 N_SLEEP_B_c_118_n N_A_27_47#_c_170_n 0.00288097f $X=0.47 $Y=1.75 $X2=0
+ $Y2=0
cc_126 N_SLEEP_B_c_113_n N_A_27_47#_c_159_n 0.00109738f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_127 N_SLEEP_B_c_112_n N_A_27_47#_c_160_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_128 N_SLEEP_B_c_114_n N_A_27_47#_c_160_n 0.00327197f $X=0.245 $Y=1.07 $X2=0
+ $Y2=0
cc_129 SLEEP_B N_A_27_47#_c_160_n 0.0311882f $X=0.21 $Y=1.275 $X2=0 $Y2=0
cc_130 N_SLEEP_B_c_116_n N_A_27_47#_c_161_n 0.00428171f $X=0.305 $Y=1.675 $X2=0
+ $Y2=0
cc_131 N_SLEEP_B_c_113_n N_A_27_47#_c_161_n 0.02077f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_132 SLEEP_B N_A_27_47#_c_161_n 0.00119742f $X=0.21 $Y=1.275 $X2=0 $Y2=0
cc_133 N_SLEEP_B_c_117_n N_VPWR_c_610_n 0.00946555f $X=0.47 $Y=1.825 $X2=0 $Y2=0
cc_134 N_SLEEP_B_c_117_n N_VPWR_c_614_n 0.00332278f $X=0.47 $Y=1.825 $X2=0 $Y2=0
cc_135 N_SLEEP_B_c_117_n N_VPWR_c_609_n 0.00484884f $X=0.47 $Y=1.825 $X2=0 $Y2=0
cc_136 N_SLEEP_B_c_111_n N_VGND_c_702_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_137 N_SLEEP_B_c_111_n N_VGND_c_707_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_138 N_SLEEP_B_c_112_n N_VGND_c_707_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_139 N_SLEEP_B_c_111_n N_VGND_c_711_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1009_g N_D_M1013_g 0.0365817f $X=2.305 $Y=2.275 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_153_n N_D_M1013_g 0.025257f $X=2.385 $Y=1.32 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_157_n N_D_M1013_g 0.00151855f $X=1.405 $Y=1.415 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_158_n N_D_M1013_g 0.0214184f $X=1.405 $Y=1.415 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_174_n N_D_M1013_g 0.0016959f $X=2.25 $Y=1.52 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_176_n N_D_M1013_g 0.0126765f $X=2.05 $Y=1.525 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_176_n N_D_c_290_n 0.0027653f $X=2.05 $Y=1.525 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_153_n D 2.15306e-19 $X=2.385 $Y=1.32 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_174_n D 0.00461433f $X=2.25 $Y=1.52 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_176_n D 0.0110081f $X=2.05 $Y=1.525 $X2=0 $Y2=0
cc_150 N_A_27_47#_M1009_g N_A_193_47#_M1003_g 0.0194476f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1002_g N_A_193_47#_c_332_n 0.00574027f $X=0.89 $Y=2.18 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_168_n N_A_193_47#_c_332_n 0.00220137f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_170_n N_A_193_47#_c_332_n 0.0219593f $X=0.695 $Y=1.795 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_157_n N_A_193_47#_c_332_n 0.0193587f $X=1.405 $Y=1.415 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_158_n N_A_193_47#_c_332_n 0.0216332f $X=1.405 $Y=1.415 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_172_n N_A_193_47#_c_332_n 0.0139021f $X=1.49 $Y=1.61 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_159_n N_A_193_47#_c_332_n 0.0230986f $X=0.725 $Y=1.295 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_161_n N_A_193_47#_c_332_n 0.00625081f $X=0.965 $Y=1.415
+ $X2=0 $Y2=0
cc_159 N_A_27_47#_M1010_g N_A_193_47#_c_333_n 0.00194826f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_155_n N_A_193_47#_c_333_n 0.00555973f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_M1002_g N_A_193_47#_c_341_n 0.00494892f $X=0.89 $Y=2.18 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_168_n N_A_193_47#_c_341_n 0.00598752f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_158_n N_A_193_47#_c_341_n 0.00141497f $X=1.405 $Y=1.415
+ $X2=0 $Y2=0
cc_164 N_A_27_47#_M1009_g N_A_193_47#_c_342_n 0.0120393f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_152_n N_A_193_47#_c_342_n 0.00283672f $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_166_n N_A_193_47#_c_342_n 9.32506e-19 $X=2.25 $Y=1.685 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_158_n N_A_193_47#_c_342_n 0.00538861f $X=1.405 $Y=1.415
+ $X2=0 $Y2=0
cc_168 N_A_27_47#_c_172_n N_A_193_47#_c_342_n 0.0115921f $X=1.49 $Y=1.61 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_176_n N_A_193_47#_c_342_n 0.0479011f $X=2.05 $Y=1.525 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1010_g N_A_193_47#_c_334_n 0.00625081f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_155_n N_A_193_47#_c_334_n 0.00490576f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_158_n N_A_193_47#_c_334_n 0.0012239f $X=1.405 $Y=1.415 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_160_n N_A_193_47#_c_334_n 0.0218122f $X=0.71 $Y=1.13 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_153_n N_A_193_47#_c_335_n 0.0197851f $X=2.385 $Y=1.32 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_M1001_g N_A_193_47#_c_335_n 0.0192833f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_174_n N_A_193_47#_c_335_n 5.32821e-19 $X=2.25 $Y=1.52 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_152_n N_A_193_47#_c_336_n 7.03475e-19 $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_153_n N_A_193_47#_c_336_n 0.00136018f $X=2.385 $Y=1.32 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1001_g N_A_193_47#_c_336_n 0.00233362f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_174_n N_A_193_47#_c_336_n 0.0018132f $X=2.25 $Y=1.52 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1009_g N_A_193_47#_c_343_n 0.00565485f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_182 N_A_27_47#_c_152_n N_A_193_47#_c_343_n 0.00429262f $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_166_n N_A_193_47#_c_343_n 0.00262328f $X=2.25 $Y=1.685 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_M1009_g N_A_193_47#_c_344_n 0.0108146f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_152_n N_A_193_47#_c_344_n 0.0184291f $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_166_n N_A_193_47#_c_344_n 0.00489663f $X=2.25 $Y=1.685 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_152_n N_A_193_47#_c_337_n 0.0127914f $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1001_g N_A_193_47#_c_337_n 0.0048515f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_174_n N_A_193_47#_c_337_n 0.0263212f $X=2.25 $Y=1.52 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_175_n N_A_193_47#_c_337_n 0.00262328f $X=2.25 $Y=1.52 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1001_g N_A_193_47#_c_338_n 0.0162516f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1001_g N_A_629_21#_M1005_g 0.0579998f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_M1009_g N_A_476_47#_c_522_n 0.00493481f $X=2.305 $Y=2.275
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_M1001_g N_A_476_47#_c_523_n 0.0119295f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1001_g N_A_476_47#_c_513_n 0.00889873f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_M1001_g N_A_476_47#_c_514_n 0.00530536f $X=2.8 $Y=0.415 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_152_n N_A_476_47#_c_520_n 6.38593e-19 $X=2.725 $Y=1.32 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_168_n N_VPWR_M1012_d 0.00176788f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_199 N_A_27_47#_M1002_g N_VPWR_c_610_n 0.0094125f $X=0.89 $Y=2.18 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_167_n N_VPWR_c_610_n 0.012721f $X=0.26 $Y=2.175 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_168_n N_VPWR_c_610_n 0.0155904f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_161_n N_VPWR_c_610_n 4.89682e-19 $X=0.965 $Y=1.415 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_167_n N_VPWR_c_614_n 0.0120313f $X=0.26 $Y=2.175 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_168_n N_VPWR_c_614_n 0.00185988f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_205 N_A_27_47#_M1002_g N_VPWR_c_615_n 0.00442511f $X=0.89 $Y=2.18 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1009_g N_VPWR_c_616_n 0.00397569f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_M1002_g N_VPWR_c_609_n 0.00889084f $X=0.89 $Y=2.18 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1009_g N_VPWR_c_609_n 0.00574885f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_167_n N_VPWR_c_609_n 0.00646745f $X=0.26 $Y=2.175 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_168_n N_VPWR_c_609_n 0.00484649f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_211 N_A_27_47#_M1002_g N_VPWR_c_620_n 0.00180726f $X=0.89 $Y=2.18 $X2=0 $Y2=0
cc_212 N_A_27_47#_M1009_g N_VPWR_c_620_n 0.00200519f $X=2.305 $Y=2.275 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_155_n N_VGND_M1015_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_27_47#_M1010_g N_VGND_c_702_n 0.00895942f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_155_n N_VGND_c_702_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_161_n N_VGND_c_702_n 4.88844e-19 $X=0.965 $Y=1.415 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_M1010_g N_VGND_c_703_n 0.00301453f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1001_g N_VGND_c_704_n 0.00182134f $X=2.8 $Y=0.415 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_280_p N_VGND_c_707_n 0.00713694f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_155_n N_VGND_c_707_n 0.00243651f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1010_g N_VGND_c_708_n 0.0046653f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_27_47#_M1001_g N_VGND_c_709_n 0.00379804f $X=2.8 $Y=0.415 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1015_s N_VGND_c_711_n 0.003754f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1010_g N_VGND_c_711_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1001_g N_VGND_c_711_n 0.00557952f $X=2.8 $Y=0.415 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_280_p N_VGND_c_711_n 0.00608739f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_155_n N_VGND_c_711_n 0.00549708f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_228 N_D_M1013_g N_A_193_47#_c_332_n 0.0064022f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_229 N_D_c_290_n N_A_193_47#_c_332_n 0.00303853f $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_230 D N_A_193_47#_c_332_n 0.00535366f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_231 N_D_c_290_n N_A_193_47#_c_333_n 0.00337468f $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_232 N_D_c_291_n N_A_193_47#_c_333_n 0.00474548f $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_233 N_D_M1013_g N_A_193_47#_c_341_n 0.0046822f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_234 N_D_M1013_g N_A_193_47#_c_342_n 0.0135107f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_235 D N_A_193_47#_c_334_n 0.00448013f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_236 N_D_c_290_n N_A_193_47#_c_335_n 0.0144205f $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_237 D N_A_193_47#_c_335_n 0.00193086f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_238 N_D_c_290_n N_A_193_47#_c_336_n 4.46416e-19 $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_239 D N_A_193_47#_c_336_n 0.0218559f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_240 N_D_M1013_g N_A_193_47#_c_337_n 0.00370009f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_241 N_D_c_290_n N_A_193_47#_c_337_n 2.6569e-19 $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_242 D N_A_193_47#_c_337_n 0.00271645f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_243 N_D_c_291_n N_A_193_47#_c_338_n 0.025355f $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_244 N_D_M1013_g N_A_476_47#_c_522_n 5.30748e-19 $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_245 N_D_c_291_n N_A_476_47#_c_523_n 6.01098e-19 $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_246 N_D_M1013_g N_VPWR_c_616_n 0.00155868f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_247 N_D_M1013_g N_VPWR_c_609_n 0.00240573f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_248 N_D_M1013_g N_VPWR_c_620_n 0.0141656f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_249 N_D_c_291_n N_VGND_c_703_n 0.010947f $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_250 D N_VGND_c_703_n 0.00136609f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_251 N_D_c_290_n N_VGND_c_709_n 0.00120761f $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_252 N_D_c_291_n N_VGND_c_709_n 0.0046653f $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_253 N_D_c_290_n N_VGND_c_711_n 0.00158512f $X=1.835 $Y=0.93 $X2=0 $Y2=0
cc_254 N_D_c_291_n N_VGND_c_711_n 0.00440885f $X=1.835 $Y=0.73 $X2=0 $Y2=0
cc_255 D N_VGND_c_711_n 0.0122902f $X=1.92 $Y=0.925 $X2=0 $Y2=0
cc_256 N_A_193_47#_c_337_n N_A_629_21#_M1005_g 9.87052e-19 $X=2.675 $Y=1.575
+ $X2=0 $Y2=0
cc_257 N_A_193_47#_M1003_g N_A_629_21#_M1011_g 0.0256604f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_258 N_A_193_47#_c_343_n N_A_629_21#_M1011_g 5.33856e-19 $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_259 N_A_193_47#_c_343_n N_A_629_21#_c_456_n 3.93081e-19 $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_260 N_A_193_47#_c_344_n N_A_629_21#_c_456_n 0.0157438f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_261 N_A_193_47#_c_342_n N_A_476_47#_M1009_d 7.42631e-19 $X=2.505 $Y=2 $X2=0
+ $Y2=0
cc_262 N_A_193_47#_c_343_n N_A_476_47#_M1009_d 9.73695e-19 $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_263 N_A_193_47#_M1003_g N_A_476_47#_c_522_n 0.00825554f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_264 N_A_193_47#_c_342_n N_A_476_47#_c_522_n 0.00915594f $X=2.505 $Y=2 $X2=0
+ $Y2=0
cc_265 N_A_193_47#_c_343_n N_A_476_47#_c_522_n 0.0172353f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_266 N_A_193_47#_c_344_n N_A_476_47#_c_522_n 0.00219621f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_267 N_A_193_47#_c_335_n N_A_476_47#_c_523_n 0.00290172f $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_268 N_A_193_47#_c_336_n N_A_476_47#_c_523_n 0.0191754f $X=2.59 $Y=0.87 $X2=0
+ $Y2=0
cc_269 N_A_193_47#_c_338_n N_A_476_47#_c_523_n 0.00414073f $X=2.372 $Y=0.705
+ $X2=0 $Y2=0
cc_270 N_A_193_47#_c_335_n N_A_476_47#_c_513_n 2.21473e-19 $X=2.38 $Y=0.87 $X2=0
+ $Y2=0
cc_271 N_A_193_47#_c_336_n N_A_476_47#_c_513_n 0.0199815f $X=2.59 $Y=0.87 $X2=0
+ $Y2=0
cc_272 N_A_193_47#_c_338_n N_A_476_47#_c_513_n 7.79765e-19 $X=2.372 $Y=0.705
+ $X2=0 $Y2=0
cc_273 N_A_193_47#_c_336_n N_A_476_47#_c_514_n 0.00299408f $X=2.59 $Y=0.87 $X2=0
+ $Y2=0
cc_274 N_A_193_47#_c_344_n N_A_476_47#_c_514_n 0.00165865f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_275 N_A_193_47#_c_337_n N_A_476_47#_c_514_n 0.0173781f $X=2.675 $Y=1.575
+ $X2=0 $Y2=0
cc_276 N_A_193_47#_M1003_g N_A_476_47#_c_520_n 0.00404596f $X=2.725 $Y=2.275
+ $X2=0 $Y2=0
cc_277 N_A_193_47#_c_343_n N_A_476_47#_c_520_n 0.0385017f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_278 N_A_193_47#_c_344_n N_A_476_47#_c_520_n 0.00171665f $X=2.76 $Y=1.74 $X2=0
+ $Y2=0
cc_279 N_A_193_47#_c_337_n N_A_476_47#_c_520_n 0.0113314f $X=2.675 $Y=1.575
+ $X2=0 $Y2=0
cc_280 N_A_193_47#_c_342_n N_VPWR_M1013_s 0.00514852f $X=2.505 $Y=2 $X2=0 $Y2=0
cc_281 N_A_193_47#_c_341_n N_VPWR_c_610_n 0.012721f $X=1.1 $Y=2.085 $X2=0 $Y2=0
cc_282 N_A_193_47#_c_341_n N_VPWR_c_615_n 0.0120336f $X=1.1 $Y=2.085 $X2=0 $Y2=0
cc_283 N_A_193_47#_c_342_n N_VPWR_c_615_n 0.00489589f $X=2.505 $Y=2 $X2=0 $Y2=0
cc_284 N_A_193_47#_M1003_g N_VPWR_c_616_n 0.00366111f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_285 N_A_193_47#_c_342_n N_VPWR_c_616_n 0.00701778f $X=2.505 $Y=2 $X2=0 $Y2=0
cc_286 N_A_193_47#_M1003_g N_VPWR_c_609_n 0.00547563f $X=2.725 $Y=2.275 $X2=0
+ $Y2=0
cc_287 N_A_193_47#_c_341_n N_VPWR_c_609_n 0.00743166f $X=1.1 $Y=2.085 $X2=0
+ $Y2=0
cc_288 N_A_193_47#_c_342_n N_VPWR_c_609_n 0.0221401f $X=2.505 $Y=2 $X2=0 $Y2=0
cc_289 N_A_193_47#_c_341_n N_VPWR_c_620_n 0.0119531f $X=1.1 $Y=2.085 $X2=0 $Y2=0
cc_290 N_A_193_47#_c_342_n N_VPWR_c_620_n 0.0252484f $X=2.505 $Y=2 $X2=0 $Y2=0
cc_291 N_A_193_47#_c_342_n A_381_369# 0.00588287f $X=2.505 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_292 N_A_193_47#_c_333_n N_VGND_c_703_n 0.00672221f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_293 N_A_193_47#_c_338_n N_VGND_c_703_n 0.00190318f $X=2.372 $Y=0.705 $X2=0
+ $Y2=0
cc_294 N_A_193_47#_c_333_n N_VGND_c_708_n 0.00730936f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_295 N_A_193_47#_c_334_n N_VGND_c_708_n 5.63036e-19 $X=1.082 $Y=0.91 $X2=0
+ $Y2=0
cc_296 N_A_193_47#_c_336_n N_VGND_c_709_n 0.00124133f $X=2.59 $Y=0.87 $X2=0
+ $Y2=0
cc_297 N_A_193_47#_c_338_n N_VGND_c_709_n 0.00500228f $X=2.372 $Y=0.705 $X2=0
+ $Y2=0
cc_298 N_A_193_47#_M1010_d N_VGND_c_711_n 0.00430317f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_299 N_A_193_47#_c_333_n N_VGND_c_711_n 0.00615829f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_300 N_A_193_47#_c_334_n N_VGND_c_711_n 9.46686e-19 $X=1.082 $Y=0.91 $X2=0
+ $Y2=0
cc_301 N_A_193_47#_c_336_n N_VGND_c_711_n 0.00244809f $X=2.59 $Y=0.87 $X2=0
+ $Y2=0
cc_302 N_A_193_47#_c_338_n N_VGND_c_711_n 0.00848363f $X=2.372 $Y=0.705 $X2=0
+ $Y2=0
cc_303 N_A_629_21#_c_452_n N_A_476_47#_c_509_n 0.00836312f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_304 N_A_629_21#_c_465_p N_A_476_47#_c_509_n 0.004107f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_305 N_A_629_21#_c_456_n N_A_476_47#_M1007_g 0.00407044f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_306 N_A_629_21#_c_452_n N_A_476_47#_M1007_g 0.00765951f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_307 N_A_629_21#_c_468_p N_A_476_47#_M1007_g 0.012841f $X=3.96 $Y=1.755 $X2=0
+ $Y2=0
cc_308 N_A_629_21#_c_465_p N_A_476_47#_c_510_n 0.00134898f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_309 N_A_629_21#_c_452_n N_A_476_47#_M1000_g 0.00103487f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_310 N_A_629_21#_M1005_g N_A_476_47#_c_511_n 0.0196785f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_311 N_A_629_21#_c_455_n N_A_476_47#_c_511_n 0.00564215f $X=3.835 $Y=1.7 $X2=0
+ $Y2=0
cc_312 N_A_629_21#_c_456_n N_A_476_47#_c_511_n 0.00731287f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_313 N_A_629_21#_c_452_n N_A_476_47#_c_511_n 0.0156359f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_314 N_A_629_21#_c_465_p N_A_476_47#_c_511_n 0.00423679f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_315 N_A_629_21#_c_468_p N_A_476_47#_c_511_n 0.00489524f $X=3.96 $Y=1.755
+ $X2=0 $Y2=0
cc_316 N_A_629_21#_c_452_n N_A_476_47#_c_512_n 0.0148261f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_317 N_A_629_21#_M1011_g N_A_476_47#_c_522_n 0.00475392f $X=3.22 $Y=2.275
+ $X2=0 $Y2=0
cc_318 N_A_629_21#_M1005_g N_A_476_47#_c_523_n 0.00148126f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_319 N_A_629_21#_M1005_g N_A_476_47#_c_513_n 0.0102149f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_320 N_A_629_21#_M1005_g N_A_476_47#_c_514_n 0.00629975f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_321 N_A_629_21#_M1005_g N_A_476_47#_c_520_n 0.0114592f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_322 N_A_629_21#_M1011_g N_A_476_47#_c_520_n 0.0108058f $X=3.22 $Y=2.275 $X2=0
+ $Y2=0
cc_323 N_A_629_21#_c_455_n N_A_476_47#_c_520_n 0.0193224f $X=3.835 $Y=1.7 $X2=0
+ $Y2=0
cc_324 N_A_629_21#_c_456_n N_A_476_47#_c_520_n 0.00911775f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_325 N_A_629_21#_c_468_p N_A_476_47#_c_520_n 0.00684055f $X=3.96 $Y=1.755
+ $X2=0 $Y2=0
cc_326 N_A_629_21#_M1005_g N_A_476_47#_c_515_n 0.0162449f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_327 N_A_629_21#_c_455_n N_A_476_47#_c_515_n 0.0238221f $X=3.835 $Y=1.7 $X2=0
+ $Y2=0
cc_328 N_A_629_21#_c_456_n N_A_476_47#_c_515_n 0.00748228f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_329 N_A_629_21#_c_452_n N_A_476_47#_c_515_n 0.0250354f $X=4.037 $Y=1.535
+ $X2=0 $Y2=0
cc_330 N_A_629_21#_M1011_g N_VPWR_c_611_n 0.00622935f $X=3.22 $Y=2.275 $X2=0
+ $Y2=0
cc_331 N_A_629_21#_c_455_n N_VPWR_c_611_n 0.00562825f $X=3.835 $Y=1.7 $X2=0
+ $Y2=0
cc_332 N_A_629_21#_c_456_n N_VPWR_c_611_n 0.00481721f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_333 N_A_629_21#_c_468_p N_VPWR_c_611_n 0.0145939f $X=3.96 $Y=1.755 $X2=0
+ $Y2=0
cc_334 N_A_629_21#_c_468_p N_VPWR_c_612_n 0.0152489f $X=3.96 $Y=1.755 $X2=0
+ $Y2=0
cc_335 N_A_629_21#_M1011_g N_VPWR_c_616_n 0.00526858f $X=3.22 $Y=2.275 $X2=0
+ $Y2=0
cc_336 N_A_629_21#_M1007_s N_VPWR_c_609_n 0.00210766f $X=3.835 $Y=1.485 $X2=0
+ $Y2=0
cc_337 N_A_629_21#_M1011_g N_VPWR_c_609_n 0.010697f $X=3.22 $Y=2.275 $X2=0 $Y2=0
cc_338 N_A_629_21#_c_455_n N_VPWR_c_609_n 0.0111384f $X=3.835 $Y=1.7 $X2=0 $Y2=0
cc_339 N_A_629_21#_c_456_n N_VPWR_c_609_n 0.00394376f $X=3.505 $Y=1.7 $X2=0
+ $Y2=0
cc_340 N_A_629_21#_c_468_p N_VPWR_c_609_n 0.0107834f $X=3.96 $Y=1.755 $X2=0
+ $Y2=0
cc_341 N_A_629_21#_M1005_g N_VGND_c_704_n 0.0113477f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_342 N_A_629_21#_c_465_p N_VGND_c_704_n 0.00727213f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_343 N_A_629_21#_c_465_p N_VGND_c_705_n 0.00872062f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_344 N_A_629_21#_M1005_g N_VGND_c_709_n 0.0046653f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_345 N_A_629_21#_M1008_s N_VGND_c_711_n 0.00232147f $X=3.835 $Y=0.235 $X2=0
+ $Y2=0
cc_346 N_A_629_21#_M1005_g N_VGND_c_711_n 0.00799591f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_347 N_A_629_21#_c_465_p N_VGND_c_711_n 0.00985818f $X=3.96 $Y=0.58 $X2=0
+ $Y2=0
cc_348 N_A_476_47#_M1007_g N_VPWR_c_611_n 0.00248972f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_476_47#_c_522_n N_VPWR_c_611_n 0.0133617f $X=3.015 $Y=2.34 $X2=0
+ $Y2=0
cc_350 N_A_476_47#_c_520_n N_VPWR_c_611_n 0.00839059f $X=3.1 $Y=2.255 $X2=0
+ $Y2=0
cc_351 N_A_476_47#_M1007_g N_VPWR_c_612_n 0.0054256f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_476_47#_M1007_g N_VPWR_c_613_n 0.00355205f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_476_47#_M1000_g N_VPWR_c_613_n 0.00355205f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_476_47#_c_512_n N_VPWR_c_613_n 0.00369023f $X=4.59 $Y=1.16 $X2=0
+ $Y2=0
cc_355 N_A_476_47#_c_522_n N_VPWR_c_616_n 0.0392604f $X=3.015 $Y=2.34 $X2=0
+ $Y2=0
cc_356 N_A_476_47#_M1000_g N_VPWR_c_617_n 0.00585385f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_476_47#_M1009_d N_VPWR_c_609_n 0.00216803f $X=2.38 $Y=2.065 $X2=0
+ $Y2=0
cc_358 N_A_476_47#_M1007_g N_VPWR_c_609_n 0.0109193f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_359 N_A_476_47#_M1000_g N_VPWR_c_609_n 0.0114913f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_476_47#_c_522_n N_VPWR_c_609_n 0.0306707f $X=3.015 $Y=2.34 $X2=0
+ $Y2=0
cc_361 N_A_476_47#_c_522_n N_VPWR_c_620_n 0.0060411f $X=3.015 $Y=2.34 $X2=0
+ $Y2=0
cc_362 N_A_476_47#_c_522_n A_560_413# 0.00670962f $X=3.015 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_363 N_A_476_47#_c_520_n A_560_413# 0.00218612f $X=3.1 $Y=2.255 $X2=-0.19
+ $Y2=-0.24
cc_364 N_A_476_47#_c_510_n N_Q_c_691_n 0.0309426f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A_476_47#_c_523_n N_VGND_c_703_n 0.00278933f $X=2.87 $Y=0.45 $X2=0
+ $Y2=0
cc_366 N_A_476_47#_c_509_n N_VGND_c_704_n 0.006368f $X=4.17 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A_476_47#_c_511_n N_VGND_c_704_n 0.00141221f $X=4.095 $Y=1.16 $X2=0
+ $Y2=0
cc_368 N_A_476_47#_c_523_n N_VGND_c_704_n 0.0109522f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_369 N_A_476_47#_c_515_n N_VGND_c_704_n 0.0120502f $X=3.695 $Y=1.16 $X2=0
+ $Y2=0
cc_370 N_A_476_47#_c_509_n N_VGND_c_705_n 0.00547395f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_371 N_A_476_47#_c_509_n N_VGND_c_706_n 0.0031786f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_476_47#_c_510_n N_VGND_c_706_n 0.0031786f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_476_47#_c_512_n N_VGND_c_706_n 0.0035554f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_476_47#_c_523_n N_VGND_c_709_n 0.0220682f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_375 N_A_476_47#_c_510_n N_VGND_c_710_n 0.00585385f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_476_47#_M1014_d N_VGND_c_711_n 0.00293225f $X=2.38 $Y=0.235 $X2=0
+ $Y2=0
cc_377 N_A_476_47#_c_509_n N_VGND_c_711_n 0.0110218f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A_476_47#_c_510_n N_VGND_c_711_n 0.0116795f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_476_47#_c_523_n N_VGND_c_711_n 0.0224235f $X=2.87 $Y=0.45 $X2=0 $Y2=0
cc_380 N_A_476_47#_c_523_n A_575_47# 0.00288367f $X=2.87 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_381 N_A_476_47#_c_513_n A_575_47# 6.59707e-19 $X=2.955 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_382 N_VPWR_c_609_n A_381_369# 0.00381236f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_383 N_VPWR_c_609_n A_560_413# 0.00280095f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_384 N_VPWR_c_609_n N_Q_M1000_d 0.002964f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_617_n Q 0.0177571f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_609_n Q 0.0108473f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_387 Q N_VGND_c_710_n 0.00913062f $X=4.77 $Y=0.425 $X2=0 $Y2=0
cc_388 N_Q_M1006_d N_VGND_c_711_n 0.00321007f $X=4.665 $Y=0.235 $X2=0 $Y2=0
cc_389 Q N_VGND_c_711_n 0.00983854f $X=4.77 $Y=0.425 $X2=0 $Y2=0
cc_390 N_VGND_c_711_n A_381_47# 0.00748004f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_391 N_VGND_c_711_n A_575_47# 0.00588947f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o21a_4.spice
* Created: Thu Aug 27 14:35:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21a_4.pex.spice"
.subckt sky130_fd_sc_hd__o21a_4  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_80_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1005_d N_A_80_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_A_80_21#_M1009_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_X_M1009_d N_A_80_21#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_80_21#_M1012_d N_B1_M1012_g N_A_475_47#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1019 N_A_80_21#_M1012_d N_B1_M1019_g N_A_475_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.117 PD=0.93 PS=1.01 NRD=0 NRS=14.76 M=1 R=4.33333
+ SA=75000.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_475_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.117 PD=1.01 PS=1.01 NRD=12.912 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_475_47#_M1010_d N_A2_M1010_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.117 PD=0.93 PS=1.01 NRD=0 NRS=1.836 M=1 R=4.33333 SA=75001.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1016 N_A_475_47#_M1010_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1016_s N_A1_M1017_g N_A_475_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_80_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_21#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75004
+ A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1002_d N_A_80_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75003.6
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A_80_21#_M1013_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1013_d N_B1_M1008_g N_A_80_21#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1014_d N_B1_M1014_g N_A_80_21#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.31 AS=0.14 PD=1.62 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1001 A_934_297# N_A1_M1001_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.31 PD=1.28 PS=1.62 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75003.1 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1015 N_A_80_21#_M1015_d N_A2_M1015_g A_934_297# VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75003.6 SB=75001.1
+ A=0.15 P=2.3 MULT=1
MM1004 N_A_80_21#_M1015_d N_A2_M1004_g A_762_297# VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75004 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1011 A_762_297# N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.285 PD=1.28 PS=2.57 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75004.4 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
c_82 VPB 0 1.78828e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o21a_4.pxi.spice"
*
.ends
*
*

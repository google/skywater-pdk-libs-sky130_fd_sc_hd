* File: sky130_fd_sc_hd__nor3_2.pxi.spice
* Created: Thu Aug 27 14:32:06 2020
* 
x_PM_SKY130_FD_SC_HD__NOR3_2%A N_A_c_55_n N_A_M1002_g N_A_M1000_g N_A_c_56_n
+ N_A_M1004_g N_A_M1009_g A A N_A_c_58_n PM_SKY130_FD_SC_HD__NOR3_2%A
x_PM_SKY130_FD_SC_HD__NOR3_2%B N_B_c_95_n N_B_M1001_g N_B_M1005_g N_B_c_96_n
+ N_B_M1003_g N_B_M1007_g B B N_B_c_98_n PM_SKY130_FD_SC_HD__NOR3_2%B
x_PM_SKY130_FD_SC_HD__NOR3_2%C N_C_c_142_n N_C_M1010_g N_C_M1006_g N_C_c_143_n
+ N_C_M1011_g N_C_M1008_g C C N_C_c_168_p N_C_c_145_n N_C_c_146_n
+ PM_SKY130_FD_SC_HD__NOR3_2%C
x_PM_SKY130_FD_SC_HD__NOR3_2%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1009_s
+ N_A_27_297#_M1007_d N_A_27_297#_c_188_n N_A_27_297#_c_208_p
+ N_A_27_297#_c_189_n N_A_27_297#_c_209_p N_A_27_297#_c_190_n
+ N_A_27_297#_c_191_n N_A_27_297#_c_192_n PM_SKY130_FD_SC_HD__NOR3_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR3_2%VPWR N_VPWR_M1000_d N_VPWR_c_224_n VPWR
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_223_n N_VPWR_c_228_n
+ PM_SKY130_FD_SC_HD__NOR3_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR3_2%A_281_297# N_A_281_297#_M1005_s
+ N_A_281_297#_M1006_d N_A_281_297#_M1008_d N_A_281_297#_c_274_n
+ N_A_281_297#_c_264_n N_A_281_297#_c_284_n N_A_281_297#_c_267_n
+ N_A_281_297#_c_265_n N_A_281_297#_c_293_p N_A_281_297#_c_288_n
+ PM_SKY130_FD_SC_HD__NOR3_2%A_281_297#
x_PM_SKY130_FD_SC_HD__NOR3_2%Y N_Y_M1002_s N_Y_M1001_d N_Y_M1010_s N_Y_M1006_s
+ N_Y_c_302_n N_Y_c_295_n N_Y_c_296_n N_Y_c_310_n N_Y_c_297_n N_Y_c_325_n
+ N_Y_c_298_n N_Y_c_299_n Y N_Y_c_344_n PM_SKY130_FD_SC_HD__NOR3_2%Y
x_PM_SKY130_FD_SC_HD__NOR3_2%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1003_s
+ N_VGND_M1010_d N_VGND_M1011_d N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n
+ N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n VGND
+ N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n
+ PM_SKY130_FD_SC_HD__NOR3_2%VGND
cc_1 VNB N_A_c_55_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_56_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB A 0.0161137f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_A_c_58_n 0.0382849f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_5 VNB N_B_c_95_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_96_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_7 VNB B 0.0156327f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_B_c_98_n 0.0365012f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_9 VNB N_C_c_142_n 0.0214684f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_C_c_143_n 0.0198049f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_11 VNB C 3.24615e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_12 VNB N_C_c_145_n 0.0404997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_C_c_146_n 0.00465382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_223_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_15 VNB N_Y_c_295_n 0.00338427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_296_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_297_n 0.0167605f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_18 VNB N_Y_c_298_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_299_n 0.0132181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB Y 0.0197285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_370_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_22 VNB N_VGND_c_371_n 0.0344379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_372_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_24 VNB N_VGND_c_373_n 0.0118683f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_25 VNB N_VGND_c_374_n 0.0181293f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_26 VNB N_VGND_c_375_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_376_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_377_n 0.0166866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_378_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_379_n 0.0263734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_380_n 0.19896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_M1000_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_33 VPB N_A_M1009_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_34 VPB N_A_c_58_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_35 VPB N_B_M1005_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_36 VPB N_B_M1007_g 0.0229477f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_37 VPB N_B_c_98_n 0.00440018f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_38 VPB N_C_M1006_g 0.0229841f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_39 VPB N_C_M1008_g 0.0228354f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_40 VPB C 0.00290811f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_41 VPB N_C_c_145_n 0.00448221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_297#_c_188_n 0.00371072f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_43 VPB N_A_27_297#_c_189_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_297#_c_190_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_297#_c_191_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_297#_c_192_n 0.00268826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_224_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_48 VPB N_VPWR_c_225_n 0.0180608f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_49 VPB N_VPWR_c_226_n 0.0709757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_223_n 0.0526883f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_51 VPB N_VPWR_c_228_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_52 VPB N_A_281_297#_c_264_n 0.0128761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_281_297#_c_265_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB Y 0.0236791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_A_c_56_n N_B_c_95_n 0.0194931f $X=0.91 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_56 N_A_M1009_g N_B_M1005_g 0.0194931f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_57 A B 0.0185436f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_58_n B 0.00160637f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_59 A N_B_c_98_n 2.03927e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A_c_58_n N_B_c_98_n 0.0194931f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_61 A N_A_27_297#_c_188_n 0.021852f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_A_27_297#_c_189_n 0.0134951f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1009_g N_A_27_297#_c_189_n 0.0134675f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_64 A N_A_27_297#_c_189_n 0.0396361f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_c_58_n N_A_27_297#_c_189_n 0.00211509f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_M1000_g N_VPWR_c_224_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1009_g N_VPWR_c_224_n 0.00302074f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_68 N_A_M1000_g N_VPWR_c_225_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_M1009_g N_VPWR_c_226_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_VPWR_c_223_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_71 N_A_M1009_g N_VPWR_c_223_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_c_55_n N_Y_c_302_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_56_n N_Y_c_302_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A_c_56_n N_Y_c_295_n 0.00890517f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_75 A N_Y_c_295_n 0.00688575f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_55_n N_Y_c_296_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_c_56_n N_Y_c_296_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_78 A N_Y_c_296_n 0.0266272f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_58_n N_Y_c_296_n 0.00230339f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_56_n N_Y_c_310_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_55_n N_VGND_c_371_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_82 A N_VGND_c_371_n 0.019624f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_c_56_n N_VGND_c_372_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_c_55_n N_VGND_c_375_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_c_56_n N_VGND_c_375_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_c_55_n N_VGND_c_380_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_c_56_n N_VGND_c_380_n 0.0057435f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B_M1007_g C 3.95514e-19 $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_89 N_B_c_98_n C 0.00427961f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_90 B N_C_c_145_n 9.27479e-19 $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_91 B N_C_c_146_n 0.0178149f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_92 N_B_c_98_n N_C_c_146_n 7.64149e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_M1005_g N_A_27_297#_c_190_n 0.0132199f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_94 N_B_M1007_g N_A_27_297#_c_190_n 0.0112055f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_95 B N_A_27_297#_c_190_n 0.0417417f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B_c_98_n N_A_27_297#_c_190_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_97 B N_A_27_297#_c_191_n 0.00942636f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_98 B N_A_27_297#_c_192_n 0.0213978f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B_M1005_g N_VPWR_c_226_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B_M1007_g N_VPWR_c_226_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B_M1005_g N_VPWR_c_223_n 0.0106871f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B_M1007_g N_VPWR_c_223_n 0.00660224f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B_M1007_g N_A_281_297#_c_264_n 0.0119904f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_A_281_297#_c_267_n 0.00417384f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B_c_95_n N_Y_c_302_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_95_n N_Y_c_295_n 0.00865686f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_107 B N_Y_c_295_n 0.0174927f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_108 N_B_c_95_n N_Y_c_310_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_c_96_n N_Y_c_310_n 0.0109565f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B_c_96_n N_Y_c_297_n 0.0109318f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_111 B N_Y_c_297_n 0.0359387f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B_c_95_n N_Y_c_298_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_96_n N_Y_c_298_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_114 B N_Y_c_298_n 0.0266272f $X=1.99 $Y=1.105 $X2=0 $Y2=0
cc_115 N_B_c_98_n N_Y_c_298_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B_c_95_n N_VGND_c_372_n 0.00146339f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_95_n N_VGND_c_378_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B_c_96_n N_VGND_c_378_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B_c_96_n N_VGND_c_379_n 0.00336341f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B_c_95_n N_VGND_c_380_n 0.0057435f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_96_n N_VGND_c_380_n 0.0070399f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_122 N_C_M1006_g N_A_27_297#_c_192_n 0.00526396f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_123 C N_A_27_297#_c_192_n 0.00971294f $X=2.47 $Y=1.445 $X2=0 $Y2=0
cc_124 N_C_M1006_g N_VPWR_c_226_n 0.00357877f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_125 N_C_M1008_g N_VPWR_c_226_n 0.00357877f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_126 N_C_M1006_g N_VPWR_c_223_n 0.00655123f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_127 N_C_M1008_g N_VPWR_c_223_n 0.00624775f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_128 C N_A_281_297#_M1006_d 0.00494976f $X=2.47 $Y=1.445 $X2=0 $Y2=0
cc_129 C N_A_281_297#_c_264_n 0.0010936f $X=2.47 $Y=1.445 $X2=0 $Y2=0
cc_130 C N_A_281_297#_c_267_n 0.0143639f $X=2.47 $Y=1.445 $X2=0 $Y2=0
cc_131 N_C_M1006_g N_A_281_297#_c_265_n 0.011972f $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_132 N_C_M1008_g N_A_281_297#_c_265_n 0.00988743f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C_c_142_n N_Y_c_297_n 0.0109316f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_134 N_C_c_168_p N_Y_c_297_n 0.0231006f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_135 N_C_c_146_n N_Y_c_297_n 0.0220432f $X=2.507 $Y=1.285 $X2=0 $Y2=0
cc_136 N_C_c_142_n N_Y_c_325_n 0.0110885f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C_c_143_n N_Y_c_325_n 0.0110634f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C_c_142_n N_Y_c_299_n 0.00127098f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C_c_143_n N_Y_c_299_n 0.0120145f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C_c_145_n N_Y_c_299_n 0.00222133f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C_c_142_n Y 4.73214e-19 $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C_M1006_g Y 6.50781e-19 $X=2.71 $Y=1.985 $X2=0 $Y2=0
cc_143 N_C_c_143_n Y 0.00409446f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_144 N_C_M1008_g Y 0.0183118f $X=3.13 $Y=1.985 $X2=0 $Y2=0
cc_145 C Y 0.012011f $X=2.47 $Y=1.445 $X2=0 $Y2=0
cc_146 N_C_c_168_p Y 0.026269f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_147 N_C_c_145_n Y 0.0190383f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_148 N_C_c_143_n N_VGND_c_374_n 0.00323103f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_149 N_C_c_142_n N_VGND_c_377_n 0.0042235f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_150 N_C_c_143_n N_VGND_c_377_n 0.0042235f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_151 N_C_c_142_n N_VGND_c_379_n 0.00336341f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C_c_142_n N_VGND_c_380_n 0.00705454f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_153 N_C_c_143_n N_VGND_c_380_n 0.00675353f $X=3.13 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_27_297#_c_189_n N_VPWR_M1000_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_155 N_A_27_297#_c_189_n N_VPWR_c_224_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_156 N_A_27_297#_c_208_p N_VPWR_c_225_n 0.0161885f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_157 N_A_27_297#_c_209_p N_VPWR_c_226_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_158 N_A_27_297#_M1000_s N_VPWR_c_223_n 0.00315976f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_159 N_A_27_297#_M1009_s N_VPWR_c_223_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_27_297#_M1007_d N_VPWR_c_223_n 0.00226545f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_161 N_A_27_297#_c_208_p N_VPWR_c_223_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_162 N_A_27_297#_c_209_p N_VPWR_c_223_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_163 N_A_27_297#_c_190_n N_A_281_297#_M1005_s 0.00165831f $X=1.835 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_164 N_A_27_297#_c_190_n N_A_281_297#_c_274_n 0.0126766f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_165 N_A_27_297#_M1007_d N_A_281_297#_c_264_n 0.00593473f $X=1.825 $Y=1.485
+ $X2=0 $Y2=0
cc_166 N_A_27_297#_c_190_n N_A_281_297#_c_264_n 0.00320918f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_167 N_A_27_297#_c_192_n N_A_281_297#_c_264_n 0.0153739f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_168 N_A_27_297#_c_192_n N_A_281_297#_c_267_n 0.0153956f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_169 N_A_27_297#_c_189_n N_Y_c_295_n 8.37688e-19 $X=0.995 $Y=1.54 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_191_n N_Y_c_295_n 0.00524452f $X=1.12 $Y=1.62 $X2=0 $Y2=0
cc_171 N_VPWR_c_223_n N_A_281_297#_M1005_s 0.00246446f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_172 N_VPWR_c_223_n N_A_281_297#_M1006_d 0.00209324f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_223_n N_A_281_297#_M1008_d 0.0020932f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_226_n N_A_281_297#_c_264_n 0.0455751f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_223_n N_A_281_297#_c_264_n 0.02717f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_176 N_VPWR_c_226_n N_A_281_297#_c_284_n 0.0142933f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_223_n N_A_281_297#_c_284_n 0.00962421f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_226_n N_A_281_297#_c_265_n 0.0489446f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_223_n N_A_281_297#_c_265_n 0.0300869f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_226_n N_A_281_297#_c_288_n 0.0131175f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_223_n N_A_281_297#_c_288_n 0.00808434f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_223_n N_Y_M1006_s 0.00216833f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_183 N_A_281_297#_c_265_n N_Y_M1006_s 0.00312348f $X=3.215 $Y=2.38 $X2=0 $Y2=0
cc_184 N_A_281_297#_M1008_d Y 0.00276279f $X=3.205 $Y=1.485 $X2=0 $Y2=0
cc_185 N_A_281_297#_c_265_n Y 0.00320918f $X=3.215 $Y=2.38 $X2=0 $Y2=0
cc_186 N_A_281_297#_c_293_p Y 0.0164145f $X=3.34 $Y=1.96 $X2=0 $Y2=0
cc_187 N_A_281_297#_c_265_n N_Y_c_344_n 0.0116103f $X=3.215 $Y=2.38 $X2=0 $Y2=0
cc_188 N_Y_c_295_n N_VGND_M1004_d 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_189 N_Y_c_297_n N_VGND_M1003_s 0.00281828f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_190 N_Y_c_297_n N_VGND_M1010_d 0.00281828f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_191 N_Y_c_299_n N_VGND_M1011_d 0.0028133f $X=3.365 $Y=0.905 $X2=0 $Y2=0
cc_192 N_Y_c_296_n N_VGND_c_371_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_193 N_Y_c_295_n N_VGND_c_372_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_194 N_Y_c_299_n N_VGND_c_373_n 7.67289e-19 $X=3.365 $Y=0.905 $X2=0 $Y2=0
cc_195 N_Y_c_299_n N_VGND_c_374_n 0.0223917f $X=3.365 $Y=0.905 $X2=0 $Y2=0
cc_196 N_Y_c_302_n N_VGND_c_375_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_197 N_Y_c_295_n N_VGND_c_375_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_198 N_Y_c_297_n N_VGND_c_377_n 0.00400646f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_199 N_Y_c_325_n N_VGND_c_377_n 0.0185141f $X=2.92 $Y=0.39 $X2=0 $Y2=0
cc_200 N_Y_c_295_n N_VGND_c_378_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_201 N_Y_c_310_n N_VGND_c_378_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_202 N_Y_c_297_n N_VGND_c_378_n 0.00198695f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_203 N_Y_c_297_n N_VGND_c_379_n 0.0552675f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_204 N_Y_M1002_s N_VGND_c_380_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_205 N_Y_M1001_d N_VGND_c_380_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_206 N_Y_M1010_s N_VGND_c_380_n 0.00215201f $X=2.785 $Y=0.235 $X2=0 $Y2=0
cc_207 N_Y_c_302_n N_VGND_c_380_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_208 N_Y_c_295_n N_VGND_c_380_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_209 N_Y_c_310_n N_VGND_c_380_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_210 N_Y_c_297_n N_VGND_c_380_n 0.014311f $X=2.755 $Y=0.815 $X2=0 $Y2=0
cc_211 N_Y_c_325_n N_VGND_c_380_n 0.0121046f $X=2.92 $Y=0.39 $X2=0 $Y2=0
cc_212 N_Y_c_299_n N_VGND_c_380_n 0.00246308f $X=3.365 $Y=0.905 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__mux2_1.spice
* Created: Thu Aug 27 14:27:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__mux2_1.pex.spice"
.subckt sky130_fd_sc_hd__mux2_1  VNB VPB S A1 A0 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_76_199#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.137107 AS=0.169 PD=1.26963 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1004 A_218_47# N_S_M1004_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0885925 PD=0.75 PS=0.820374 NRD=31.428 NRS=34.284 M=1 R=2.8 SA=75000.7
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_76_199#_M1005_d N_A1_M1005_g A_218_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.09975 AS=0.0693 PD=0.895 PS=0.75 NRD=1.428 NRS=31.428 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1011 A_439_47# N_A0_M1011_g N_A_76_199#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.09975 PD=0.75 PS=0.895 NRD=31.428 NRS=54.276 M=1 R=2.8
+ SA=75001.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_505_21#_M1000_g A_439_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0693 PD=1.11 PS=0.75 NRD=21.42 NRS=31.428 M=1 R=2.8 SA=75002.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 N_A_505_21#_M1008_d N_S_M1008_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1449 PD=1.36 PS=1.11 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_76_199#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.223028 AS=0.26 PD=1.96479 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1003 A_218_374# N_S_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07665 AS=0.0936718 PD=0.785 PS=0.825211 NRD=59.7895 NRS=57.4452 M=1 R=2.8
+ SA=75000.7 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_76_199#_M1001_d N_A0_M1001_g A_218_374# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1932 AS=0.07665 PD=1.34 PS=0.785 NRD=53.9386 NRS=59.7895 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 A_535_374# N_A1_M1006_g N_A_76_199#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1932 PD=0.63 PS=1.34 NRD=23.443 NRS=70.3487 M=1 R=2.8
+ SA=75002.3 SB=75001 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_505_21#_M1002_g A_535_374# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0693 AS=0.0441 PD=0.75 PS=0.63 NRD=21.0987 NRS=23.443 M=1 R=2.8
+ SA=75002.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_505_21#_M1009_d N_S_M1009_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0693 PD=1.4 PS=0.75 NRD=0 NRS=2.3443 M=1 R=2.8 SA=75003.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_38 VNB 0 1.9931e-19 $X=0.42 $Y=-0.085
*
.include "sky130_fd_sc_hd__mux2_1.pxi.spice"
*
.ends
*
*

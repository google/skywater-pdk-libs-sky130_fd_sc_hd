* File: sky130_fd_sc_hd__or2b_4.pxi.spice
* Created: Thu Aug 27 14:43:10 2020
* 
x_PM_SKY130_FD_SC_HD__OR2B_4%B_N N_B_N_M1002_g N_B_N_M1005_g B_N B_N B_N
+ N_B_N_c_77_n PM_SKY130_FD_SC_HD__OR2B_4%B_N
x_PM_SKY130_FD_SC_HD__OR2B_4%A_27_53# N_A_27_53#_M1002_s N_A_27_53#_M1005_d
+ N_A_27_53#_c_99_n N_A_27_53#_M1012_g N_A_27_53#_M1007_g N_A_27_53#_c_100_n
+ N_A_27_53#_c_101_n N_A_27_53#_c_102_n N_A_27_53#_c_103_n N_A_27_53#_c_104_n
+ N_A_27_53#_c_105_n N_A_27_53#_c_110_n PM_SKY130_FD_SC_HD__OR2B_4%A_27_53#
x_PM_SKY130_FD_SC_HD__OR2B_4%A N_A_M1010_g N_A_M1008_g A N_A_c_158_n N_A_c_159_n
+ PM_SKY130_FD_SC_HD__OR2B_4%A
x_PM_SKY130_FD_SC_HD__OR2B_4%A_219_297# N_A_219_297#_M1012_d
+ N_A_219_297#_M1007_s N_A_219_297#_c_190_n N_A_219_297#_M1003_g
+ N_A_219_297#_M1000_g N_A_219_297#_c_191_n N_A_219_297#_M1004_g
+ N_A_219_297#_M1001_g N_A_219_297#_c_192_n N_A_219_297#_M1006_g
+ N_A_219_297#_M1011_g N_A_219_297#_c_193_n N_A_219_297#_M1009_g
+ N_A_219_297#_M1013_g N_A_219_297#_c_201_n N_A_219_297#_c_194_n
+ N_A_219_297#_c_215_n N_A_219_297#_c_203_n N_A_219_297#_c_234_n
+ N_A_219_297#_c_204_n N_A_219_297#_c_268_p N_A_219_297#_c_205_n
+ N_A_219_297#_c_195_n N_A_219_297#_c_196_n
+ PM_SKY130_FD_SC_HD__OR2B_4%A_219_297#
x_PM_SKY130_FD_SC_HD__OR2B_4%VPWR N_VPWR_M1005_s N_VPWR_M1008_d N_VPWR_M1001_s
+ N_VPWR_M1013_s N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n VPWR
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_313_n
+ PM_SKY130_FD_SC_HD__OR2B_4%VPWR
x_PM_SKY130_FD_SC_HD__OR2B_4%X N_X_M1003_d N_X_M1006_d N_X_M1000_d N_X_M1011_d
+ N_X_c_380_n N_X_c_417_n N_X_c_383_n N_X_c_371_n N_X_c_372_n N_X_c_395_n
+ N_X_c_419_n N_X_c_376_n N_X_c_373_n N_X_c_401_n N_X_c_377_n N_X_c_374_n X
+ PM_SKY130_FD_SC_HD__OR2B_4%X
x_PM_SKY130_FD_SC_HD__OR2B_4%VGND N_VGND_M1002_d N_VGND_M1010_d N_VGND_M1004_s
+ N_VGND_M1009_s N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n VGND N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ PM_SKY130_FD_SC_HD__OR2B_4%VGND
cc_1 VNB N_B_N_M1002_g 0.0403802f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB B_N 0.00936139f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_B_N_c_77_n 0.0382319f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_53#_c_99_n 0.019479f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_5 VNB N_A_27_53#_c_100_n 0.0317458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_53#_c_101_n 0.0136901f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_7 VNB N_A_27_53#_c_102_n 0.0195877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_53#_c_103_n 0.00233375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_104_n 0.00923383f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_10 VNB N_A_27_53#_c_105_n 0.0126651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB A 0.00812666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_c_158_n 0.0228975f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.785
cc_13 VNB N_A_c_159_n 0.0169647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_219_297#_c_190_n 0.016768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_15 VNB N_A_219_297#_c_191_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_219_297#_c_192_n 0.0157965f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_17 VNB N_A_219_297#_c_193_n 0.0191453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_219_297#_c_194_n 0.00212928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_219_297#_c_195_n 0.00306363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_219_297#_c_196_n 0.0644875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_313_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_371_n 0.00217862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_372_n 0.00291109f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.53
cc_24 VNB N_X_c_373_n 0.0100824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_374_n 0.00222314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0230536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_444_n 0.00613174f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_VGND_c_445_n 0.00360321f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_29 VNB N_VGND_c_446_n 0.00417234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_447_n 0.0177475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_448_n 0.00324283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_449_n 0.0171196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_450_n 0.00324283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_451_n 0.0200255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_452_n 0.0110503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_453_n 0.222559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_454_n 0.0174489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_455_n 0.020655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_456_n 0.00336608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_B_N_M1005_g 0.0666208f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_41 VPB B_N 0.0295284f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_42 VPB N_B_N_c_77_n 0.0100629f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_43 VPB N_A_27_53#_M1007_g 0.0223366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_53#_c_100_n 0.0124541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_53#_c_101_n 0.00249896f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_46 VPB N_A_27_53#_c_105_n 0.00999504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_53#_c_110_n 0.015111f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.53
cc_48 VPB N_A_M1008_g 0.0186453f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_49 VPB N_A_c_158_n 0.00407197f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.785
cc_50 VPB N_A_219_297#_M1000_g 0.0191174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_219_297#_M1001_g 0.0177993f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_52 VPB N_A_219_297#_M1011_g 0.0180899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_219_297#_M1013_g 0.0219253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_219_297#_c_201_n 0.0106203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_219_297#_c_194_n 0.00176706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_219_297#_c_203_n 0.00688428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_219_297#_c_204_n 0.0011175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_219_297#_c_205_n 0.00261924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_219_297#_c_196_n 0.0104024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_315_n 0.0190905f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_62 VPB N_VPWR_c_316_n 0.00471615f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_63 VPB N_VPWR_c_317_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_318_n 0.0154369f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.87
cc_65 VPB N_VPWR_c_319_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_320_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_321_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_322_n 0.0437467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_323_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_324_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_313_n 0.0565283f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_376_n 8.02457e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_377_n 0.00431973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB X 0.0218764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 N_B_N_c_77_n N_A_27_53#_c_100_n 0.0116586f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B_N_M1002_g N_A_27_53#_c_102_n 0.0125629f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_77 N_B_N_M1002_g N_A_27_53#_c_103_n 0.0139789f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_78 N_B_N_M1002_g N_A_27_53#_c_104_n 0.00412742f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_79 B_N N_A_27_53#_c_104_n 0.0273927f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_80 N_B_N_c_77_n N_A_27_53#_c_104_n 0.00728523f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B_N_M1002_g N_A_27_53#_c_105_n 0.00866774f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_82 B_N N_A_27_53#_c_105_n 0.0206572f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B_N_M1005_g N_A_27_53#_c_110_n 0.0195028f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_84 B_N N_A_27_53#_c_110_n 0.0473214f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_85 N_B_N_M1005_g N_VPWR_c_315_n 0.00450113f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_86 B_N N_VPWR_c_315_n 0.0223212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B_N_M1005_g N_VPWR_c_322_n 0.00585385f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_88 N_B_N_M1005_g N_VPWR_c_313_n 0.0120826f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_89 B_N N_VPWR_c_313_n 0.00407169f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B_N_M1002_g N_VGND_c_453_n 0.0073571f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_91 N_B_N_M1002_g N_VGND_c_454_n 0.00402941f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_92 N_B_N_M1002_g N_VGND_c_455_n 0.00501457f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_93 N_A_27_53#_M1007_g N_A_M1008_g 0.0498091f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_27_53#_c_101_n A 0.00143049f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_101_n N_A_c_158_n 0.0498091f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_27_53#_c_99_n N_A_c_159_n 0.011608f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_27_53#_M1007_g N_A_219_297#_c_201_n 0.0194691f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_98 N_A_27_53#_c_110_n N_A_219_297#_c_201_n 0.056389f $X=0.68 $Y=2.2 $X2=0
+ $Y2=0
cc_99 N_A_27_53#_c_99_n N_A_219_297#_c_194_n 0.0027318f $X=1.37 $Y=0.995 $X2=0
+ $Y2=0
cc_100 N_A_27_53#_M1007_g N_A_219_297#_c_194_n 0.00446933f $X=1.43 $Y=1.985
+ $X2=0 $Y2=0
cc_101 N_A_27_53#_c_100_n N_A_219_297#_c_194_n 0.00459671f $X=1.295 $Y=1.16
+ $X2=0 $Y2=0
cc_102 N_A_27_53#_c_101_n N_A_219_297#_c_194_n 0.00972263f $X=1.4 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_53#_c_105_n N_A_219_297#_c_194_n 0.0246012f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_104 N_A_27_53#_c_110_n N_A_219_297#_c_194_n 0.00410296f $X=0.68 $Y=2.2 $X2=0
+ $Y2=0
cc_105 N_A_27_53#_c_99_n N_A_219_297#_c_215_n 0.0105803f $X=1.37 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_27_53#_M1007_g N_A_219_297#_c_203_n 0.00515613f $X=1.43 $Y=1.985
+ $X2=0 $Y2=0
cc_107 N_A_27_53#_M1007_g N_A_219_297#_c_205_n 0.00226926f $X=1.43 $Y=1.985
+ $X2=0 $Y2=0
cc_108 N_A_27_53#_c_100_n N_A_219_297#_c_205_n 0.00858393f $X=1.295 $Y=1.16
+ $X2=0 $Y2=0
cc_109 N_A_27_53#_c_105_n N_A_219_297#_c_205_n 0.0109731f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_110 N_A_27_53#_c_110_n N_A_219_297#_c_205_n 0.0102314f $X=0.68 $Y=2.2 $X2=0
+ $Y2=0
cc_111 N_A_27_53#_c_99_n N_A_219_297#_c_195_n 0.00802177f $X=1.37 $Y=0.995 $X2=0
+ $Y2=0
cc_112 N_A_27_53#_c_101_n N_A_219_297#_c_195_n 0.00160921f $X=1.4 $Y=1.16 $X2=0
+ $Y2=0
cc_113 N_A_27_53#_c_105_n N_A_219_297#_c_195_n 0.00807051f $X=0.68 $Y=1.325
+ $X2=0 $Y2=0
cc_114 N_A_27_53#_M1007_g N_VPWR_c_322_n 0.00427501f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_27_53#_c_110_n N_VPWR_c_322_n 0.0116048f $X=0.68 $Y=2.2 $X2=0 $Y2=0
cc_116 N_A_27_53#_M1005_d N_VPWR_c_313_n 0.00615334f $X=0.545 $Y=2.065 $X2=0
+ $Y2=0
cc_117 N_A_27_53#_M1007_g N_VPWR_c_313_n 0.00811782f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_27_53#_c_110_n N_VPWR_c_313_n 0.00646998f $X=0.68 $Y=2.2 $X2=0 $Y2=0
cc_119 N_A_27_53#_c_99_n N_VGND_c_451_n 0.00426291f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_27_53#_c_99_n N_VGND_c_453_n 0.00708878f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_27_53#_c_102_n N_VGND_c_453_n 0.0116656f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_27_53#_c_103_n N_VGND_c_453_n 0.00384815f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_123 N_A_27_53#_c_105_n N_VGND_c_453_n 0.00106095f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_124 N_A_27_53#_c_102_n N_VGND_c_454_n 0.0183741f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_27_53#_c_103_n N_VGND_c_454_n 0.00229799f $X=0.595 $Y=0.82 $X2=0
+ $Y2=0
cc_126 N_A_27_53#_c_99_n N_VGND_c_455_n 0.00479981f $X=1.37 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_27_53#_c_100_n N_VGND_c_455_n 0.00574579f $X=1.295 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_27_53#_c_105_n N_VGND_c_455_n 0.0327468f $X=0.68 $Y=1.325 $X2=0 $Y2=0
cc_129 N_A_c_159_n N_A_219_297#_c_190_n 0.0183064f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_M1008_g N_A_219_297#_M1000_g 0.0328803f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_M1008_g N_A_219_297#_c_201_n 0.00334483f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_132 A N_A_219_297#_c_194_n 0.0159946f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_133 N_A_c_158_n N_A_219_297#_c_194_n 0.00174778f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_159_n N_A_219_297#_c_194_n 0.00165315f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_159_n N_A_219_297#_c_215_n 0.00547876f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_M1008_g N_A_219_297#_c_203_n 0.0148546f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_137 A N_A_219_297#_c_203_n 0.0501285f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_c_158_n N_A_219_297#_c_203_n 0.00285374f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_139 A N_A_219_297#_c_234_n 0.0143219f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_140 A N_A_219_297#_c_204_n 0.00217775f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A_c_158_n N_A_219_297#_c_204_n 2.16197e-19 $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_142 A N_A_219_297#_c_195_n 0.00939662f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_c_159_n N_A_219_297#_c_195_n 0.0026861f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_144 A N_A_219_297#_c_196_n 0.0136794f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_c_158_n N_A_219_297#_c_196_n 0.0218305f $X=1.85 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_VPWR_c_316_n 0.00620055f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1008_g N_VPWR_c_322_n 0.00585385f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1008_g N_VPWR_c_313_n 0.0107512f $X=1.79 $Y=1.985 $X2=0 $Y2=0
cc_149 A N_VGND_c_444_n 0.0147599f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_c_159_n N_VGND_c_444_n 0.00865803f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_159_n N_VGND_c_451_n 0.00543342f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_159_n N_VGND_c_453_n 0.00992834f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_219_297#_c_203_n N_VPWR_M1008_d 0.00268898f $X=2.49 $Y=1.53 $X2=0
+ $Y2=0
cc_154 N_A_219_297#_M1000_g N_VPWR_c_316_n 0.00170728f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_219_297#_c_203_n N_VPWR_c_316_n 0.0151808f $X=2.49 $Y=1.53 $X2=0
+ $Y2=0
cc_156 N_A_219_297#_M1001_g N_VPWR_c_317_n 0.00157837f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_219_297#_M1011_g N_VPWR_c_317_n 0.00157837f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_219_297#_M1013_g N_VPWR_c_319_n 0.00338128f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_159 N_A_219_297#_M1000_g N_VPWR_c_320_n 0.00585385f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_219_297#_M1001_g N_VPWR_c_320_n 0.00585385f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_161 N_A_219_297#_c_201_n N_VPWR_c_322_n 0.0308118f $X=1.22 $Y=1.63 $X2=0
+ $Y2=0
cc_162 N_A_219_297#_M1011_g N_VPWR_c_323_n 0.00585385f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_219_297#_M1013_g N_VPWR_c_323_n 0.00585385f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_219_297#_M1007_s N_VPWR_c_313_n 0.00209319f $X=1.095 $Y=1.485 $X2=0
+ $Y2=0
cc_165 N_A_219_297#_M1000_g N_VPWR_c_313_n 0.0106265f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_219_297#_M1001_g N_VPWR_c_313_n 0.00588483f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_219_297#_M1011_g N_VPWR_c_313_n 0.00588483f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_219_297#_M1013_g N_VPWR_c_313_n 0.0114944f $X=3.54 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_219_297#_c_201_n N_VPWR_c_313_n 0.0174754f $X=1.22 $Y=1.63 $X2=0
+ $Y2=0
cc_170 N_A_219_297#_c_203_n A_301_297# 0.00366293f $X=2.49 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_219_297#_c_203_n N_X_M1000_d 0.00167564f $X=2.49 $Y=1.53 $X2=0 $Y2=0
cc_172 N_A_219_297#_c_190_n N_X_c_380_n 0.00496583f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_219_297#_c_191_n N_X_c_380_n 0.00619772f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_219_297#_c_192_n N_X_c_380_n 5.54467e-19 $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_219_297#_c_203_n N_X_c_383_n 0.0132239f $X=2.49 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_219_297#_c_196_n N_X_c_383_n 2.80046e-19 $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_219_297#_c_191_n N_X_c_371_n 0.00844712f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_219_297#_c_192_n N_X_c_371_n 0.00850187f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_219_297#_c_234_n N_X_c_371_n 3.39565e-19 $X=2.575 $Y=1.245 $X2=0
+ $Y2=0
cc_180 N_A_219_297#_c_268_p N_X_c_371_n 0.0351744f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_219_297#_c_196_n N_X_c_371_n 0.00221825f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_219_297#_c_190_n N_X_c_372_n 0.00281545f $X=2.28 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_219_297#_c_191_n N_X_c_372_n 0.00110328f $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_219_297#_c_203_n N_X_c_372_n 0.00590182f $X=2.49 $Y=1.53 $X2=0 $Y2=0
cc_185 N_A_219_297#_c_234_n N_X_c_372_n 0.0142226f $X=2.575 $Y=1.245 $X2=0 $Y2=0
cc_186 N_A_219_297#_c_196_n N_X_c_372_n 0.00256683f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_219_297#_c_191_n N_X_c_395_n 5.54467e-19 $X=2.7 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_219_297#_c_192_n N_X_c_395_n 0.00619772f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_219_297#_c_193_n N_X_c_395_n 0.0111919f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_219_297#_M1013_g N_X_c_376_n 0.0164745f $X=3.54 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_219_297#_c_193_n N_X_c_373_n 0.0115011f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_219_297#_c_268_p N_X_c_373_n 3.05012e-19 $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_219_297#_M1001_g N_X_c_401_n 0.0109414f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_219_297#_c_203_n N_X_c_401_n 0.00254059f $X=2.49 $Y=1.53 $X2=0 $Y2=0
cc_195 N_A_219_297#_c_268_p N_X_c_401_n 0.00373137f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_219_297#_M1001_g N_X_c_377_n 0.00153039f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_219_297#_M1011_g N_X_c_377_n 0.0184398f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_198 N_A_219_297#_c_203_n N_X_c_377_n 0.00893203f $X=2.49 $Y=1.53 $X2=0 $Y2=0
cc_199 N_A_219_297#_c_268_p N_X_c_377_n 0.0454006f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_219_297#_c_196_n N_X_c_377_n 0.00449618f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_219_297#_c_192_n N_X_c_374_n 0.00110455f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_219_297#_c_193_n N_X_c_374_n 0.00110455f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_219_297#_c_268_p N_X_c_374_n 0.026132f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A_219_297#_c_196_n N_X_c_374_n 0.00229943f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_219_297#_c_193_n X 0.0223624f $X=3.54 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_219_297#_c_268_p X 0.0142614f $X=3.335 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_219_297#_c_190_n N_VGND_c_444_n 0.00172493f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_219_297#_c_215_n N_VGND_c_444_n 0.034858f $X=1.58 $Y=0.4 $X2=0 $Y2=0
cc_209 N_A_219_297#_c_191_n N_VGND_c_445_n 0.00146448f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_219_297#_c_192_n N_VGND_c_445_n 0.00146448f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_219_297#_c_193_n N_VGND_c_446_n 0.00316354f $X=3.54 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_219_297#_c_190_n N_VGND_c_447_n 0.00542757f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_219_297#_c_191_n N_VGND_c_447_n 0.00425814f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_219_297#_c_192_n N_VGND_c_449_n 0.00425814f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_219_297#_c_193_n N_VGND_c_449_n 0.00425814f $X=3.54 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_219_297#_c_215_n N_VGND_c_451_n 0.0142632f $X=1.58 $Y=0.4 $X2=0 $Y2=0
cc_217 N_A_219_297#_c_195_n N_VGND_c_451_n 0.00176441f $X=1.517 $Y=0.905 $X2=0
+ $Y2=0
cc_218 N_A_219_297#_M1012_d N_VGND_c_453_n 0.00218509f $X=1.445 $Y=0.235 $X2=0
+ $Y2=0
cc_219 N_A_219_297#_c_190_n N_VGND_c_453_n 0.00969354f $X=2.28 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_219_297#_c_191_n N_VGND_c_453_n 0.00573829f $X=2.7 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_219_297#_c_192_n N_VGND_c_453_n 0.00573829f $X=3.12 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_219_297#_c_193_n N_VGND_c_453_n 0.00679592f $X=3.54 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_219_297#_c_215_n N_VGND_c_453_n 0.0118614f $X=1.58 $Y=0.4 $X2=0 $Y2=0
cc_224 N_A_219_297#_c_195_n N_VGND_c_453_n 0.00281074f $X=1.517 $Y=0.905 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_313_n A_301_297# 0.00897657f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_226 N_VPWR_c_313_n N_X_M1000_d 0.00254126f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_313_n N_X_M1011_d 0.00251211f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_320_n N_X_c_417_n 0.0142343f $X=2.785 $Y=2.72 $X2=0 $Y2=0
cc_229 N_VPWR_c_313_n N_X_c_417_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_323_n N_X_c_419_n 0.0140073f $X=3.625 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_313_n N_X_c_419_n 0.00948039f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_232 N_VPWR_c_313_n N_X_c_401_n 0.00600321f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_233 N_VPWR_M1001_s N_X_c_377_n 0.00188877f $X=2.775 $Y=1.485 $X2=0 $Y2=0
cc_234 N_VPWR_c_317_n N_X_c_377_n 0.0126427f $X=2.91 $Y=2.3 $X2=0 $Y2=0
cc_235 N_VPWR_c_313_n N_X_c_377_n 0.00572969f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_M1013_s X 0.00474164f $X=3.615 $Y=1.485 $X2=0 $Y2=0
cc_237 N_VPWR_c_319_n X 0.0174458f $X=3.75 $Y=1.96 $X2=0 $Y2=0
cc_238 N_X_c_371_n N_VGND_M1004_s 0.00167709f $X=3.165 $Y=0.82 $X2=0 $Y2=0
cc_239 N_X_c_373_n N_VGND_M1009_s 0.00529783f $X=3.67 $Y=0.82 $X2=0 $Y2=0
cc_240 N_X_c_372_n N_VGND_c_444_n 0.00788212f $X=2.655 $Y=0.82 $X2=0 $Y2=0
cc_241 N_X_c_371_n N_VGND_c_445_n 0.0113791f $X=3.165 $Y=0.82 $X2=0 $Y2=0
cc_242 N_X_c_373_n N_VGND_c_446_n 0.0130412f $X=3.67 $Y=0.82 $X2=0 $Y2=0
cc_243 N_X_c_380_n N_VGND_c_447_n 0.0153831f $X=2.49 $Y=0.4 $X2=0 $Y2=0
cc_244 N_X_c_371_n N_VGND_c_447_n 0.00193763f $X=3.165 $Y=0.82 $X2=0 $Y2=0
cc_245 N_X_c_371_n N_VGND_c_449_n 0.00193763f $X=3.165 $Y=0.82 $X2=0 $Y2=0
cc_246 N_X_c_395_n N_VGND_c_449_n 0.0153831f $X=3.33 $Y=0.4 $X2=0 $Y2=0
cc_247 N_X_c_373_n N_VGND_c_449_n 0.00193763f $X=3.67 $Y=0.82 $X2=0 $Y2=0
cc_248 N_X_c_373_n N_VGND_c_452_n 0.00356336f $X=3.67 $Y=0.82 $X2=0 $Y2=0
cc_249 N_X_M1003_d N_VGND_c_453_n 0.00217091f $X=2.355 $Y=0.235 $X2=0 $Y2=0
cc_250 N_X_M1006_d N_VGND_c_453_n 0.00217091f $X=3.195 $Y=0.235 $X2=0 $Y2=0
cc_251 N_X_c_380_n N_VGND_c_453_n 0.0119657f $X=2.49 $Y=0.4 $X2=0 $Y2=0
cc_252 N_X_c_371_n N_VGND_c_453_n 0.00828048f $X=3.165 $Y=0.82 $X2=0 $Y2=0
cc_253 N_X_c_395_n N_VGND_c_453_n 0.0119657f $X=3.33 $Y=0.4 $X2=0 $Y2=0
cc_254 N_X_c_373_n N_VGND_c_453_n 0.0107276f $X=3.67 $Y=0.82 $X2=0 $Y2=0

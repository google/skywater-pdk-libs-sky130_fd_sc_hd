* File: sky130_fd_sc_hd__buf_4.pxi.spice
* Created: Tue Sep  1 18:59:17 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_4%A N_A_M1009_g N_A_M1005_g A N_A_c_56_n
+ PM_SKY130_FD_SC_HD__BUF_4%A
x_PM_SKY130_FD_SC_HD__BUF_4%A_27_47# N_A_27_47#_M1009_s N_A_27_47#_M1005_s
+ N_A_27_47#_M1002_g N_A_27_47#_M1000_g N_A_27_47#_M1003_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1004_g N_A_27_47#_M1006_g N_A_27_47#_M1007_g N_A_27_47#_M1008_g
+ N_A_27_47#_c_103_n N_A_27_47#_c_104_n N_A_27_47#_c_178_p N_A_27_47#_c_93_n
+ N_A_27_47#_c_94_n N_A_27_47#_c_117_n N_A_27_47#_c_95_n N_A_27_47#_c_96_n
+ N_A_27_47#_c_129_p N_A_27_47#_c_97_n N_A_27_47#_c_98_n
+ PM_SKY130_FD_SC_HD__BUF_4%A_27_47#
x_PM_SKY130_FD_SC_HD__BUF_4%VPWR N_VPWR_M1005_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_c_192_n N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_196_n
+ N_VPWR_c_197_n VPWR VPWR N_VPWR_c_198_n N_VPWR_c_199_n N_VPWR_c_200_n
+ N_VPWR_c_191_n PM_SKY130_FD_SC_HD__BUF_4%VPWR
x_PM_SKY130_FD_SC_HD__BUF_4%X N_X_M1002_d N_X_M1004_d N_X_M1000_s N_X_M1006_s
+ N_X_c_272_p N_X_c_264_n N_X_c_274_p N_X_c_266_n N_X_c_237_n N_X_c_239_n X X X
+ PM_SKY130_FD_SC_HD__BUF_4%X
x_PM_SKY130_FD_SC_HD__BUF_4%VGND N_VGND_M1009_d N_VGND_M1003_s N_VGND_M1007_s
+ N_VGND_c_281_n N_VGND_c_282_n N_VGND_c_283_n N_VGND_c_284_n N_VGND_c_285_n
+ N_VGND_c_286_n N_VGND_c_287_n N_VGND_c_288_n VGND VGND N_VGND_c_289_n
+ N_VGND_c_290_n PM_SKY130_FD_SC_HD__BUF_4%VGND
cc_1 VNB N_A_M1009_g 0.0230742f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB A 0.0104808f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_56_n 0.0345057f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_M1002_g 0.017747f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1000_g 4.62589e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_6 VNB N_A_27_47#_M1003_g 0.017008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1001_g 4.475e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1004_g 0.0160467f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1006_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1007_g 0.0233974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1008_g 7.17862e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_93_n 0.00173547f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_94_n 0.00183103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_95_n 0.00306151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_96_n 8.76075e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_97_n 9.9617e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_98_n 0.0737477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_191_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_237_n 0.00156003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.00519118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_281_n 0.00174207f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_22 VNB N_VGND_c_282_n 3.15634e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_283_n 0.0148018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_284_n 0.0317254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_285_n 0.0155583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_286_n 0.00340577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_287_n 0.0152957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_288_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_289_n 0.0118624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_290_n 0.168512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VPB N_A_M1005_g 0.0276674f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB A 0.0032877f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_c_56_n 0.00729225f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_34 VPB N_A_27_47#_M1000_g 0.0196327f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_35 VPB N_A_27_47#_M1001_g 0.018902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_47#_M1006_g 0.0177541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_M1008_g 0.0266676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_103_n 0.0088614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_104_n 0.0316012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_96_n 0.00329784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_192_n 0.00222383f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.16
cc_42 VPB N_VPWR_c_193_n 3.03604e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_194_n 0.0147759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_195_n 0.0452743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_196_n 0.0128097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_197_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_198_n 0.0178658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_199_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_200_n 0.00340355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_191_n 0.0493063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_X_c_239_n 0.00181325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB X 0.00293419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB X 0.00269983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 N_A_M1009_g N_A_27_47#_M1002_g 0.0241205f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_55 N_A_c_56_n N_A_27_47#_M1000_g 0.0270159f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_M1005_g N_A_27_47#_c_103_n 8.84614e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_57 A N_A_27_47#_c_103_n 0.0252277f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_56_n N_A_27_47#_c_103_n 0.00179954f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_A_27_47#_c_104_n 0.0101539f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_60 N_A_M1009_g N_A_27_47#_c_93_n 0.0133263f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_61 A N_A_27_47#_c_93_n 0.00885242f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_62 N_A_c_56_n N_A_27_47#_c_93_n 0.00116945f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_63 A N_A_27_47#_c_94_n 0.0139772f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_c_56_n N_A_27_47#_c_94_n 0.00413894f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1005_g N_A_27_47#_c_117_n 0.0113208f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_66 A N_A_27_47#_c_117_n 0.00309924f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_M1009_g N_A_27_47#_c_95_n 0.00384839f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_68 A N_A_27_47#_c_96_n 0.00519104f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_c_56_n N_A_27_47#_c_96_n 0.00432163f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_70 A N_A_27_47#_c_97_n 0.0141041f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_A_27_47#_c_97_n 0.00136438f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_56_n N_A_27_47#_c_98_n 0.01253f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_VPWR_c_192_n 0.00278456f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_VPWR_c_198_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_M1005_g N_VPWR_c_191_n 0.0104829f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_76 N_A_M1009_g N_VGND_c_281_n 0.008483f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_77 N_A_M1009_g N_VGND_c_285_n 0.00379842f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_78 N_A_M1009_g N_VGND_c_290_n 0.00547837f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_117_n N_VPWR_M1005_d 0.00272877f $X=0.64 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_47#_M1000_g N_VPWR_c_192_n 0.010223f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_27_47#_M1001_g N_VPWR_c_192_n 6.64064e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_117_n N_VPWR_c_192_n 0.0131184f $X=0.64 $Y=1.57 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_129_p N_VPWR_c_192_n 5.49869e-19 $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_47#_M1000_g N_VPWR_c_193_n 6.76314e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_27_47#_M1001_g N_VPWR_c_193_n 0.0111118f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_27_47#_M1006_g N_VPWR_c_193_n 0.0110866f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_27_47#_M1008_g N_VPWR_c_193_n 6.72101e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_98_n N_VPWR_c_193_n 2.63087e-19 $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1006_g N_VPWR_c_195_n 8.09353e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1008_g N_VPWR_c_195_n 0.0161847f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1000_g N_VPWR_c_196_n 0.00505556f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_27_47#_M1001_g N_VPWR_c_196_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_104_n N_VPWR_c_198_n 0.0210382f $X=0.26 $Y=2.31 $X2=0 $Y2=0
cc_94 N_A_27_47#_M1006_g N_VPWR_c_199_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_27_47#_M1008_g N_VPWR_c_199_n 0.0046653f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_27_47#_M1005_s N_VPWR_c_191_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_M1000_g N_VPWR_c_191_n 0.00858194f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1001_g N_VPWR_c_191_n 0.00796766f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1006_g N_VPWR_c_191_n 0.00796766f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_27_47#_M1008_g N_VPWR_c_191_n 0.00796766f $X=2.15 $Y=1.985 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_104_n N_VPWR_c_191_n 0.0124268f $X=0.26 $Y=2.31 $X2=0 $Y2=0
cc_102 N_A_27_47#_M1002_g N_X_c_237_n 7.06573e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_93_n N_X_c_237_n 0.00154915f $X=0.64 $Y=0.82 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_129_p N_X_c_237_n 0.0100467f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_98_n N_X_c_237_n 0.00216279f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1000_g N_X_c_239_n 6.55102e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_96_n N_X_c_239_n 0.00288331f $X=0.725 $Y=1.485 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_129_p N_X_c_239_n 0.00893131f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_98_n N_X_c_239_n 0.00213561f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_27_47#_M1003_g X 0.0158916f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1001_g X 0.00389939f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1004_g X 0.0125487f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1006_g X 0.00434593f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_27_47#_M1007_g X 0.00463984f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A_27_47#_M1008_g X 0.00437841f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_129_p X 0.00689751f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_98_n X 0.0406104f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1001_g X 0.0147808f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1006_g X 0.0120253f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1008_g X 0.0015501f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_98_n X 0.00142331f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_93_n N_VGND_M1009_d 0.00193386f $X=0.64 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_27_47#_M1002_g N_VGND_c_281_n 0.00141404f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_93_n N_VGND_c_281_n 0.0145326f $X=0.64 $Y=0.82 $X2=0 $Y2=0
cc_125 N_A_27_47#_M1002_g N_VGND_c_282_n 6.10735e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_126 N_A_27_47#_M1003_g N_VGND_c_282_n 0.00787546f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1004_g N_VGND_c_282_n 0.00768883f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1007_g N_VGND_c_282_n 5.77787e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_98_n N_VGND_c_282_n 2.53763e-19 $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1004_g N_VGND_c_284_n 7.31324e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1007_g N_VGND_c_284_n 0.0125339f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_178_p N_VGND_c_285_n 0.0115672f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_93_n N_VGND_c_285_n 0.00206869f $X=0.64 $Y=0.82 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1002_g N_VGND_c_287_n 0.00585385f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_135 N_A_27_47#_M1003_g N_VGND_c_287_n 0.00350562f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1004_g N_VGND_c_289_n 0.00350455f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1007_g N_VGND_c_289_n 0.0046653f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_138 N_A_27_47#_M1009_s N_VGND_c_290_n 0.00377256f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_M1002_g N_VGND_c_290_n 0.0106402f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_27_47#_M1003_g N_VGND_c_290_n 0.00418574f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_27_47#_M1004_g N_VGND_c_290_n 0.00418373f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A_27_47#_M1007_g N_VGND_c_290_n 0.00796766f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_178_p N_VGND_c_290_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_93_n N_VGND_c_290_n 0.00629255f $X=0.64 $Y=0.82 $X2=0 $Y2=0
cc_145 N_VPWR_c_191_n N_X_M1000_s 0.00570907f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_146 N_VPWR_c_191_n N_X_M1006_s 0.00570907f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_147 N_VPWR_c_196_n N_X_c_264_n 0.0113958f $X=1.355 $Y=2.72 $X2=0 $Y2=0
cc_148 N_VPWR_c_191_n N_X_c_264_n 0.00646998f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_149 N_VPWR_c_199_n N_X_c_266_n 0.0113958f $X=2.195 $Y=2.72 $X2=0 $Y2=0
cc_150 N_VPWR_c_191_n N_X_c_266_n 0.00646998f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_151 N_VPWR_M1001_d X 0.00187831f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_152 N_VPWR_c_193_n X 0.0146577f $X=1.52 $Y=2 $X2=0 $Y2=0
cc_153 N_VPWR_c_195_n N_VGND_c_284_n 0.00942828f $X=2.36 $Y=1.66 $X2=0 $Y2=0
cc_154 X N_VGND_M1003_s 0.00163861f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_155 X N_VGND_c_282_n 0.0171742f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_156 N_X_c_272_p N_VGND_c_287_n 0.0113595f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_157 X N_VGND_c_287_n 0.00193763f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_158 N_X_c_274_p N_VGND_c_289_n 0.0113958f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_159 X N_VGND_c_289_n 0.00209862f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_160 N_X_M1002_d N_VGND_c_290_n 0.00418657f $X=0.965 $Y=0.235 $X2=0 $Y2=0
cc_161 N_X_M1004_d N_VGND_c_290_n 0.00418582f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_162 N_X_c_272_p N_VGND_c_290_n 0.0064623f $X=1.1 $Y=0.56 $X2=0 $Y2=0
cc_163 N_X_c_274_p N_VGND_c_290_n 0.00646998f $X=1.94 $Y=0.56 $X2=0 $Y2=0
cc_164 X N_VGND_c_290_n 0.00931472f $X=1.53 $Y=0.765 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a21boi_0.pxi.spice
* Created: Thu Aug 27 14:00:23 2020
* 
x_PM_SKY130_FD_SC_HD__A21BOI_0%B1_N N_B1_N_M1003_g N_B1_N_c_61_n N_B1_N_M1002_g
+ N_B1_N_c_63_n B1_N N_B1_N_c_59_n N_B1_N_c_60_n
+ PM_SKY130_FD_SC_HD__A21BOI_0%B1_N
x_PM_SKY130_FD_SC_HD__A21BOI_0%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_93_n N_A_27_47#_c_94_n N_A_27_47#_c_95_n N_A_27_47#_M1006_g
+ N_A_27_47#_M1004_g N_A_27_47#_c_102_n N_A_27_47#_c_96_n N_A_27_47#_c_97_n
+ N_A_27_47#_c_98_n N_A_27_47#_c_103_n N_A_27_47#_c_99_n
+ PM_SKY130_FD_SC_HD__A21BOI_0%A_27_47#
x_PM_SKY130_FD_SC_HD__A21BOI_0%A1 N_A1_M1001_g N_A1_M1007_g N_A1_c_152_n
+ N_A1_c_153_n N_A1_c_154_n A1 N_A1_c_155_n N_A1_c_156_n
+ PM_SKY130_FD_SC_HD__A21BOI_0%A1
x_PM_SKY130_FD_SC_HD__A21BOI_0%A2 N_A2_M1000_g N_A2_c_196_n N_A2_M1005_g
+ N_A2_c_197_n A2 N_A2_c_199_n N_A2_c_200_n PM_SKY130_FD_SC_HD__A21BOI_0%A2
x_PM_SKY130_FD_SC_HD__A21BOI_0%VPWR N_VPWR_M1002_d N_VPWR_M1001_d N_VPWR_c_227_n
+ N_VPWR_c_228_n VPWR N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n
+ N_VPWR_c_226_n N_VPWR_c_233_n N_VPWR_c_234_n PM_SKY130_FD_SC_HD__A21BOI_0%VPWR
x_PM_SKY130_FD_SC_HD__A21BOI_0%Y N_Y_M1006_d N_Y_M1004_s N_Y_c_268_n N_Y_c_269_n
+ Y PM_SKY130_FD_SC_HD__A21BOI_0%Y
x_PM_SKY130_FD_SC_HD__A21BOI_0%A_300_369# N_A_300_369#_M1004_d
+ N_A_300_369#_M1005_d N_A_300_369#_c_301_n N_A_300_369#_c_302_n
+ N_A_300_369#_c_303_n PM_SKY130_FD_SC_HD__A21BOI_0%A_300_369#
x_PM_SKY130_FD_SC_HD__A21BOI_0%VGND N_VGND_M1003_d N_VGND_M1000_d N_VGND_c_330_n
+ N_VGND_c_331_n VGND N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n
+ PM_SKY130_FD_SC_HD__A21BOI_0%VGND
cc_1 VNB N_B1_N_M1003_g 0.0514486f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_B1_N_c_59_n 0.00860684f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.4
cc_3 VNB N_B1_N_c_60_n 0.00357717f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.4
cc_4 VNB N_A_27_47#_c_93_n 0.0513882f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.885
cc_5 VNB N_A_27_47#_c_94_n 0.0209875f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_6 VNB N_A_27_47#_c_95_n 0.0205569f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_7 VNB N_A_27_47#_c_96_n 0.0208554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_97_n 0.00808219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_98_n 0.0145959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_99_n 0.0133528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_152_n 0.0114193f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_12 VNB N_A1_c_153_n 0.017814f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_13 VNB N_A1_c_154_n 2.80507e-19 $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.885
cc_14 VNB N_A1_c_155_n 0.0223112f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.4
cc_15 VNB N_A1_c_156_n 0.0077197f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.4
cc_16 VNB N_A2_c_196_n 0.0256553f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.44
cc_17 VNB N_A2_c_197_n 0.00416751f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A2 0.0219075f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.885
cc_19 VNB N_A2_c_199_n 0.0209972f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.4
cc_20 VNB N_A2_c_200_n 0.0207577f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=1.4
cc_21 VNB N_VPWR_c_226_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_268_n 9.34776e-19 $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.885
cc_23 VNB N_Y_c_269_n 0.00408859f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_24 VNB N_VGND_c_330_n 0.0103398f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.885
cc_25 VNB N_VGND_c_331_n 0.0182339f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=2.275
cc_26 VNB N_VGND_c_332_n 0.0356652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_333_n 0.0339017f $X=-0.19 $Y=-0.24 $X2=0.682 $Y2=1.4
cc_28 VNB N_VGND_c_334_n 0.161677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_B1_N_c_61_n 0.0198716f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.71
cc_30 VPB N_B1_N_M1002_g 0.0269148f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.275
cc_31 VPB N_B1_N_c_63_n 0.0202113f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.885
cc_32 VPB N_B1_N_c_59_n 0.00987419f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_33 VPB N_B1_N_c_60_n 0.00786316f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_34 VPB N_A_27_47#_c_94_n 0.0105617f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.275
cc_35 VPB N_A_27_47#_M1004_g 0.0235039f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.4
cc_36 VPB N_A_27_47#_c_102_n 0.0331956f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_37 VPB N_A_27_47#_c_103_n 0.0145863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_99_n 0.0377476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A1_M1001_g 0.0315647f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.445
cc_40 VPB N_A1_c_154_n 0.0108075f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.885
cc_41 VPB N_A1_c_156_n 0.00498526f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_42 VPB N_A2_M1005_g 0.0463711f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.275
cc_43 VPB N_A2_c_197_n 0.0168297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB A2 0.00808647f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.885
cc_45 VPB N_VPWR_c_227_n 0.00621036f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.275
cc_46 VPB N_VPWR_c_228_n 0.00474108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_229_n 0.0153759f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.265
cc_48 VPB N_VPWR_c_230_n 0.0293736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_231_n 0.0171491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_226_n 0.0519058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_233_n 0.00510584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_234_n 0.00362058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_Y_c_268_n 0.00333792f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.885
cc_54 VPB Y 0.00912866f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_55 VPB N_A_300_369#_c_301_n 0.0035954f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=2.275
cc_56 VPB N_A_300_369#_c_302_n 0.00655518f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.4
cc_57 VPB N_A_300_369#_c_303_n 0.0302695f $X=-0.19 $Y=1.305 $X2=0.585 $Y2=1.4
cc_58 N_B1_N_M1003_g N_A_27_47#_c_93_n 0.0133739f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_59 N_B1_N_c_60_n N_A_27_47#_c_93_n 0.00184543f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_60 N_B1_N_M1003_g N_A_27_47#_c_94_n 0.00613729f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_61 N_B1_N_c_59_n N_A_27_47#_c_94_n 0.0100287f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_62 N_B1_N_c_60_n N_A_27_47#_c_94_n 0.00386066f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_63 N_B1_N_M1003_g N_A_27_47#_c_95_n 0.00618331f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_64 N_B1_N_c_61_n N_A_27_47#_M1004_g 0.00247065f $X=0.575 $Y=1.71 $X2=0 $Y2=0
cc_65 N_B1_N_c_61_n N_A_27_47#_c_102_n 0.0100287f $X=0.575 $Y=1.71 $X2=0 $Y2=0
cc_66 N_B1_N_M1003_g N_A_27_47#_c_96_n 0.00561773f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_67 N_B1_N_M1003_g N_A_27_47#_c_97_n 0.0192495f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_68 N_B1_N_c_59_n N_A_27_47#_c_97_n 0.00120624f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_69 N_B1_N_c_60_n N_A_27_47#_c_97_n 0.0357041f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_70 N_B1_N_M1003_g N_A_27_47#_c_99_n 0.0293802f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_71 N_B1_N_c_60_n N_A_27_47#_c_99_n 0.0585201f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_72 N_B1_N_M1002_g N_VPWR_c_227_n 0.0100685f $X=0.475 $Y=2.275 $X2=0 $Y2=0
cc_73 N_B1_N_c_63_n N_VPWR_c_227_n 0.00110929f $X=0.575 $Y=1.885 $X2=0 $Y2=0
cc_74 N_B1_N_c_60_n N_VPWR_c_227_n 0.0211297f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_75 N_B1_N_M1002_g N_VPWR_c_229_n 0.00486043f $X=0.475 $Y=2.275 $X2=0 $Y2=0
cc_76 N_B1_N_M1002_g N_VPWR_c_226_n 0.0074654f $X=0.475 $Y=2.275 $X2=0 $Y2=0
cc_77 N_B1_N_c_60_n N_VPWR_c_226_n 0.00505156f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_78 N_B1_N_c_59_n N_Y_c_268_n 3.48912e-19 $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_79 N_B1_N_c_60_n N_Y_c_268_n 0.0380762f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_80 N_B1_N_c_61_n Y 6.17107e-19 $X=0.575 $Y=1.71 $X2=0 $Y2=0
cc_81 N_B1_N_M1002_g Y 0.00488856f $X=0.475 $Y=2.275 $X2=0 $Y2=0
cc_82 N_B1_N_c_60_n Y 0.0247793f $X=0.585 $Y=1.4 $X2=0 $Y2=0
cc_83 N_B1_N_M1003_g N_VGND_c_332_n 0.00986672f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_84 N_B1_N_M1003_g N_VGND_c_334_n 0.00767637f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_102_n N_A1_M1001_g 0.0243907f $X=1.255 $Y=1.68 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_93_n N_A1_c_152_n 0.0181128f $X=1.255 $Y=1.065 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_95_n N_A1_c_153_n 0.00819422f $X=1.245 $Y=0.77 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_94_n N_A1_c_155_n 0.0181128f $X=1.255 $Y=1.435 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_93_n N_A1_c_156_n 4.015e-19 $X=1.255 $Y=1.065 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_94_n N_A1_c_156_n 4.05015e-19 $X=1.255 $Y=1.435 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1004_g N_VPWR_c_227_n 0.00304341f $X=1.425 $Y=2.165 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_c_103_n N_VPWR_c_229_n 0.0176892f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1004_g N_VPWR_c_230_n 0.0054895f $X=1.425 $Y=2.165 $X2=0 $Y2=0
cc_94 N_A_27_47#_M1002_s N_VPWR_c_226_n 0.00369639f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_M1004_g N_VPWR_c_226_n 0.0113139f $X=1.425 $Y=2.165 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_103_n N_VPWR_c_226_n 0.00990583f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_94_n N_Y_c_268_n 0.0222339f $X=1.255 $Y=1.435 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_102_n N_Y_c_268_n 0.0208697f $X=1.255 $Y=1.68 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_97_n N_Y_c_268_n 0.00602972f $X=0.98 $Y=0.93 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_93_n N_Y_c_269_n 0.0161454f $X=1.255 $Y=1.065 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_94_n N_Y_c_269_n 0.00941342f $X=1.255 $Y=1.435 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_95_n N_Y_c_269_n 0.011696f $X=1.245 $Y=0.77 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_97_n N_Y_c_269_n 0.0197003f $X=0.98 $Y=0.93 $X2=0 $Y2=0
cc_104 N_A_27_47#_M1004_g Y 0.00850081f $X=1.425 $Y=2.165 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_102_n Y 0.00786461f $X=1.255 $Y=1.68 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1004_g N_A_300_369#_c_302_n 0.00758233f $X=1.425 $Y=2.165
+ $X2=0 $Y2=0
cc_107 N_A_27_47#_c_93_n N_VGND_c_332_n 0.00239528f $X=1.255 $Y=1.065 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_95_n N_VGND_c_332_n 0.00381759f $X=1.245 $Y=0.77 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_96_n N_VGND_c_332_n 0.0161283f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_97_n N_VGND_c_332_n 0.0451257f $X=0.98 $Y=0.93 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_93_n N_VGND_c_333_n 3.8293e-19 $X=1.255 $Y=1.065 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_95_n N_VGND_c_333_n 0.00579312f $X=1.245 $Y=0.77 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1003_s N_VGND_c_334_n 0.00226047f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_93_n N_VGND_c_334_n 6.40452e-19 $X=1.255 $Y=1.065 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_95_n N_VGND_c_334_n 0.0116953f $X=1.245 $Y=0.77 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_96_n N_VGND_c_334_n 0.010767f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_97_n N_VGND_c_334_n 0.0073992f $X=0.98 $Y=0.93 $X2=0 $Y2=0
cc_118 N_A1_c_155_n N_A2_c_196_n 0.0206196f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_119 N_A1_M1001_g N_A2_M1005_g 0.0379996f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_120 N_A1_c_154_n N_A2_c_197_n 0.0206196f $X=1.865 $Y=1.435 $X2=0 $Y2=0
cc_121 N_A1_c_152_n A2 5.03093e-19 $X=1.865 $Y=0.9 $X2=0 $Y2=0
cc_122 N_A1_c_156_n A2 0.0529629f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_123 N_A1_c_152_n N_A2_c_199_n 0.0206196f $X=1.865 $Y=0.9 $X2=0 $Y2=0
cc_124 N_A1_c_156_n N_A2_c_199_n 0.0101957f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_125 N_A1_c_153_n N_A2_c_200_n 0.0206196f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_126 N_A1_M1001_g N_VPWR_c_228_n 0.00275982f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_127 N_A1_M1001_g N_VPWR_c_230_n 0.00424868f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_128 N_A1_M1001_g N_VPWR_c_226_n 0.00581442f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_129 N_A1_M1001_g N_Y_c_268_n 0.00212966f $X=1.855 $Y=2.165 $X2=0 $Y2=0
cc_130 N_A1_c_155_n N_Y_c_268_n 0.0015651f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_131 N_A1_c_156_n N_Y_c_268_n 0.0346076f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_132 N_A1_c_152_n N_Y_c_269_n 0.00274346f $X=1.865 $Y=0.9 $X2=0 $Y2=0
cc_133 N_A1_c_153_n N_Y_c_269_n 0.0118895f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_134 N_A1_c_156_n N_Y_c_269_n 0.0345029f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_135 N_A1_M1001_g N_A_300_369#_c_301_n 0.00916243f $X=1.855 $Y=2.165 $X2=0
+ $Y2=0
cc_136 N_A1_c_154_n N_A_300_369#_c_301_n 3.16357e-19 $X=1.865 $Y=1.435 $X2=0
+ $Y2=0
cc_137 N_A1_c_156_n N_A_300_369#_c_301_n 0.0254973f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_138 N_A1_M1001_g N_A_300_369#_c_302_n 0.00707734f $X=1.855 $Y=2.165 $X2=0
+ $Y2=0
cc_139 N_A1_c_154_n N_A_300_369#_c_302_n 0.00187511f $X=1.865 $Y=1.435 $X2=0
+ $Y2=0
cc_140 N_A1_c_156_n N_A_300_369#_c_302_n 0.00170493f $X=1.865 $Y=0.93 $X2=0
+ $Y2=0
cc_141 N_A1_M1001_g N_A_300_369#_c_303_n 5.16893e-19 $X=1.855 $Y=2.165 $X2=0
+ $Y2=0
cc_142 N_A1_c_153_n N_VGND_c_331_n 0.00292002f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_143 N_A1_c_152_n N_VGND_c_333_n 0.00149925f $X=1.865 $Y=0.9 $X2=0 $Y2=0
cc_144 N_A1_c_153_n N_VGND_c_333_n 0.00585385f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_145 N_A1_c_152_n N_VGND_c_334_n 0.00133936f $X=1.865 $Y=0.9 $X2=0 $Y2=0
cc_146 N_A1_c_153_n N_VGND_c_334_n 0.00662154f $X=1.865 $Y=0.765 $X2=0 $Y2=0
cc_147 N_A1_c_156_n N_VGND_c_334_n 0.0148028f $X=1.865 $Y=0.93 $X2=0 $Y2=0
cc_148 N_A2_M1005_g N_VPWR_c_228_n 0.00275982f $X=2.285 $Y=2.165 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_VPWR_c_231_n 0.00424868f $X=2.285 $Y=2.165 $X2=0 $Y2=0
cc_150 N_A2_M1005_g N_VPWR_c_226_n 0.00672169f $X=2.285 $Y=2.165 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_A_300_369#_c_301_n 0.0127871f $X=2.285 $Y=2.165 $X2=0
+ $Y2=0
cc_152 N_A2_M1005_g N_A_300_369#_c_302_n 5.16893e-19 $X=2.285 $Y=2.165 $X2=0
+ $Y2=0
cc_153 N_A2_M1005_g N_A_300_369#_c_303_n 0.00756041f $X=2.285 $Y=2.165 $X2=0
+ $Y2=0
cc_154 N_A2_c_197_n N_A_300_369#_c_303_n 0.00145273f $X=2.39 $Y=1.435 $X2=0
+ $Y2=0
cc_155 A2 N_A_300_369#_c_303_n 0.0130978f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_156 A2 N_VGND_c_331_n 0.0206335f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_157 N_A2_c_199_n N_VGND_c_331_n 0.00146533f $X=2.435 $Y=0.93 $X2=0 $Y2=0
cc_158 N_A2_c_200_n N_VGND_c_331_n 0.0126065f $X=2.39 $Y=0.765 $X2=0 $Y2=0
cc_159 N_A2_c_200_n N_VGND_c_333_n 0.00486043f $X=2.39 $Y=0.765 $X2=0 $Y2=0
cc_160 A2 N_VGND_c_334_n 0.00101891f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_161 N_A2_c_200_n N_VGND_c_334_n 0.00814024f $X=2.39 $Y=0.765 $X2=0 $Y2=0
cc_162 N_VPWR_c_226_n N_Y_M1004_s 0.00373913f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_227_n Y 0.0203341f $X=0.69 $Y=2.3 $X2=0 $Y2=0
cc_164 N_VPWR_c_230_n Y 0.0163792f $X=1.975 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_c_226_n Y 0.0091658f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_226_n N_A_300_369#_M1004_d 0.00223231f $X=2.53 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_167 N_VPWR_c_226_n N_A_300_369#_M1005_d 0.00213418f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_VPWR_M1001_d N_A_300_369#_c_301_n 0.00172254f $X=1.93 $Y=1.845 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_228_n N_A_300_369#_c_301_n 0.0130079f $X=2.07 $Y=2.34 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_230_n N_A_300_369#_c_301_n 0.0020606f $X=1.975 $Y=2.72 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_231_n N_A_300_369#_c_301_n 0.0020606f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_226_n N_A_300_369#_c_301_n 0.00846507f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_230_n N_A_300_369#_c_302_n 0.0188597f $X=1.975 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_226_n N_A_300_369#_c_302_n 0.0122476f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_231_n N_A_300_369#_c_303_n 0.0209643f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_226_n N_A_300_369#_c_303_n 0.0124297f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_177 N_Y_c_268_n N_A_300_369#_c_302_n 0.0119468f $X=1.462 $Y=1.2 $X2=0 $Y2=0
cc_178 Y N_A_300_369#_c_302_n 0.00833879f $X=1.065 $Y=2.125 $X2=0 $Y2=0
cc_179 N_Y_c_269_n N_VGND_c_333_n 0.0185768f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_180 N_Y_M1006_d N_VGND_c_334_n 0.00946742f $X=1.32 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_c_269_n N_VGND_c_334_n 0.0112558f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_182 N_VGND_c_334_n A_400_47# 0.00404825f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__sdfbbp_1.pxi.spice
* Created: Tue Sep  1 19:29:44 2020
* 
x_PM_SKY130_FD_SC_HD__SDFBBP_1%CLK N_CLK_c_305_n N_CLK_c_300_n N_CLK_M1045_g
+ N_CLK_c_306_n N_CLK_M1026_g N_CLK_c_301_n N_CLK_c_307_n CLK CLK N_CLK_c_303_n
+ N_CLK_c_304_n PM_SKY130_FD_SC_HD__SDFBBP_1%CLK
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_27_47# N_A_27_47#_M1045_s N_A_27_47#_M1026_s
+ N_A_27_47#_M1027_g N_A_27_47#_M1000_g N_A_27_47#_c_345_n N_A_27_47#_M1043_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1033_g N_A_27_47#_c_346_n N_A_27_47#_c_347_n
+ N_A_27_47#_M1025_g N_A_27_47#_c_598_p N_A_27_47#_c_349_n N_A_27_47#_c_350_n
+ N_A_27_47#_c_360_n N_A_27_47#_c_476_p N_A_27_47#_c_351_n N_A_27_47#_c_352_n
+ N_A_27_47#_c_353_n N_A_27_47#_c_363_n N_A_27_47#_c_364_n N_A_27_47#_c_365_n
+ N_A_27_47#_c_366_n N_A_27_47#_c_367_n N_A_27_47#_c_368_n N_A_27_47#_c_354_n
+ N_A_27_47#_c_370_n N_A_27_47#_c_371_n N_A_27_47#_c_372_n N_A_27_47#_c_373_n
+ N_A_27_47#_c_374_n PM_SKY130_FD_SC_HD__SDFBBP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%SCD N_SCD_M1007_g N_SCD_M1034_g SCD SCD
+ N_SCD_c_613_n PM_SKY130_FD_SC_HD__SDFBBP_1%SCD
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_423_315# N_A_423_315#_M1012_s
+ N_A_423_315#_M1035_s N_A_423_315#_c_652_n N_A_423_315#_M1040_g
+ N_A_423_315#_c_653_n N_A_423_315#_c_654_n N_A_423_315#_M1020_g
+ N_A_423_315#_c_655_n N_A_423_315#_c_707_p N_A_423_315#_c_656_n
+ N_A_423_315#_c_645_n N_A_423_315#_c_646_n N_A_423_315#_c_647_n
+ N_A_423_315#_c_648_n N_A_423_315#_c_649_n N_A_423_315#_c_658_n
+ N_A_423_315#_c_650_n N_A_423_315#_c_651_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_423_315#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%SCE N_SCE_c_749_n N_SCE_M1022_g N_SCE_c_750_n
+ N_SCE_c_751_n N_SCE_M1012_g N_SCE_c_752_n N_SCE_c_759_n N_SCE_M1035_g
+ N_SCE_c_760_n N_SCE_c_761_n N_SCE_M1019_g N_SCE_c_753_n N_SCE_c_762_n
+ N_SCE_c_754_n SCE SCE SCE N_SCE_c_757_n PM_SKY130_FD_SC_HD__SDFBBP_1%SCE
x_PM_SKY130_FD_SC_HD__SDFBBP_1%D N_D_M1023_g N_D_M1014_g D D N_D_c_851_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%D
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_193_47# N_A_193_47#_M1027_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1041_g N_A_193_47#_c_889_n N_A_193_47#_c_890_n
+ N_A_193_47#_M1015_g N_A_193_47#_c_892_n N_A_193_47#_c_893_n
+ N_A_193_47#_M1009_g N_A_193_47#_M1017_g N_A_193_47#_c_894_n
+ N_A_193_47#_c_895_n N_A_193_47#_c_896_n N_A_193_47#_c_911_n
+ N_A_193_47#_c_912_n N_A_193_47#_c_897_n N_A_193_47#_c_898_n
+ N_A_193_47#_c_899_n N_A_193_47#_c_900_n N_A_193_47#_c_901_n
+ N_A_193_47#_c_902_n N_A_193_47#_c_903_n N_A_193_47#_c_904_n
+ N_A_193_47#_c_905_n N_A_193_47#_c_906_n PM_SKY130_FD_SC_HD__SDFBBP_1%A_193_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_1107_21# N_A_1107_21#_M1029_d
+ N_A_1107_21#_M1011_d N_A_1107_21#_M1038_g N_A_1107_21#_M1036_g
+ N_A_1107_21#_M1047_g N_A_1107_21#_c_1121_n N_A_1107_21#_M1003_g
+ N_A_1107_21#_c_1130_n N_A_1107_21#_c_1179_p N_A_1107_21#_c_1143_n
+ N_A_1107_21#_c_1122_n N_A_1107_21#_c_1123_n N_A_1107_21#_c_1124_n
+ N_A_1107_21#_c_1132_n N_A_1107_21#_c_1133_n N_A_1107_21#_c_1148_n
+ N_A_1107_21#_c_1125_n N_A_1107_21#_c_1126_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_1107_21#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%SET_B N_SET_B_c_1266_n N_SET_B_M1011_g
+ N_SET_B_M1044_g N_SET_B_M1004_g N_SET_B_M1008_g SET_B N_SET_B_c_1272_n
+ N_SET_B_c_1273_n N_SET_B_c_1274_n N_SET_B_c_1275_n N_SET_B_c_1276_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%SET_B
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_931_47# N_A_931_47#_M1043_d N_A_931_47#_M1041_d
+ N_A_931_47#_M1029_g N_A_931_47#_M1037_g N_A_931_47#_c_1405_n
+ N_A_931_47#_c_1411_n N_A_931_47#_c_1401_n N_A_931_47#_c_1396_n
+ N_A_931_47#_c_1397_n N_A_931_47#_c_1398_n N_A_931_47#_c_1399_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_931_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_1400_21# N_A_1400_21#_M1013_s
+ N_A_1400_21#_M1006_s N_A_1400_21#_c_1500_n N_A_1400_21#_M1028_g
+ N_A_1400_21#_c_1501_n N_A_1400_21#_M1032_g N_A_1400_21#_M1030_g
+ N_A_1400_21#_M1031_g N_A_1400_21#_c_1503_n N_A_1400_21#_c_1504_n
+ N_A_1400_21#_c_1512_n N_A_1400_21#_c_1513_n N_A_1400_21#_c_1505_n
+ N_A_1400_21#_c_1506_n N_A_1400_21#_c_1515_n N_A_1400_21#_c_1516_n
+ N_A_1400_21#_c_1517_n N_A_1400_21#_c_1518_n N_A_1400_21#_c_1507_n
+ N_A_1400_21#_c_1508_n PM_SKY130_FD_SC_HD__SDFBBP_1%A_1400_21#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_1887_21# N_A_1887_21#_M1018_d
+ N_A_1887_21#_M1008_d N_A_1887_21#_M1005_g N_A_1887_21#_M1042_g
+ N_A_1887_21#_c_1659_n N_A_1887_21#_M1001_g N_A_1887_21#_M1039_g
+ N_A_1887_21#_c_1660_n N_A_1887_21#_c_1661_n N_A_1887_21#_c_1662_n
+ N_A_1887_21#_c_1663_n N_A_1887_21#_c_1664_n N_A_1887_21#_M1046_g
+ N_A_1887_21#_c_1674_n N_A_1887_21#_M1021_g N_A_1887_21#_c_1665_n
+ N_A_1887_21#_c_1666_n N_A_1887_21#_c_1675_n N_A_1887_21#_c_1676_n
+ N_A_1887_21#_c_1677_n N_A_1887_21#_c_1678_n N_A_1887_21#_c_1735_p
+ N_A_1887_21#_c_1783_p N_A_1887_21#_c_1706_n N_A_1887_21#_c_1667_n
+ N_A_1887_21#_c_1680_n N_A_1887_21#_c_1681_n N_A_1887_21#_c_1723_n
+ N_A_1887_21#_c_1699_n N_A_1887_21#_c_1726_n N_A_1887_21#_c_1668_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_1887_21#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_1714_47# N_A_1714_47#_M1009_d
+ N_A_1714_47#_M1033_d N_A_1714_47#_M1018_g N_A_1714_47#_M1024_g
+ N_A_1714_47#_c_1852_n N_A_1714_47#_c_1855_n N_A_1714_47#_c_1841_n
+ N_A_1714_47#_c_1847_n N_A_1714_47#_c_1842_n N_A_1714_47#_c_1843_n
+ N_A_1714_47#_c_1844_n N_A_1714_47#_c_1845_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_1714_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%RESET_B N_RESET_B_M1013_g N_RESET_B_M1006_g
+ RESET_B N_RESET_B_c_1940_n PM_SKY130_FD_SC_HD__SDFBBP_1%RESET_B
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_2596_47# N_A_2596_47#_M1046_s
+ N_A_2596_47#_M1021_s N_A_2596_47#_M1016_g N_A_2596_47#_M1002_g
+ N_A_2596_47#_c_1974_n N_A_2596_47#_c_1980_n N_A_2596_47#_c_1975_n
+ N_A_2596_47#_c_1976_n N_A_2596_47#_c_1977_n N_A_2596_47#_c_1978_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_2596_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%VPWR N_VPWR_M1026_d N_VPWR_M1034_s N_VPWR_M1035_d
+ N_VPWR_M1036_d N_VPWR_M1032_d N_VPWR_M1042_d N_VPWR_M1030_d N_VPWR_M1006_d
+ N_VPWR_M1021_d N_VPWR_c_2027_n N_VPWR_c_2028_n N_VPWR_c_2029_n N_VPWR_c_2030_n
+ N_VPWR_c_2031_n N_VPWR_c_2032_n N_VPWR_c_2033_n N_VPWR_c_2034_n
+ N_VPWR_c_2035_n N_VPWR_c_2036_n VPWR VPWR N_VPWR_c_2037_n N_VPWR_c_2038_n
+ N_VPWR_c_2039_n N_VPWR_c_2040_n N_VPWR_c_2041_n N_VPWR_c_2042_n
+ N_VPWR_c_2043_n N_VPWR_c_2044_n N_VPWR_c_2026_n N_VPWR_c_2046_n
+ N_VPWR_c_2047_n N_VPWR_c_2048_n N_VPWR_c_2049_n N_VPWR_c_2050_n
+ N_VPWR_c_2051_n N_VPWR_c_2052_n PM_SKY130_FD_SC_HD__SDFBBP_1%VPWR
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_453_363# N_A_453_363#_M1022_d
+ N_A_453_363#_M1023_d N_A_453_363#_M1040_d N_A_453_363#_M1014_d
+ N_A_453_363#_c_2238_n N_A_453_363#_c_2246_n N_A_453_363#_c_2247_n
+ N_A_453_363#_c_2239_n N_A_453_363#_c_2240_n N_A_453_363#_c_2241_n
+ N_A_453_363#_c_2242_n N_A_453_363#_c_2243_n N_A_453_363#_c_2244_n
+ N_A_453_363#_c_2245_n PM_SKY130_FD_SC_HD__SDFBBP_1%A_453_363#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%Q_N N_Q_N_M1001_d N_Q_N_M1039_d N_Q_N_c_2374_n
+ N_Q_N_c_2371_n Q_N Q_N Q_N N_Q_N_c_2373_n Q_N PM_SKY130_FD_SC_HD__SDFBBP_1%Q_N
x_PM_SKY130_FD_SC_HD__SDFBBP_1%Q N_Q_M1016_d N_Q_M1002_d N_Q_c_2402_n
+ N_Q_c_2405_n N_Q_c_2403_n Q Q Q PM_SKY130_FD_SC_HD__SDFBBP_1%Q
x_PM_SKY130_FD_SC_HD__SDFBBP_1%VGND N_VGND_M1045_d N_VGND_M1007_s N_VGND_M1012_d
+ N_VGND_M1038_d N_VGND_M1003_s N_VGND_M1005_d N_VGND_M1013_d N_VGND_M1046_d
+ N_VGND_c_2418_n N_VGND_c_2419_n N_VGND_c_2420_n N_VGND_c_2421_n
+ N_VGND_c_2422_n N_VGND_c_2423_n N_VGND_c_2424_n N_VGND_c_2425_n
+ N_VGND_c_2426_n N_VGND_c_2427_n N_VGND_c_2428_n N_VGND_c_2429_n
+ N_VGND_c_2430_n N_VGND_c_2431_n VGND VGND N_VGND_c_2432_n N_VGND_c_2433_n
+ N_VGND_c_2434_n N_VGND_c_2435_n N_VGND_c_2436_n N_VGND_c_2437_n
+ N_VGND_c_2438_n N_VGND_c_2439_n N_VGND_c_2440_n N_VGND_c_2441_n
+ N_VGND_c_2442_n N_VGND_c_2443_n PM_SKY130_FD_SC_HD__SDFBBP_1%VGND
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_1251_47# N_A_1251_47#_M1044_d
+ N_A_1251_47#_M1028_d N_A_1251_47#_c_2632_n N_A_1251_47#_c_2635_n
+ N_A_1251_47#_c_2642_n PM_SKY130_FD_SC_HD__SDFBBP_1%A_1251_47#
x_PM_SKY130_FD_SC_HD__SDFBBP_1%A_2026_47# N_A_2026_47#_M1004_d
+ N_A_2026_47#_M1031_d N_A_2026_47#_c_2665_n N_A_2026_47#_c_2662_n
+ PM_SKY130_FD_SC_HD__SDFBBP_1%A_2026_47#
cc_1 VNB N_CLK_c_300_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_CLK_c_301_n 0.0233701f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB CLK 0.0187448f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_303_n 0.0195341f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_c_304_n 0.0141401f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1027_g 0.0365281f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_345_n 0.0180417f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_8 VNB N_A_27_47#_c_346_n 0.0123509f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_9 VNB N_A_27_47#_c_347_n 0.00338667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1025_g 0.0470486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_349_n 0.00157584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_350_n 0.00643757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_351_n 0.00246572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_352_n 0.0042958f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_353_n 0.0326251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_354_n 0.0229605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCD_M1007_g 0.0516583f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_18 VNB SCD 0.00798024f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_19 VNB N_A_423_315#_c_645_n 0.00300075f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_20 VNB N_A_423_315#_c_646_n 6.21324e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_21 VNB N_A_423_315#_c_647_n 0.00186605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_423_315#_c_648_n 0.0282104f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_23 VNB N_A_423_315#_c_649_n 0.00348698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_423_315#_c_650_n 0.00275863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_423_315#_c_651_n 0.0162167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_SCE_c_749_n 0.0172164f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_27 VNB N_SCE_c_750_n 0.0483627f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.59
cc_28 VNB N_SCE_c_751_n 0.0183888f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_29 VNB N_SCE_c_752_n 0.0274276f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_30 VNB N_SCE_c_753_n 0.00477854f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_31 VNB N_SCE_c_754_n 0.00357502f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_32 VNB SCE 0.00199642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB SCE 0.00480114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_SCE_c_757_n 0.0272237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_D_M1023_g 0.0472628f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_36 VNB N_A_193_47#_c_889_n 0.0133397f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_37 VNB N_A_193_47#_c_890_n 0.00420241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_193_47#_M1015_g 0.0199586f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_39 VNB N_A_193_47#_c_892_n 0.00878847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_193_47#_c_893_n 0.0180676f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_41 VNB N_A_193_47#_c_894_n 0.00302102f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_42 VNB N_A_193_47#_c_895_n 0.0312104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_193_47#_c_896_n 0.00454848f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_44 VNB N_A_193_47#_c_897_n 0.0292214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_193_47#_c_898_n 0.00651836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_193_47#_c_899_n 0.0012554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_193_47#_c_900_n 0.0218885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_193_47#_c_901_n 0.00235584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_193_47#_c_902_n 0.00200585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_193_47#_c_903_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_193_47#_c_904_n 0.0249277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_193_47#_c_905_n 0.00497848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_193_47#_c_906_n 0.0184534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1107_21#_M1038_g 0.0422736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_55 VNB N_A_1107_21#_c_1121_n 0.0192941f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_56 VNB N_A_1107_21#_c_1122_n 0.0018362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1107_21#_c_1123_n 0.00420076f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_58 VNB N_A_1107_21#_c_1124_n 0.0112435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1107_21#_c_1125_n 0.00590578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1107_21#_c_1126_n 0.0321305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_1266_n 0.0324101f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_62 VNB N_SET_B_M1011_g 0.00696184f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_63 VNB N_SET_B_M1044_g 0.0203534f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_64 VNB N_SET_B_M1004_g 0.02059f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_65 VNB N_SET_B_M1008_g 0.00796403f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_66 VNB SET_B 0.0076612f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.665
cc_67 VNB N_SET_B_c_1272_n 0.0154416f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_68 VNB N_SET_B_c_1273_n 0.00192349f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_69 VNB N_SET_B_c_1274_n 0.00323141f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_70 VNB N_SET_B_c_1275_n 0.00433788f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_71 VNB N_SET_B_c_1276_n 0.0319099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_931_47#_M1029_g 0.0258208f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_73 VNB N_A_931_47#_c_1396_n 0.00430594f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_74 VNB N_A_931_47#_c_1397_n 0.00789989f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_75 VNB N_A_931_47#_c_1398_n 0.00392752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_931_47#_c_1399_n 0.0143193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1400_21#_c_1500_n 0.0176574f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_78 VNB N_A_1400_21#_c_1501_n 0.034268f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_79 VNB N_A_1400_21#_M1031_g 0.0279648f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_80 VNB N_A_1400_21#_c_1503_n 0.011123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1400_21#_c_1504_n 0.00216927f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_82 VNB N_A_1400_21#_c_1505_n 0.00257402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1400_21#_c_1506_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1400_21#_c_1507_n 0.0195979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1400_21#_c_1508_n 0.00516344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1887_21#_M1005_g 0.0454209f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_87 VNB N_A_1887_21#_c_1659_n 0.0204896f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_88 VNB N_A_1887_21#_c_1660_n 0.0628379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1887_21#_c_1661_n 0.0171658f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_90 VNB N_A_1887_21#_c_1662_n 0.00811852f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_91 VNB N_A_1887_21#_c_1663_n 4.80417e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_92 VNB N_A_1887_21#_c_1664_n 0.0183894f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_93 VNB N_A_1887_21#_c_1665_n 0.0180366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_1887_21#_c_1666_n 0.00820903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_1887_21#_c_1667_n 0.0032181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_1887_21#_c_1668_n 0.00274082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_1714_47#_M1018_g 0.0219016f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_98 VNB N_A_1714_47#_c_1841_n 0.0117442f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_99 VNB N_A_1714_47#_c_1842_n 0.0114112f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_100 VNB N_A_1714_47#_c_1843_n 4.78869e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_1714_47#_c_1844_n 0.00186596f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_102 VNB N_A_1714_47#_c_1845_n 0.0176532f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_RESET_B_M1013_g 0.0349691f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.4
cc_104 VNB RESET_B 0.00386832f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_105 VNB N_RESET_B_c_1940_n 0.0287645f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.665
cc_106 VNB N_A_2596_47#_c_1974_n 0.0072656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_A_2596_47#_c_1975_n 0.00526785f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_108 VNB N_A_2596_47#_c_1976_n 0.0261462f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_109 VNB N_A_2596_47#_c_1977_n 2.8602e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_110 VNB N_A_2596_47#_c_1978_n 0.0201038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VPWR_c_2026_n 0.592346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_A_453_363#_c_2238_n 0.00615118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_A_453_363#_c_2239_n 0.00639648f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_114 VNB N_A_453_363#_c_2240_n 0.00623774f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_115 VNB N_A_453_363#_c_2241_n 0.00860491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_A_453_363#_c_2242_n 0.00211397f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_117 VNB N_A_453_363#_c_2243_n 0.00637751f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_453_363#_c_2244_n 0.00279367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_A_453_363#_c_2245_n 0.0142904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_Q_N_c_2371_n 0.00376073f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_121 VNB Q_N 0.00140118f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_122 VNB N_Q_N_c_2373_n 0.00366681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_Q_c_2402_n 0.00494099f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_124 VNB N_Q_c_2403_n 0.0229347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB Q 0.0170421f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_126 VNB N_VGND_c_2418_n 4.12476e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_127 VNB N_VGND_c_2419_n 0.00892979f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_128 VNB N_VGND_c_2420_n 0.00280508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2421_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2422_n 0.00556104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2423_n 0.00245603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2424_n 0.00557257f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2425_n 0.00259569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2426_n 0.0568827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2427_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2428_n 0.0383919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2429_n 0.00513816f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2430_n 0.0404697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2431_n 0.0037591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2432_n 0.0153564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2433_n 0.0165418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2434_n 0.0446468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2435_n 0.0540331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2436_n 0.0289512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2437_n 0.0150576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2438_n 0.66078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2439_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2440_n 0.00478425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2441_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2442_n 0.00510472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2443_n 0.00430718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VPB N_CLK_c_305_n 0.0118979f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_153 VPB N_CLK_c_306_n 0.0184083f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_154 VPB N_CLK_c_307_n 0.0238007f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_155 VPB CLK 0.0178201f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_156 VPB N_CLK_c_303_n 0.0100928f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_157 VPB N_A_27_47#_M1000_g 0.0379063f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_158 VPB N_A_27_47#_M1010_g 0.0215869f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_159 VPB N_A_27_47#_M1033_g 0.020906f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_160 VPB N_A_27_47#_c_346_n 0.017753f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_161 VPB N_A_27_47#_c_347_n 0.00403587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_27_47#_c_360_n 0.00103857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_27_47#_c_351_n 0.00335104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_27_47#_c_352_n 0.00245106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_27_47#_c_363_n 0.00362242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_27_47#_c_364_n 0.0330865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_27_47#_c_365_n 0.00181346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_27_47#_c_366_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_27_47#_c_367_n 0.00165292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_27_47#_c_368_n 0.00361706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_27_47#_c_354_n 0.0119282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_27_47#_c_370_n 0.0269269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_27_47#_c_371_n 0.00575159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_27_47#_c_372_n 0.0282388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_27_47#_c_373_n 0.00514398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_27_47#_c_374_n 0.0125285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_SCD_M1007_g 0.00110945f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_178 VPB N_SCD_M1034_g 0.0216594f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_179 VPB SCD 0.0054215f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_180 VPB N_SCD_c_613_n 0.04309f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_181 VPB N_A_423_315#_c_652_n 0.0180058f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_182 VPB N_A_423_315#_c_653_n 0.0628939f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_183 VPB N_A_423_315#_c_654_n 0.00770302f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_184 VPB N_A_423_315#_c_655_n 0.00300738f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_185 VPB N_A_423_315#_c_656_n 0.00841999f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_186 VPB N_A_423_315#_c_649_n 0.00556026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_423_315#_c_658_n 0.00654809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_SCE_c_752_n 0.0321372f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_189 VPB N_SCE_c_759_n 0.0173506f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_190 VPB N_SCE_c_760_n 0.0252061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_SCE_c_761_n 0.0144423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_SCE_c_762_n 0.00545787f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_193 VPB SCE 0.0076776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_D_M1023_g 0.00324838f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_195 VPB N_D_M1014_g 0.036057f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_196 VPB D 0.0116166f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_197 VPB N_D_c_851_n 0.0385655f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_198 VPB N_A_193_47#_M1041_g 0.0466077f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_199 VPB N_A_193_47#_c_889_n 0.0183248f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_200 VPB N_A_193_47#_c_890_n 0.00338145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_193_47#_M1017_g 0.0221986f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_202 VPB N_A_193_47#_c_911_n 0.0038403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_193_47#_c_912_n 0.0288235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_193_47#_c_903_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_193_47#_c_906_n 0.0187495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1107_21#_M1038_g 0.0150734f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_207 VPB N_A_1107_21#_M1036_g 0.0210587f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_208 VPB N_A_1107_21#_M1047_g 0.0317411f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_209 VPB N_A_1107_21#_c_1130_n 0.0055347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_A_1107_21#_c_1123_n 0.00619371f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_211 VPB N_A_1107_21#_c_1132_n 0.00575673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1107_21#_c_1133_n 0.0308181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1107_21#_c_1126_n 0.00659461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_SET_B_M1011_g 0.0508831f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_215 VPB N_SET_B_M1008_g 0.0496972f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_216 VPB N_A_931_47#_M1037_g 0.0203673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_217 VPB N_A_931_47#_c_1401_n 0.0121994f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_218 VPB N_A_931_47#_c_1397_n 0.00789134f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_219 VPB N_A_931_47#_c_1398_n 0.00271559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_931_47#_c_1399_n 0.0166794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1400_21#_c_1501_n 0.0218089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_222 VPB N_A_1400_21#_M1032_g 0.0205161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1400_21#_M1030_g 0.0210669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1400_21#_c_1512_n 0.0018943f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_225 VPB N_A_1400_21#_c_1513_n 0.0051975f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_226 VPB N_A_1400_21#_c_1506_n 0.00162652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1400_21#_c_1515_n 0.0327539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1400_21#_c_1516_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_1400_21#_c_1517_n 0.00737873f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_A_1400_21#_c_1518_n 0.00331979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1400_21#_c_1507_n 0.025869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_1400_21#_c_1508_n 0.00361429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_1887_21#_M1005_g 0.0159956f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_234 VPB N_A_1887_21#_M1042_g 0.021027f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_235 VPB N_A_1887_21#_M1039_g 0.0245592f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_236 VPB N_A_1887_21#_c_1661_n 0.00533941f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_237 VPB N_A_1887_21#_c_1663_n 0.0131679f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_238 VPB N_A_1887_21#_c_1674_n 0.0188715f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_239 VPB N_A_1887_21#_c_1675_n 0.0180753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_1887_21#_c_1676_n 0.00423323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_1887_21#_c_1677_n 0.0329665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_A_1887_21#_c_1678_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_A_1887_21#_c_1667_n 0.00331106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_A_1887_21#_c_1680_n 0.0072909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_A_1887_21#_c_1681_n 0.0016887f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_A_1887_21#_c_1668_n 2.41561e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_A_1714_47#_M1024_g 0.021833f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_248 VPB N_A_1714_47#_c_1847_n 0.0117899f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_249 VPB N_A_1714_47#_c_1842_n 0.00583428f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_250 VPB N_A_1714_47#_c_1843_n 7.45241e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_A_1714_47#_c_1844_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_252 VPB N_A_1714_47#_c_1845_n 0.00898586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_RESET_B_M1006_g 0.0248581f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_254 VPB RESET_B 9.55576e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_255 VPB N_RESET_B_c_1940_n 0.00925958f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_256 VPB N_A_2596_47#_M1002_g 0.0242997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_A_2596_47#_c_1980_n 0.013369f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_258 VPB N_A_2596_47#_c_1975_n 0.00520524f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_259 VPB N_A_2596_47#_c_1976_n 0.00598454f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_260 VPB N_VPWR_c_2027_n 0.00106376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_2028_n 0.00822796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_2029_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_2030_n 0.00313724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_2031_n 0.00562862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_2032_n 0.00358969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_2033_n 0.0292737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_2034_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_2035_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_2036_n 0.022998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_2037_n 0.0154511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_2038_n 0.0164006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_2039_n 0.0423496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_2040_n 0.0534515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_2041_n 0.0591311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_2042_n 0.0306954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_2043_n 0.0291788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_2044_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_2026_n 0.0758686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_2046_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_2047_n 0.00531184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_2048_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_2049_n 0.00609488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_2050_n 0.00928062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_2051_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_2052_n 0.00440561f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_286 VPB N_A_453_363#_c_2246_n 0.00565224f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.445
cc_287 VPB N_A_453_363#_c_2247_n 0.00638424f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_A_453_363#_c_2240_n 0.00227448f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_289 VPB N_A_453_363#_c_2242_n 3.39779e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_290 VPB N_A_453_363#_c_2243_n 0.00336519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB N_A_453_363#_c_2244_n 8.04394e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_292 VPB N_A_453_363#_c_2245_n 0.0146808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_293 VPB N_Q_N_c_2374_n 0.00137514f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_294 VPB N_Q_N_c_2371_n 0.00384084f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_295 VPB Q_N 0.00760446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_296 VPB N_Q_c_2405_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_297 VPB N_Q_c_2403_n 0.0137089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_298 VPB Q 0.0280643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_299 N_CLK_c_300_n N_A_27_47#_M1027_g 0.0200643f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_300 CLK N_A_27_47#_M1027_g 3.07529e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_301 N_CLK_c_304_n N_A_27_47#_M1027_g 0.00498861f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_302 N_CLK_c_307_n N_A_27_47#_M1000_g 0.0280586f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_303 CLK N_A_27_47#_M1000_g 5.68848e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_304 N_CLK_c_303_n N_A_27_47#_M1000_g 0.00521293f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_305 N_CLK_c_300_n N_A_27_47#_c_349_n 0.00685438f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_306 N_CLK_c_301_n N_A_27_47#_c_349_n 0.00799602f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_307 CLK N_A_27_47#_c_349_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_308 N_CLK_c_301_n N_A_27_47#_c_350_n 0.00621081f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_309 CLK N_A_27_47#_c_350_n 0.0148236f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_310 N_CLK_c_303_n N_A_27_47#_c_350_n 3.2891e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_311 N_CLK_c_306_n N_A_27_47#_c_360_n 0.0129431f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_312 N_CLK_c_307_n N_A_27_47#_c_360_n 0.0013404f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_313 CLK N_A_27_47#_c_360_n 0.00690269f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_314 N_CLK_c_301_n N_A_27_47#_c_351_n 0.00191059f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_315 N_CLK_c_307_n N_A_27_47#_c_351_n 0.00441254f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_316 CLK N_A_27_47#_c_351_n 0.0517134f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_317 N_CLK_c_303_n N_A_27_47#_c_351_n 0.00100166f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_318 N_CLK_c_304_n N_A_27_47#_c_351_n 0.00247465f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_319 N_CLK_c_306_n N_A_27_47#_c_363_n 2.18052e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_320 N_CLK_c_307_n N_A_27_47#_c_363_n 0.00374438f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_321 CLK N_A_27_47#_c_363_n 0.0157801f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_322 N_CLK_c_303_n N_A_27_47#_c_363_n 2.59784e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_323 N_CLK_c_306_n N_A_27_47#_c_365_n 0.00106507f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_324 CLK N_A_27_47#_c_354_n 0.00162145f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_325 N_CLK_c_303_n N_A_27_47#_c_354_n 0.0169859f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_326 N_CLK_c_306_n N_VPWR_c_2027_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_327 N_CLK_c_306_n N_VPWR_c_2037_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_328 N_CLK_c_306_n N_VPWR_c_2026_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_329 N_CLK_c_300_n N_VGND_c_2418_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_330 N_CLK_c_300_n N_VGND_c_2432_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_331 N_CLK_c_301_n N_VGND_c_2432_n 4.87495e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_332 N_CLK_c_300_n N_VGND_c_2438_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_364_n N_SCD_M1034_g 0.00922354f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_364_n SCD 0.00832905f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_364_n N_SCD_c_613_n 8.81844e-19 $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_336 N_A_27_47#_c_354_n N_SCD_c_613_n 0.00498361f $X=0.89 $Y=1.235 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_364_n N_A_423_315#_c_652_n 0.00654011f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_364_n N_A_423_315#_c_653_n 0.0080054f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_364_n N_A_423_315#_c_655_n 0.00712494f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_364_n N_A_423_315#_c_656_n 0.0146914f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_c_364_n N_A_423_315#_c_658_n 0.0162289f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_c_364_n N_SCE_c_752_n 0.0020833f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_343 N_A_27_47#_c_364_n N_SCE_c_760_n 0.0106145f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_344 N_A_27_47#_c_364_n N_SCE_c_762_n 0.00392465f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_345 N_A_27_47#_c_364_n SCE 0.0117724f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_345_n N_D_M1023_g 0.0212393f $X=4.58 $Y=0.705 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_364_n N_D_M1014_g 0.00707191f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_348 N_A_27_47#_c_364_n D 0.0200936f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_364_n N_D_c_851_n 9.34945e-19 $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_350 N_A_27_47#_c_364_n N_A_193_47#_M1000_d 6.81311e-19 $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_M1010_g N_A_193_47#_M1041_g 0.0190155f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_352_n N_A_193_47#_M1041_g 0.00534395f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_353 N_A_27_47#_c_364_n N_A_193_47#_M1041_g 0.00696374f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_367_n N_A_193_47#_M1041_g 5.24592e-19 $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_370_n N_A_193_47#_M1041_g 0.0174486f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_371_n N_A_193_47#_M1041_g 0.00867228f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_352_n N_A_193_47#_c_889_n 0.010154f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_366_n N_A_193_47#_c_889_n 3.83457e-19 $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_c_370_n N_A_193_47#_c_889_n 0.0212221f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_371_n N_A_193_47#_c_889_n 0.00654686f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_352_n N_A_193_47#_c_890_n 0.00203307f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_353_n N_A_193_47#_c_890_n 0.0232669f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_345_n N_A_193_47#_M1015_g 0.0127842f $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_352_n N_A_193_47#_M1015_g 4.45841e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_353_n N_A_193_47#_M1015_g 0.0214266f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1025_g N_A_193_47#_c_893_n 0.0131194f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_368_n N_A_193_47#_M1017_g 0.00133927f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_372_n N_A_193_47#_M1017_g 0.0192968f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_373_n N_A_193_47#_M1017_g 6.52047e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_347_n N_A_193_47#_c_894_n 2.62384e-19 $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_M1025_g N_A_193_47#_c_894_n 0.00310082f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_347_n N_A_193_47#_c_895_n 0.0206253f $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_M1025_g N_A_193_47#_c_895_n 0.0213524f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_346_n N_A_193_47#_c_896_n 0.0110233f $X=8.96 $Y=1.32 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_347_n N_A_193_47#_c_896_n 0.00356667f $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_M1025_g N_A_193_47#_c_896_n 0.00638693f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_373_n N_A_193_47#_c_896_n 0.00682571f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_346_n N_A_193_47#_c_911_n 0.00852739f $X=8.96 $Y=1.32 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_368_n N_A_193_47#_c_911_n 0.00483121f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_372_n N_A_193_47#_c_911_n 5.88448e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_373_n N_A_193_47#_c_911_n 0.0168759f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_374_n N_A_193_47#_c_911_n 0.00347329f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_346_n N_A_193_47#_c_912_n 0.0213022f $X=8.96 $Y=1.32 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_368_n N_A_193_47#_c_912_n 0.00219663f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_372_n N_A_193_47#_c_912_n 0.0169266f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_373_n N_A_193_47#_c_912_n 0.00153059f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_352_n N_A_193_47#_c_897_n 0.0155618f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_353_n N_A_193_47#_c_897_n 0.00553622f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_M1027_g N_A_193_47#_c_898_n 0.00656242f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_349_n N_A_193_47#_c_898_n 0.00215974f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_351_n N_A_193_47#_c_898_n 0.00508333f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_352_n N_A_193_47#_c_899_n 0.00934078f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_372_n N_A_193_47#_c_900_n 2.37019e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_366_n N_A_193_47#_c_901_n 0.111295f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_352_n N_A_193_47#_c_902_n 4.74166e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_346_n N_A_193_47#_c_903_n 3.23054e-19 $X=8.96 $Y=1.32 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_347_n N_A_193_47#_c_903_n 9.01357e-19 $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_373_n N_A_193_47#_c_903_n 0.00149027f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_352_n N_A_193_47#_c_904_n 0.00674133f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_345_n N_A_193_47#_c_905_n 4.90539e-19 $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_352_n N_A_193_47#_c_905_n 0.0210004f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_353_n N_A_193_47#_c_905_n 0.00154674f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_403 N_A_27_47#_c_370_n N_A_193_47#_c_905_n 3.18577e-19 $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_404 N_A_27_47#_c_371_n N_A_193_47#_c_905_n 0.00339609f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_405 N_A_27_47#_M1027_g N_A_193_47#_c_906_n 0.0233345f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_349_n N_A_193_47#_c_906_n 0.0115937f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_407 N_A_27_47#_c_476_p N_A_193_47#_c_906_n 0.00802121f $X=0.72 $Y=1.795 $X2=0
+ $Y2=0
cc_408 N_A_27_47#_c_351_n N_A_193_47#_c_906_n 0.0685543f $X=0.75 $Y=1.235 $X2=0
+ $Y2=0
cc_409 N_A_27_47#_c_364_n N_A_193_47#_c_906_n 0.0268048f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_410 N_A_27_47#_c_365_n N_A_193_47#_c_906_n 0.00184875f $X=0.835 $Y=1.87 $X2=0
+ $Y2=0
cc_411 N_A_27_47#_c_352_n N_A_1107_21#_M1038_g 5.35023e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_412 N_A_27_47#_c_366_n N_A_1107_21#_M1036_g 0.00197541f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_M1033_g N_A_1107_21#_M1047_g 0.0164618f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_414 N_A_27_47#_c_347_n N_A_1107_21#_M1047_g 0.00557814f $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_c_366_n N_A_1107_21#_M1047_g 0.00750594f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_372_n N_A_1107_21#_M1047_g 0.00910409f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_373_n N_A_1107_21#_M1047_g 0.00264318f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_366_n N_A_1107_21#_c_1130_n 0.0240118f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_419 N_A_27_47#_c_366_n N_A_1107_21#_c_1143_n 0.0279846f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_c_366_n N_A_1107_21#_c_1132_n 0.0141612f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_421 N_A_27_47#_M1010_g N_A_1107_21#_c_1133_n 0.0161827f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_366_n N_A_1107_21#_c_1133_n 0.00193898f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_370_n N_A_1107_21#_c_1133_n 0.00927772f $X=5.04 $Y=1.74
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_366_n N_A_1107_21#_c_1148_n 0.00959465f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_425 N_A_27_47#_c_347_n N_A_1107_21#_c_1126_n 0.0027239f $X=8.58 $Y=1.32 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_M1025_g N_SET_B_c_1272_n 0.00574114f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_M1010_g N_A_931_47#_c_1405_n 0.0091014f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_364_n N_A_931_47#_c_1405_n 2.09728e-19 $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_366_n N_A_931_47#_c_1405_n 0.00506942f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_367_n N_A_931_47#_c_1405_n 0.00303545f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_370_n N_A_931_47#_c_1405_n 0.00186639f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_432 N_A_27_47#_c_371_n N_A_931_47#_c_1405_n 0.0152514f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_433 N_A_27_47#_c_352_n N_A_931_47#_c_1411_n 0.00676006f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_434 N_A_27_47#_c_353_n N_A_931_47#_c_1411_n 9.25786e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_435 N_A_27_47#_M1010_g N_A_931_47#_c_1401_n 0.00650943f $X=5.01 $Y=2.275
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_352_n N_A_931_47#_c_1401_n 0.00666284f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_366_n N_A_931_47#_c_1401_n 0.013911f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_438 N_A_27_47#_c_367_n N_A_931_47#_c_1401_n 0.00149623f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_370_n N_A_931_47#_c_1401_n 0.00203066f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_440 N_A_27_47#_c_371_n N_A_931_47#_c_1401_n 0.0282877f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_366_n N_A_931_47#_c_1397_n 0.00350894f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_352_n N_A_931_47#_c_1398_n 0.00728915f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_443 N_A_27_47#_c_366_n N_A_931_47#_c_1398_n 0.00456576f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_366_n N_A_1400_21#_M1032_g 0.00576309f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_366_n N_A_1400_21#_c_1506_n 0.00477237f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_346_n N_A_1400_21#_c_1515_n 0.00385681f $X=8.96 $Y=1.32
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_c_366_n N_A_1400_21#_c_1515_n 0.0139809f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_448 N_A_27_47#_c_368_n N_A_1400_21#_c_1515_n 0.0255925f $X=8.51 $Y=1.87 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_372_n N_A_1400_21#_c_1515_n 0.00176885f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_c_373_n N_A_1400_21#_c_1515_n 0.00661378f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_c_374_n N_A_1400_21#_c_1515_n 0.00371524f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_c_366_n N_A_1400_21#_c_1516_n 0.0264578f $X=8.365 $Y=1.87
+ $X2=0 $Y2=0
cc_453 N_A_27_47#_c_372_n N_A_1400_21#_c_1516_n 7.96394e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_454 N_A_27_47#_c_373_n N_A_1400_21#_c_1516_n 0.00130051f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_455 N_A_27_47#_c_374_n N_A_1400_21#_c_1516_n 7.27878e-19 $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_456 N_A_27_47#_c_366_n N_A_1400_21#_c_1517_n 0.020032f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_372_n N_A_1400_21#_c_1517_n 6.45403e-19 $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_458 N_A_27_47#_c_373_n N_A_1400_21#_c_1517_n 0.00461622f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_459 N_A_27_47#_c_374_n N_A_1400_21#_c_1517_n 0.00148716f $X=8.445 $Y=1.575
+ $X2=0 $Y2=0
cc_460 N_A_27_47#_M1025_g N_A_1887_21#_M1005_g 0.0428093f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_461 N_A_27_47#_M1033_g N_A_1714_47#_c_1852_n 0.00496872f $X=8.505 $Y=2.275
+ $X2=0 $Y2=0
cc_462 N_A_27_47#_c_368_n N_A_1714_47#_c_1852_n 0.00187313f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_463 N_A_27_47#_c_373_n N_A_1714_47#_c_1852_n 0.00141396f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_464 N_A_27_47#_M1025_g N_A_1714_47#_c_1855_n 0.00969843f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_465 N_A_27_47#_M1025_g N_A_1714_47#_c_1841_n 0.0106063f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_466 N_A_27_47#_c_368_n N_A_1714_47#_c_1847_n 0.00214622f $X=8.51 $Y=1.87
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_c_373_n N_A_1714_47#_c_1847_n 0.0013353f $X=8.445 $Y=1.74
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_M1025_g N_A_1714_47#_c_1843_n 0.00155103f $X=9.035 $Y=0.415
+ $X2=0 $Y2=0
cc_469 N_A_27_47#_c_476_p N_VPWR_M1026_d 7.14517e-19 $X=0.72 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_470 N_A_27_47#_c_365_n N_VPWR_M1026_d 0.00181761f $X=0.835 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_471 N_A_27_47#_c_366_n N_VPWR_M1032_d 0.00670518f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_M1000_g N_VPWR_c_2027_n 0.00837918f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_360_n N_VPWR_c_2027_n 0.00328949f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_476_p N_VPWR_c_2027_n 0.0133733f $X=0.72 $Y=1.795 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_363_n N_VPWR_c_2027_n 0.0127225f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_364_n N_VPWR_c_2027_n 2.78216e-19 $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_365_n N_VPWR_c_2027_n 0.00348405f $X=0.835 $Y=1.87 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_M1000_g N_VPWR_c_2028_n 0.00230379f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_364_n N_VPWR_c_2028_n 0.0156468f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_480 N_A_27_47#_c_364_n N_VPWR_c_2029_n 0.00411755f $X=4.685 $Y=1.87 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_366_n N_VPWR_c_2030_n 0.00160449f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_366_n N_VPWR_c_2031_n 0.0137399f $X=8.365 $Y=1.87 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_360_n N_VPWR_c_2037_n 0.0018545f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_363_n N_VPWR_c_2037_n 0.0123893f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_485 N_A_27_47#_M1000_g N_VPWR_c_2038_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_M1010_g N_VPWR_c_2040_n 0.00367119f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_487 N_A_27_47#_M1033_g N_VPWR_c_2041_n 0.00424681f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_373_n N_VPWR_c_2041_n 0.00254851f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_M1000_g N_VPWR_c_2026_n 0.00536257f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_M1010_g N_VPWR_c_2026_n 0.00562272f $X=5.01 $Y=2.275 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_M1033_g N_VPWR_c_2026_n 0.0061745f $X=8.505 $Y=2.275 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_360_n N_VPWR_c_2026_n 0.00394611f $X=0.605 $Y=1.88 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_363_n N_VPWR_c_2026_n 0.00665993f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_364_n N_VPWR_c_2026_n 0.18557f $X=4.685 $Y=1.87 $X2=0 $Y2=0
cc_495 N_A_27_47#_c_365_n N_VPWR_c_2026_n 0.01448f $X=0.835 $Y=1.87 $X2=0 $Y2=0
cc_496 N_A_27_47#_c_366_n N_VPWR_c_2026_n 0.159156f $X=8.365 $Y=1.87 $X2=0 $Y2=0
cc_497 N_A_27_47#_c_367_n N_VPWR_c_2026_n 0.0160117f $X=4.975 $Y=1.87 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_c_368_n N_VPWR_c_2026_n 0.0148451f $X=8.51 $Y=1.87 $X2=0 $Y2=0
cc_499 N_A_27_47#_c_371_n N_VPWR_c_2026_n 3.19863e-19 $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_372_n N_VPWR_c_2026_n 3.05853e-19 $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_373_n N_VPWR_c_2026_n 0.00131252f $X=8.445 $Y=1.74 $X2=0
+ $Y2=0
cc_502 N_A_27_47#_c_364_n A_381_363# 0.00298073f $X=4.685 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_503 N_A_27_47#_c_364_n N_A_453_363#_c_2246_n 0.0156835f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_504 N_A_27_47#_c_364_n N_A_453_363#_c_2247_n 0.0104101f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_505 N_A_27_47#_c_364_n N_A_453_363#_c_2240_n 0.00714524f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_506 N_A_27_47#_c_364_n N_A_453_363#_c_2241_n 0.0497172f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_507 N_A_27_47#_c_364_n N_A_453_363#_c_2242_n 0.0128797f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_508 N_A_27_47#_c_364_n N_A_453_363#_c_2243_n 0.00118055f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_509 N_A_27_47#_c_352_n N_A_453_363#_c_2244_n 0.00749938f $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_510 N_A_27_47#_c_353_n N_A_453_363#_c_2244_n 2.04896e-19 $X=4.71 $Y=0.87
+ $X2=0 $Y2=0
cc_511 N_A_27_47#_c_364_n N_A_453_363#_c_2244_n 0.0130335f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_512 N_A_27_47#_c_345_n N_A_453_363#_c_2245_n 0.00475032f $X=4.58 $Y=0.705
+ $X2=0 $Y2=0
cc_513 N_A_27_47#_c_352_n N_A_453_363#_c_2245_n 0.0620374f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_364_n N_A_453_363#_c_2245_n 0.0188924f $X=4.685 $Y=1.87
+ $X2=0 $Y2=0
cc_515 N_A_27_47#_c_367_n N_A_453_363#_c_2245_n 0.00185048f $X=4.975 $Y=1.87
+ $X2=0 $Y2=0
cc_516 N_A_27_47#_c_371_n N_A_453_363#_c_2245_n 0.0281945f $X=5.04 $Y=1.74 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_366_n A_1351_329# 0.00110713f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_518 N_A_27_47#_c_366_n A_1572_329# 0.00532504f $X=8.365 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_519 N_A_27_47#_c_349_n N_VGND_M1045_d 0.00162876f $X=0.605 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_520 N_A_27_47#_M1027_g N_VGND_c_2418_n 0.00826882f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_349_n N_VGND_c_2418_n 0.0165953f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_354_n N_VGND_c_2418_n 5.88506e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_M1027_g N_VGND_c_2419_n 0.00319233f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_524 N_A_27_47#_M1025_g N_VGND_c_2423_n 0.00124887f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_525 N_A_27_47#_c_345_n N_VGND_c_2426_n 0.00556304f $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_526 N_A_27_47#_c_352_n N_VGND_c_2426_n 0.00113905f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_527 N_A_27_47#_c_353_n N_VGND_c_2426_n 2.48118e-19 $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_528 N_A_27_47#_M1025_g N_VGND_c_2430_n 0.00359964f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_529 N_A_27_47#_c_598_p N_VGND_c_2432_n 0.00735289f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_530 N_A_27_47#_c_349_n N_VGND_c_2432_n 0.00243651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_531 N_A_27_47#_M1027_g N_VGND_c_2433_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_532 N_A_27_47#_M1045_s N_VGND_c_2438_n 0.00358206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_A_27_47#_M1027_g N_VGND_c_2438_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_534 N_A_27_47#_c_345_n N_VGND_c_2438_n 0.00678262f $X=4.58 $Y=0.705 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_M1025_g N_VGND_c_2438_n 0.00563077f $X=9.035 $Y=0.415 $X2=0
+ $Y2=0
cc_536 N_A_27_47#_c_598_p N_VGND_c_2438_n 0.00626856f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_537 N_A_27_47#_c_349_n N_VGND_c_2438_n 0.0057651f $X=0.605 $Y=0.72 $X2=0
+ $Y2=0
cc_538 N_A_27_47#_c_352_n N_VGND_c_2438_n 0.00122477f $X=4.71 $Y=0.87 $X2=0
+ $Y2=0
cc_539 N_SCD_M1034_g N_A_423_315#_c_652_n 0.0310295f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_540 N_SCD_c_613_n N_A_423_315#_c_654_n 0.0310295f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_541 N_SCD_M1007_g N_SCE_c_749_n 0.033964f $X=1.83 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_542 N_SCD_M1007_g N_SCE_c_754_n 0.00423581f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_543 N_SCD_M1007_g SCE 0.00547993f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_544 N_SCD_M1007_g SCE 0.0141807f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_545 SCD SCE 0.0399718f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_546 N_SCD_M1007_g N_SCE_c_757_n 0.0205263f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_547 N_SCD_M1007_g N_A_193_47#_c_897_n 0.0122391f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_548 SCD N_A_193_47#_c_897_n 0.00983418f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_549 N_SCD_c_613_n N_A_193_47#_c_897_n 7.56832e-19 $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_550 N_SCD_M1007_g N_A_193_47#_c_898_n 0.00180888f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_551 N_SCD_M1007_g N_A_193_47#_c_906_n 0.00844652f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_552 N_SCD_M1034_g N_A_193_47#_c_906_n 0.00452759f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_553 SCD N_A_193_47#_c_906_n 0.0470439f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_554 N_SCD_c_613_n N_A_193_47#_c_906_n 0.00114684f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_555 N_SCD_M1034_g N_VPWR_c_2028_n 0.0156084f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_556 SCD N_VPWR_c_2028_n 0.0157864f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_557 N_SCD_c_613_n N_VPWR_c_2028_n 0.00226856f $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_558 N_SCD_M1034_g N_VPWR_c_2039_n 0.00442511f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_559 N_SCD_M1034_g N_VPWR_c_2026_n 0.00418686f $X=1.83 $Y=2.135 $X2=0 $Y2=0
cc_560 N_SCD_M1034_g N_A_453_363#_c_2246_n 0.00148049f $X=1.83 $Y=2.135 $X2=0
+ $Y2=0
cc_561 N_SCD_M1007_g N_VGND_c_2419_n 0.00525265f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_562 SCD N_VGND_c_2419_n 0.00628942f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_563 N_SCD_c_613_n N_VGND_c_2419_n 8.59131e-19 $X=1.83 $Y=1.49 $X2=0 $Y2=0
cc_564 N_SCD_M1007_g N_VGND_c_2434_n 0.00585385f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_565 N_SCD_M1007_g N_VGND_c_2438_n 0.00764087f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_566 N_A_423_315#_c_653_n N_SCE_c_750_n 0.00587794f $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_567 N_A_423_315#_c_656_n N_SCE_c_750_n 4.1633e-19 $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_568 N_A_423_315#_c_645_n N_SCE_c_750_n 0.00142101f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_569 N_A_423_315#_c_646_n N_SCE_c_750_n 0.00721303f $X=3.125 $Y=0.71 $X2=0
+ $Y2=0
cc_570 N_A_423_315#_c_645_n N_SCE_c_751_n 0.007706f $X=3.475 $Y=0.71 $X2=0 $Y2=0
cc_571 N_A_423_315#_c_651_n N_SCE_c_751_n 0.0157579f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_572 N_A_423_315#_c_653_n N_SCE_c_752_n 0.0213525f $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_573 N_A_423_315#_c_656_n N_SCE_c_752_n 0.0109878f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_574 N_A_423_315#_c_658_n N_SCE_c_752_n 0.010066f $X=2.905 $Y=1.66 $X2=0 $Y2=0
cc_575 N_A_423_315#_c_650_n N_SCE_c_752_n 0.00695886f $X=3.622 $Y=1.095 $X2=0
+ $Y2=0
cc_576 N_A_423_315#_c_656_n N_SCE_c_760_n 0.00779447f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_577 N_A_423_315#_c_645_n N_SCE_c_753_n 0.00574578f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_578 N_A_423_315#_c_647_n N_SCE_c_753_n 0.00695886f $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_579 N_A_423_315#_c_648_n N_SCE_c_753_n 0.0207451f $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_580 N_A_423_315#_c_651_n N_SCE_c_753_n 9.51141e-19 $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_581 N_A_423_315#_c_655_n N_SCE_c_762_n 0.00990576f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_582 N_A_423_315#_c_654_n N_SCE_c_754_n 9.48832e-19 $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_583 N_A_423_315#_c_654_n SCE 0.00531279f $X=2.265 $Y=1.65 $X2=0 $Y2=0
cc_584 N_A_423_315#_c_654_n N_SCE_c_757_n 0.00742685f $X=2.265 $Y=1.65 $X2=0
+ $Y2=0
cc_585 N_A_423_315#_c_647_n N_D_M1023_g 0.00105116f $X=3.685 $Y=0.93 $X2=0 $Y2=0
cc_586 N_A_423_315#_c_649_n N_D_M1023_g 0.00175438f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_587 N_A_423_315#_c_651_n N_D_M1023_g 0.0616329f $X=3.685 $Y=0.765 $X2=0 $Y2=0
cc_588 N_A_423_315#_c_656_n D 0.0135689f $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_589 N_A_423_315#_c_649_n D 0.017414f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_590 N_A_423_315#_c_656_n N_D_c_851_n 4.98039e-19 $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_591 N_A_423_315#_c_648_n N_D_c_851_n 0.00265425f $X=3.685 $Y=0.93 $X2=0 $Y2=0
cc_592 N_A_423_315#_c_649_n N_D_c_851_n 0.00200746f $X=3.56 $Y=1.575 $X2=0 $Y2=0
cc_593 N_A_423_315#_c_645_n N_A_193_47#_c_897_n 0.0197158f $X=3.475 $Y=0.71
+ $X2=0 $Y2=0
cc_594 N_A_423_315#_c_646_n N_A_193_47#_c_897_n 0.00794081f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_595 N_A_423_315#_c_647_n N_A_193_47#_c_897_n 0.014943f $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_596 N_A_423_315#_c_648_n N_A_193_47#_c_897_n 0.00180177f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_597 N_A_423_315#_c_652_n N_VPWR_c_2028_n 0.0027725f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_598 N_A_423_315#_c_655_n N_VPWR_c_2029_n 0.0139381f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_599 N_A_423_315#_c_656_n N_VPWR_c_2029_n 0.00494232f $X=3.475 $Y=1.66 $X2=0
+ $Y2=0
cc_600 N_A_423_315#_c_652_n N_VPWR_c_2039_n 0.00516156f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_601 N_A_423_315#_c_655_n N_VPWR_c_2039_n 0.0118139f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_602 N_A_423_315#_M1035_s N_VPWR_c_2026_n 0.00335142f $X=2.855 $Y=2.065 $X2=0
+ $Y2=0
cc_603 N_A_423_315#_c_652_n N_VPWR_c_2026_n 0.00685533f $X=2.19 $Y=1.725 $X2=0
+ $Y2=0
cc_604 N_A_423_315#_c_653_n N_VPWR_c_2026_n 2.96327e-19 $X=2.695 $Y=1.65 $X2=0
+ $Y2=0
cc_605 N_A_423_315#_c_655_n N_VPWR_c_2026_n 0.00308197f $X=2.98 $Y=2.3 $X2=0
+ $Y2=0
cc_606 N_A_423_315#_c_658_n N_VPWR_c_2026_n 0.00196684f $X=2.905 $Y=1.66 $X2=0
+ $Y2=0
cc_607 N_A_423_315#_c_707_p N_A_453_363#_c_2238_n 0.00220863f $X=3.04 $Y=0.47
+ $X2=0 $Y2=0
cc_608 N_A_423_315#_c_646_n N_A_453_363#_c_2238_n 0.0137055f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_609 N_A_423_315#_c_652_n N_A_453_363#_c_2246_n 0.00894778f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_610 N_A_423_315#_c_653_n N_A_453_363#_c_2246_n 0.00237707f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_611 N_A_423_315#_c_655_n N_A_453_363#_c_2246_n 0.0230656f $X=2.98 $Y=2.3
+ $X2=0 $Y2=0
cc_612 N_A_423_315#_c_652_n N_A_453_363#_c_2247_n 0.00320876f $X=2.19 $Y=1.725
+ $X2=0 $Y2=0
cc_613 N_A_423_315#_c_653_n N_A_453_363#_c_2247_n 0.0175674f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_614 N_A_423_315#_c_658_n N_A_453_363#_c_2247_n 0.0225881f $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_615 N_A_423_315#_c_707_p N_A_453_363#_c_2239_n 0.0232733f $X=3.04 $Y=0.47
+ $X2=0 $Y2=0
cc_616 N_A_423_315#_c_653_n N_A_453_363#_c_2240_n 0.00532216f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_617 N_A_423_315#_c_658_n N_A_453_363#_c_2240_n 6.00227e-19 $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_618 N_A_423_315#_c_656_n N_A_453_363#_c_2241_n 0.00811555f $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_619 N_A_423_315#_c_645_n N_A_453_363#_c_2241_n 0.00315275f $X=3.475 $Y=0.71
+ $X2=0 $Y2=0
cc_620 N_A_423_315#_c_648_n N_A_453_363#_c_2241_n 3.93982e-19 $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_621 N_A_423_315#_c_649_n N_A_453_363#_c_2241_n 0.0158823f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_622 N_A_423_315#_c_650_n N_A_453_363#_c_2241_n 0.00384754f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_623 N_A_423_315#_c_656_n N_A_453_363#_c_2242_n 0.00169392f $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_624 N_A_423_315#_c_646_n N_A_453_363#_c_2242_n 0.00141688f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_625 N_A_423_315#_c_649_n N_A_453_363#_c_2242_n 0.0011872f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_626 N_A_423_315#_c_658_n N_A_453_363#_c_2242_n 9.72289e-19 $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_627 N_A_423_315#_c_650_n N_A_453_363#_c_2242_n 0.00120978f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_628 N_A_423_315#_c_653_n N_A_453_363#_c_2243_n 0.00101345f $X=2.695 $Y=1.65
+ $X2=0 $Y2=0
cc_629 N_A_423_315#_c_656_n N_A_453_363#_c_2243_n 5.57877e-19 $X=3.475 $Y=1.66
+ $X2=0 $Y2=0
cc_630 N_A_423_315#_c_646_n N_A_453_363#_c_2243_n 0.00610396f $X=3.125 $Y=0.71
+ $X2=0 $Y2=0
cc_631 N_A_423_315#_c_658_n N_A_453_363#_c_2243_n 0.0185169f $X=2.905 $Y=1.66
+ $X2=0 $Y2=0
cc_632 N_A_423_315#_c_650_n N_A_453_363#_c_2243_n 0.00944685f $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_633 N_A_423_315#_c_649_n N_A_453_363#_c_2244_n 0.00152543f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_634 N_A_423_315#_c_650_n N_A_453_363#_c_2244_n 4.68942e-19 $X=3.622 $Y=1.095
+ $X2=0 $Y2=0
cc_635 N_A_423_315#_c_645_n N_A_453_363#_c_2245_n 0.00482345f $X=3.475 $Y=0.71
+ $X2=0 $Y2=0
cc_636 N_A_423_315#_c_647_n N_A_453_363#_c_2245_n 0.00870657f $X=3.685 $Y=0.93
+ $X2=0 $Y2=0
cc_637 N_A_423_315#_c_649_n N_A_453_363#_c_2245_n 0.00442233f $X=3.56 $Y=1.575
+ $X2=0 $Y2=0
cc_638 N_A_423_315#_c_645_n N_VGND_M1012_d 0.00246138f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_639 N_A_423_315#_c_645_n N_VGND_c_2420_n 0.0177928f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_640 N_A_423_315#_c_648_n N_VGND_c_2420_n 4.49423e-19 $X=3.685 $Y=0.93 $X2=0
+ $Y2=0
cc_641 N_A_423_315#_c_651_n N_VGND_c_2420_n 0.00914963f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_642 N_A_423_315#_c_651_n N_VGND_c_2426_n 0.0046653f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_643 N_A_423_315#_c_707_p N_VGND_c_2434_n 0.0101366f $X=3.04 $Y=0.47 $X2=0
+ $Y2=0
cc_644 N_A_423_315#_c_645_n N_VGND_c_2434_n 0.00345019f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_645 N_A_423_315#_M1012_s N_VGND_c_2438_n 0.00190491f $X=2.915 $Y=0.235 $X2=0
+ $Y2=0
cc_646 N_A_423_315#_c_707_p N_VGND_c_2438_n 0.00346716f $X=3.04 $Y=0.47 $X2=0
+ $Y2=0
cc_647 N_A_423_315#_c_645_n N_VGND_c_2438_n 0.00513527f $X=3.475 $Y=0.71 $X2=0
+ $Y2=0
cc_648 N_A_423_315#_c_651_n N_VGND_c_2438_n 0.00398879f $X=3.685 $Y=0.765 $X2=0
+ $Y2=0
cc_649 N_SCE_c_752_n N_D_M1023_g 0.00323589f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_650 N_SCE_c_752_n N_D_M1014_g 0.00214944f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_651 N_SCE_c_760_n N_D_M1014_g 0.0334116f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_652 N_SCE_c_752_n D 0.00166353f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_653 N_SCE_c_760_n D 0.0100165f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_654 N_SCE_c_752_n N_D_c_851_n 0.00552281f $X=3.265 $Y=1.835 $X2=0 $Y2=0
cc_655 N_SCE_c_750_n N_A_193_47#_c_897_n 0.0053068f $X=3.175 $Y=0.81 $X2=0 $Y2=0
cc_656 N_SCE_c_752_n N_A_193_47#_c_897_n 0.00239268f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_657 N_SCE_c_753_n N_A_193_47#_c_897_n 4.50186e-19 $X=3.257 $Y=0.81 $X2=0
+ $Y2=0
cc_658 N_SCE_c_754_n N_A_193_47#_c_897_n 0.0203775f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_659 SCE N_A_193_47#_c_897_n 0.0107956f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_660 SCE N_A_193_47#_c_897_n 0.00156771f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_661 N_SCE_c_757_n N_A_193_47#_c_897_n 0.00314883f $X=2.25 $Y=0.81 $X2=0 $Y2=0
cc_662 N_SCE_c_759_n N_VPWR_c_2029_n 0.00953982f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_663 N_SCE_c_760_n N_VPWR_c_2029_n 0.00200314f $X=3.61 $Y=1.91 $X2=0 $Y2=0
cc_664 N_SCE_c_761_n N_VPWR_c_2029_n 0.00920451f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_665 N_SCE_c_759_n N_VPWR_c_2039_n 0.0046653f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_666 N_SCE_c_761_n N_VPWR_c_2040_n 0.0046653f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_667 N_SCE_c_759_n N_VPWR_c_2026_n 0.00581646f $X=3.265 $Y=1.985 $X2=0 $Y2=0
cc_668 N_SCE_c_761_n N_VPWR_c_2026_n 0.00446764f $X=3.685 $Y=1.985 $X2=0 $Y2=0
cc_669 N_SCE_c_749_n N_A_453_363#_c_2238_n 0.00215187f $X=2.22 $Y=0.735 $X2=0
+ $Y2=0
cc_670 N_SCE_c_750_n N_A_453_363#_c_2238_n 0.0135177f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_671 N_SCE_c_751_n N_A_453_363#_c_2238_n 3.61202e-19 $X=3.25 $Y=0.735 $X2=0
+ $Y2=0
cc_672 N_SCE_c_752_n N_A_453_363#_c_2238_n 0.00458533f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_673 N_SCE_c_754_n N_A_453_363#_c_2238_n 0.0127619f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_674 SCE N_A_453_363#_c_2238_n 0.00830792f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_675 SCE N_A_453_363#_c_2238_n 0.00226589f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_676 N_SCE_c_757_n N_A_453_363#_c_2238_n 0.00224421f $X=2.25 $Y=0.81 $X2=0
+ $Y2=0
cc_677 N_SCE_c_752_n N_A_453_363#_c_2247_n 0.00460376f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_678 SCE N_A_453_363#_c_2247_n 0.0248247f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_679 N_SCE_c_750_n N_A_453_363#_c_2239_n 0.00657992f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_680 N_SCE_c_751_n N_A_453_363#_c_2239_n 8.04587e-19 $X=3.25 $Y=0.735 $X2=0
+ $Y2=0
cc_681 N_SCE_c_754_n N_A_453_363#_c_2239_n 0.00267477f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_682 N_SCE_c_750_n N_A_453_363#_c_2240_n 0.00119558f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_683 N_SCE_c_754_n N_A_453_363#_c_2240_n 0.00490238f $X=2.25 $Y=0.93 $X2=0
+ $Y2=0
cc_684 SCE N_A_453_363#_c_2240_n 0.0204381f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_685 N_SCE_c_757_n N_A_453_363#_c_2240_n 9.25794e-19 $X=2.25 $Y=0.81 $X2=0
+ $Y2=0
cc_686 N_SCE_c_752_n N_A_453_363#_c_2241_n 0.00696234f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_687 N_SCE_c_760_n N_A_453_363#_c_2241_n 5.63442e-19 $X=3.61 $Y=1.91 $X2=0
+ $Y2=0
cc_688 N_SCE_c_750_n N_A_453_363#_c_2242_n 0.00100011f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_689 N_SCE_c_752_n N_A_453_363#_c_2242_n 0.00229563f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_690 N_SCE_c_750_n N_A_453_363#_c_2243_n 0.0056856f $X=3.175 $Y=0.81 $X2=0
+ $Y2=0
cc_691 N_SCE_c_752_n N_A_453_363#_c_2243_n 0.00631075f $X=3.265 $Y=1.835 $X2=0
+ $Y2=0
cc_692 N_SCE_c_751_n N_VGND_c_2420_n 0.00409489f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_693 N_SCE_c_749_n N_VGND_c_2434_n 0.00537877f $X=2.22 $Y=0.735 $X2=0 $Y2=0
cc_694 N_SCE_c_750_n N_VGND_c_2434_n 0.00315686f $X=3.175 $Y=0.81 $X2=0 $Y2=0
cc_695 N_SCE_c_751_n N_VGND_c_2434_n 0.0042361f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_696 SCE N_VGND_c_2434_n 0.00824495f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_697 N_SCE_c_749_n N_VGND_c_2438_n 0.00695567f $X=2.22 $Y=0.735 $X2=0 $Y2=0
cc_698 N_SCE_c_750_n N_VGND_c_2438_n 0.00211039f $X=3.175 $Y=0.81 $X2=0 $Y2=0
cc_699 N_SCE_c_751_n N_VGND_c_2438_n 0.00704136f $X=3.25 $Y=0.735 $X2=0 $Y2=0
cc_700 N_SCE_c_754_n N_VGND_c_2438_n 0.00197531f $X=2.25 $Y=0.93 $X2=0 $Y2=0
cc_701 SCE N_VGND_c_2438_n 0.00364093f $X=2.01 $Y=0.425 $X2=0 $Y2=0
cc_702 SCE A_381_47# 0.00150833f $X=2.01 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_703 N_D_c_851_n N_A_193_47#_M1041_g 0.0186046f $X=4.105 $Y=1.49 $X2=0 $Y2=0
cc_704 N_D_M1023_g N_A_193_47#_c_890_n 0.0186046f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_705 N_D_M1023_g N_A_193_47#_c_897_n 0.00630058f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_706 N_D_M1014_g N_VPWR_c_2029_n 0.0014636f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_707 D N_VPWR_c_2029_n 0.0112011f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_708 N_D_M1014_g N_VPWR_c_2040_n 0.00585385f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_709 D N_VPWR_c_2040_n 0.00771405f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_710 N_D_M1014_g N_VPWR_c_2026_n 0.00659811f $X=4.105 $Y=2.275 $X2=0 $Y2=0
cc_711 D N_VPWR_c_2026_n 0.00345538f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_712 N_D_M1023_g N_A_453_363#_c_2241_n 0.00796014f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_713 D N_A_453_363#_c_2241_n 0.00855055f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_714 N_D_c_851_n N_A_453_363#_c_2241_n 5.10457e-19 $X=4.105 $Y=1.49 $X2=0
+ $Y2=0
cc_715 N_D_M1023_g N_A_453_363#_c_2244_n 0.00192517f $X=4.105 $Y=0.445 $X2=0
+ $Y2=0
cc_716 N_D_M1023_g N_A_453_363#_c_2245_n 0.017252f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_717 D N_A_453_363#_c_2245_n 0.0480833f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_718 D A_752_413# 0.00729005f $X=3.825 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_719 N_D_M1023_g N_VGND_c_2420_n 0.00188039f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_720 N_D_M1023_g N_VGND_c_2426_n 0.00585385f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_721 N_D_M1023_g N_VGND_c_2438_n 0.00646586f $X=4.105 $Y=0.445 $X2=0 $Y2=0
cc_722 N_A_193_47#_M1015_g N_A_1107_21#_M1038_g 0.0245694f $X=5.13 $Y=0.415
+ $X2=0 $Y2=0
cc_723 N_A_193_47#_c_892_n N_A_1107_21#_M1038_g 0.0105189f $X=5.13 $Y=1.245
+ $X2=0 $Y2=0
cc_724 N_A_193_47#_c_900_n N_A_1107_21#_M1038_g 7.74803e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_725 N_A_193_47#_c_902_n N_A_1107_21#_M1038_g 0.00642269f $X=5.29 $Y=0.85
+ $X2=0 $Y2=0
cc_726 N_A_193_47#_c_904_n N_A_1107_21#_M1038_g 0.0200662f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_727 N_A_193_47#_c_905_n N_A_1107_21#_M1038_g 0.00189958f $X=5.19 $Y=0.93
+ $X2=0 $Y2=0
cc_728 N_A_193_47#_c_893_n N_A_1107_21#_c_1121_n 0.0350413f $X=8.495 $Y=0.705
+ $X2=0 $Y2=0
cc_729 N_A_193_47#_c_894_n N_A_1107_21#_c_1121_n 0.00163029f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_730 N_A_193_47#_c_900_n N_A_1107_21#_c_1130_n 0.00196084f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_731 N_A_193_47#_c_900_n N_A_1107_21#_c_1143_n 0.00348372f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_732 N_A_193_47#_c_900_n N_A_1107_21#_c_1122_n 0.00149139f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_733 N_A_193_47#_c_900_n N_A_1107_21#_c_1123_n 0.016449f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_734 N_A_193_47#_c_900_n N_A_1107_21#_c_1124_n 0.00917755f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_735 N_A_193_47#_c_900_n N_A_1107_21#_c_1132_n 8.24776e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_736 N_A_193_47#_c_900_n N_A_1107_21#_c_1148_n 6.83984e-19 $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_737 N_A_193_47#_c_894_n N_A_1107_21#_c_1125_n 0.0111636f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_738 N_A_193_47#_c_895_n N_A_1107_21#_c_1125_n 9.16922e-19 $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_739 N_A_193_47#_c_896_n N_A_1107_21#_c_1125_n 0.00462764f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_740 N_A_193_47#_c_900_n N_A_1107_21#_c_1125_n 0.0153364f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_741 N_A_193_47#_c_903_n N_A_1107_21#_c_1125_n 0.00129536f $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_742 N_A_193_47#_c_894_n N_A_1107_21#_c_1126_n 5.74798e-19 $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_743 N_A_193_47#_c_895_n N_A_1107_21#_c_1126_n 0.00181008f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_744 N_A_193_47#_c_896_n N_A_1107_21#_c_1126_n 0.00174717f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_745 N_A_193_47#_c_900_n N_A_1107_21#_c_1126_n 0.00365485f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_746 N_A_193_47#_c_903_n N_A_1107_21#_c_1126_n 6.8647e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_747 N_A_193_47#_c_900_n N_SET_B_c_1266_n 0.00391814f $X=8.365 $Y=1.19
+ $X2=-0.19 $Y2=-0.24
cc_748 N_A_193_47#_c_900_n N_SET_B_M1011_g 0.00116968f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_749 N_A_193_47#_c_900_n SET_B 0.00593372f $X=8.365 $Y=1.19 $X2=0 $Y2=0
cc_750 N_A_193_47#_c_894_n N_SET_B_c_1272_n 0.0194369f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_751 N_A_193_47#_c_895_n N_SET_B_c_1272_n 0.00227773f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_752 N_A_193_47#_c_896_n N_SET_B_c_1272_n 0.00534882f $X=8.937 $Y=1.305 $X2=0
+ $Y2=0
cc_753 N_A_193_47#_c_900_n N_SET_B_c_1272_n 0.158118f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_754 N_A_193_47#_c_903_n N_SET_B_c_1272_n 0.0254944f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_755 N_A_193_47#_c_900_n N_SET_B_c_1273_n 0.0265126f $X=8.365 $Y=1.19 $X2=0
+ $Y2=0
cc_756 N_A_193_47#_c_900_n N_A_931_47#_M1029_g 0.00190185f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_757 N_A_193_47#_M1041_g N_A_931_47#_c_1405_n 0.00264322f $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_758 N_A_193_47#_M1015_g N_A_931_47#_c_1411_n 0.00883573f $X=5.13 $Y=0.415
+ $X2=0 $Y2=0
cc_759 N_A_193_47#_c_897_n N_A_931_47#_c_1411_n 0.00579266f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_760 N_A_193_47#_c_902_n N_A_931_47#_c_1411_n 0.00257401f $X=5.29 $Y=0.85
+ $X2=0 $Y2=0
cc_761 N_A_193_47#_c_904_n N_A_931_47#_c_1411_n 5.24878e-19 $X=5.19 $Y=0.93
+ $X2=0 $Y2=0
cc_762 N_A_193_47#_c_905_n N_A_931_47#_c_1411_n 0.0194937f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_763 N_A_193_47#_M1041_g N_A_931_47#_c_1401_n 8.73767e-19 $X=4.59 $Y=2.275
+ $X2=0 $Y2=0
cc_764 N_A_193_47#_c_901_n N_A_931_47#_c_1401_n 3.03433e-19 $X=5.435 $Y=1.19
+ $X2=0 $Y2=0
cc_765 N_A_193_47#_M1015_g N_A_931_47#_c_1396_n 0.00119254f $X=5.13 $Y=0.415
+ $X2=0 $Y2=0
cc_766 N_A_193_47#_c_892_n N_A_931_47#_c_1396_n 8.54957e-19 $X=5.13 $Y=1.245
+ $X2=0 $Y2=0
cc_767 N_A_193_47#_c_900_n N_A_931_47#_c_1396_n 0.0145635f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_768 N_A_193_47#_c_902_n N_A_931_47#_c_1396_n 0.0138897f $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_769 N_A_193_47#_c_904_n N_A_931_47#_c_1396_n 7.78235e-19 $X=5.19 $Y=0.93
+ $X2=0 $Y2=0
cc_770 N_A_193_47#_c_905_n N_A_931_47#_c_1396_n 0.0244377f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_771 N_A_193_47#_c_900_n N_A_931_47#_c_1397_n 0.0379564f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_772 N_A_193_47#_c_892_n N_A_931_47#_c_1398_n 0.00268952f $X=5.13 $Y=1.245
+ $X2=0 $Y2=0
cc_773 N_A_193_47#_c_900_n N_A_931_47#_c_1398_n 0.0109965f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_774 N_A_193_47#_c_901_n N_A_931_47#_c_1398_n 0.00666557f $X=5.435 $Y=1.19
+ $X2=0 $Y2=0
cc_775 N_A_193_47#_c_904_n N_A_931_47#_c_1398_n 5.70846e-19 $X=5.19 $Y=0.93
+ $X2=0 $Y2=0
cc_776 N_A_193_47#_c_905_n N_A_931_47#_c_1398_n 0.0053097f $X=5.19 $Y=0.93 $X2=0
+ $Y2=0
cc_777 N_A_193_47#_c_900_n N_A_931_47#_c_1399_n 0.00390921f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_778 N_A_193_47#_c_900_n N_A_1400_21#_c_1501_n 0.00768602f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_779 N_A_193_47#_c_900_n N_A_1400_21#_c_1506_n 0.0122882f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_780 N_A_193_47#_c_896_n N_A_1400_21#_c_1515_n 0.00715591f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_781 N_A_193_47#_c_911_n N_A_1400_21#_c_1515_n 0.0157692f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_782 N_A_193_47#_c_912_n N_A_1400_21#_c_1515_n 0.00190553f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_783 N_A_193_47#_c_900_n N_A_1400_21#_c_1515_n 0.014133f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_784 N_A_193_47#_c_903_n N_A_1400_21#_c_1515_n 0.027417f $X=8.51 $Y=1.19 $X2=0
+ $Y2=0
cc_785 N_A_193_47#_c_900_n N_A_1400_21#_c_1516_n 0.0276968f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_786 N_A_193_47#_c_911_n N_A_1400_21#_c_1517_n 0.00264766f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_787 N_A_193_47#_c_900_n N_A_1400_21#_c_1517_n 0.00618009f $X=8.365 $Y=1.19
+ $X2=0 $Y2=0
cc_788 N_A_193_47#_c_911_n N_A_1887_21#_M1005_g 3.55913e-19 $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_789 N_A_193_47#_M1017_g N_A_1887_21#_M1042_g 0.0155835f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_790 N_A_193_47#_M1017_g N_A_1887_21#_c_1677_n 6.56548e-19 $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_791 N_A_193_47#_c_912_n N_A_1887_21#_c_1677_n 0.00900453f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_792 N_A_193_47#_M1017_g N_A_1714_47#_c_1852_n 0.00935459f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_793 N_A_193_47#_c_911_n N_A_1714_47#_c_1852_n 0.00669245f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_794 N_A_193_47#_c_912_n N_A_1714_47#_c_1852_n 0.0028948f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_795 N_A_193_47#_c_894_n N_A_1714_47#_c_1855_n 0.00390894f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_796 N_A_193_47#_c_895_n N_A_1714_47#_c_1855_n 0.00171906f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_797 N_A_193_47#_c_896_n N_A_1714_47#_c_1855_n 0.00314176f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_798 N_A_193_47#_c_894_n N_A_1714_47#_c_1841_n 0.011772f $X=8.615 $Y=0.87
+ $X2=0 $Y2=0
cc_799 N_A_193_47#_c_896_n N_A_1714_47#_c_1841_n 0.00837617f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_800 N_A_193_47#_c_903_n N_A_1714_47#_c_1841_n 6.65017e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_801 N_A_193_47#_M1017_g N_A_1714_47#_c_1847_n 0.00655842f $X=8.925 $Y=2.275
+ $X2=0 $Y2=0
cc_802 N_A_193_47#_c_911_n N_A_1714_47#_c_1847_n 0.0359925f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_803 N_A_193_47#_c_912_n N_A_1714_47#_c_1847_n 0.0021011f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_804 N_A_193_47#_c_896_n N_A_1714_47#_c_1843_n 0.00588727f $X=8.937 $Y=1.305
+ $X2=0 $Y2=0
cc_805 N_A_193_47#_c_911_n N_A_1714_47#_c_1843_n 0.00820582f $X=8.955 $Y=1.74
+ $X2=0 $Y2=0
cc_806 N_A_193_47#_c_903_n N_A_1714_47#_c_1843_n 2.68785e-19 $X=8.51 $Y=1.19
+ $X2=0 $Y2=0
cc_807 N_A_193_47#_c_906_n N_VPWR_c_2027_n 0.0127357f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_808 N_A_193_47#_c_906_n N_VPWR_c_2028_n 0.0391685f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_809 N_A_193_47#_c_906_n N_VPWR_c_2038_n 0.015988f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_810 N_A_193_47#_M1041_g N_VPWR_c_2040_n 0.00541732f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_811 N_A_193_47#_M1017_g N_VPWR_c_2041_n 0.00367119f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_812 N_A_193_47#_M1041_g N_VPWR_c_2026_n 0.00632491f $X=4.59 $Y=2.275 $X2=0
+ $Y2=0
cc_813 N_A_193_47#_M1017_g N_VPWR_c_2026_n 0.00567418f $X=8.925 $Y=2.275 $X2=0
+ $Y2=0
cc_814 N_A_193_47#_c_906_n N_VPWR_c_2026_n 0.00409094f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_815 N_A_193_47#_c_897_n N_A_453_363#_c_2238_n 0.0192415f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_816 N_A_193_47#_c_897_n N_A_453_363#_c_2239_n 0.00367673f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_817 N_A_193_47#_c_897_n N_A_453_363#_c_2240_n 0.00548406f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_818 N_A_193_47#_c_897_n N_A_453_363#_c_2241_n 0.0879477f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_819 N_A_193_47#_c_897_n N_A_453_363#_c_2242_n 0.0279145f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_820 N_A_193_47#_c_897_n N_A_453_363#_c_2243_n 0.00550979f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_821 N_A_193_47#_c_890_n N_A_453_363#_c_2244_n 0.00125006f $X=4.665 $Y=1.32
+ $X2=0 $Y2=0
cc_822 N_A_193_47#_c_897_n N_A_453_363#_c_2244_n 0.0256464f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_823 N_A_193_47#_c_890_n N_A_453_363#_c_2245_n 0.0156881f $X=4.665 $Y=1.32
+ $X2=0 $Y2=0
cc_824 N_A_193_47#_c_897_n N_A_453_363#_c_2245_n 0.0170158f $X=5.145 $Y=0.85
+ $X2=0 $Y2=0
cc_825 N_A_193_47#_c_905_n N_A_453_363#_c_2245_n 0.00205629f $X=5.19 $Y=0.93
+ $X2=0 $Y2=0
cc_826 N_A_193_47#_c_897_n N_VGND_c_2419_n 0.00411431f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_827 N_A_193_47#_c_906_n N_VGND_c_2419_n 0.0194875f $X=1.1 $Y=0.51 $X2=0 $Y2=0
cc_828 N_A_193_47#_c_897_n N_VGND_c_2420_n 0.00131319f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_829 N_A_193_47#_c_893_n N_VGND_c_2422_n 0.00175149f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_830 N_A_193_47#_M1015_g N_VGND_c_2426_n 0.00359964f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_831 N_A_193_47#_c_893_n N_VGND_c_2430_n 0.00435972f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_832 N_A_193_47#_c_894_n N_VGND_c_2430_n 0.00288727f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_833 N_A_193_47#_c_895_n N_VGND_c_2430_n 2.15978e-19 $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_834 N_A_193_47#_c_906_n N_VGND_c_2433_n 0.00978627f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_835 N_A_193_47#_M1027_d N_VGND_c_2438_n 0.00324958f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_836 N_A_193_47#_M1015_g N_VGND_c_2438_n 0.00564268f $X=5.13 $Y=0.415 $X2=0
+ $Y2=0
cc_837 N_A_193_47#_c_893_n N_VGND_c_2438_n 0.00616326f $X=8.495 $Y=0.705 $X2=0
+ $Y2=0
cc_838 N_A_193_47#_c_894_n N_VGND_c_2438_n 0.00224883f $X=8.615 $Y=0.87 $X2=0
+ $Y2=0
cc_839 N_A_193_47#_c_897_n N_VGND_c_2438_n 0.183568f $X=5.145 $Y=0.85 $X2=0
+ $Y2=0
cc_840 N_A_193_47#_c_898_n N_VGND_c_2438_n 0.0151383f $X=1.295 $Y=0.85 $X2=0
+ $Y2=0
cc_841 N_A_193_47#_c_902_n N_VGND_c_2438_n 0.0153531f $X=5.29 $Y=0.85 $X2=0
+ $Y2=0
cc_842 N_A_193_47#_c_906_n N_VGND_c_2438_n 0.00372614f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_843 N_A_193_47#_c_905_n A_1041_47# 0.00109904f $X=5.19 $Y=0.93 $X2=-0.19
+ $Y2=-0.24
cc_844 N_A_1107_21#_M1038_g N_SET_B_c_1266_n 0.0189927f $X=5.61 $Y=0.445
+ $X2=-0.19 $Y2=-0.24
cc_845 N_A_1107_21#_M1038_g N_SET_B_M1011_g 0.0137896f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_846 N_A_1107_21#_M1036_g N_SET_B_M1011_g 0.0101628f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_847 N_A_1107_21#_c_1130_n N_SET_B_M1011_g 0.0159332f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_848 N_A_1107_21#_c_1179_p N_SET_B_M1011_g 0.00507112f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_849 N_A_1107_21#_c_1132_n N_SET_B_M1011_g 0.00473578f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_850 N_A_1107_21#_c_1133_n N_SET_B_M1011_g 0.020182f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_851 N_A_1107_21#_M1038_g N_SET_B_M1044_g 0.0145491f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_852 N_A_1107_21#_c_1122_n N_SET_B_M1044_g 7.07383e-19 $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_853 N_A_1107_21#_M1038_g SET_B 0.00110276f $X=5.61 $Y=0.445 $X2=0 $Y2=0
cc_854 N_A_1107_21#_c_1122_n SET_B 0.00826425f $X=6.9 $Y=1.065 $X2=0 $Y2=0
cc_855 N_A_1107_21#_M1029_d N_SET_B_c_1272_n 5.47499e-19 $X=6.73 $Y=0.235 $X2=0
+ $Y2=0
cc_856 N_A_1107_21#_c_1121_n N_SET_B_c_1272_n 0.00505121f $X=8.015 $Y=0.985
+ $X2=0 $Y2=0
cc_857 N_A_1107_21#_c_1122_n N_SET_B_c_1272_n 0.0207654f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_858 N_A_1107_21#_c_1124_n N_SET_B_c_1272_n 0.0210775f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_859 N_A_1107_21#_c_1125_n N_SET_B_c_1272_n 0.0109336f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_860 N_A_1107_21#_c_1122_n N_SET_B_c_1273_n 0.0023059f $X=6.9 $Y=1.065 $X2=0
+ $Y2=0
cc_861 N_A_1107_21#_c_1122_n N_A_931_47#_M1029_g 0.00713446f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_862 N_A_1107_21#_c_1123_n N_A_931_47#_M1029_g 0.00191756f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_863 N_A_1107_21#_c_1143_n N_A_931_47#_M1037_g 0.0126258f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_864 N_A_1107_21#_M1036_g N_A_931_47#_c_1405_n 0.00191115f $X=5.61 $Y=2.275
+ $X2=0 $Y2=0
cc_865 N_A_1107_21#_M1038_g N_A_931_47#_c_1411_n 0.00853561f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_866 N_A_1107_21#_M1038_g N_A_931_47#_c_1401_n 0.0154362f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_867 N_A_1107_21#_c_1132_n N_A_931_47#_c_1401_n 0.0330453f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_868 N_A_1107_21#_M1038_g N_A_931_47#_c_1396_n 0.0188177f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_869 N_A_1107_21#_c_1130_n N_A_931_47#_c_1397_n 0.0141289f $X=6.385 $Y=1.91
+ $X2=0 $Y2=0
cc_870 N_A_1107_21#_c_1143_n N_A_931_47#_c_1397_n 0.00218253f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_871 N_A_1107_21#_c_1123_n N_A_931_47#_c_1397_n 0.0246731f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_872 N_A_1107_21#_c_1148_n N_A_931_47#_c_1397_n 0.00650509f $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_873 N_A_1107_21#_M1038_g N_A_931_47#_c_1398_n 0.0109165f $X=5.61 $Y=0.445
+ $X2=0 $Y2=0
cc_874 N_A_1107_21#_c_1132_n N_A_931_47#_c_1398_n 0.0169843f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_875 N_A_1107_21#_c_1133_n N_A_931_47#_c_1398_n 0.0011995f $X=5.72 $Y=1.74
+ $X2=0 $Y2=0
cc_876 N_A_1107_21#_c_1123_n N_A_931_47#_c_1399_n 0.00939619f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_877 N_A_1107_21#_c_1148_n N_A_931_47#_c_1399_n 9.09922e-19 $X=6.47 $Y=1.87
+ $X2=0 $Y2=0
cc_878 N_A_1107_21#_c_1122_n N_A_1400_21#_c_1500_n 0.0078099f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_879 N_A_1107_21#_c_1124_n N_A_1400_21#_c_1500_n 0.00387485f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_880 N_A_1107_21#_c_1122_n N_A_1400_21#_c_1501_n 0.00166514f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_881 N_A_1107_21#_c_1123_n N_A_1400_21#_c_1501_n 0.00752116f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_882 N_A_1107_21#_c_1124_n N_A_1400_21#_c_1501_n 0.0118467f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_883 N_A_1107_21#_c_1125_n N_A_1400_21#_c_1501_n 0.00205483f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_884 N_A_1107_21#_c_1126_n N_A_1400_21#_c_1501_n 0.0187813f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_885 N_A_1107_21#_M1047_g N_A_1400_21#_M1032_g 0.0153539f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_886 N_A_1107_21#_c_1143_n N_A_1400_21#_M1032_g 0.00219889f $X=6.815 $Y=1.91
+ $X2=0 $Y2=0
cc_887 N_A_1107_21#_M1047_g N_A_1400_21#_c_1506_n 2.86505e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_888 N_A_1107_21#_c_1123_n N_A_1400_21#_c_1506_n 0.0309286f $X=6.9 $Y=1.785
+ $X2=0 $Y2=0
cc_889 N_A_1107_21#_c_1124_n N_A_1400_21#_c_1506_n 0.0205152f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_890 N_A_1107_21#_c_1126_n N_A_1400_21#_c_1506_n 0.00382982f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_891 N_A_1107_21#_c_1125_n N_A_1400_21#_c_1516_n 9.59092e-19 $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_892 N_A_1107_21#_c_1126_n N_A_1400_21#_c_1516_n 0.00358318f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_893 N_A_1107_21#_M1047_g N_A_1400_21#_c_1517_n 0.0143059f $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_894 N_A_1107_21#_c_1124_n N_A_1400_21#_c_1517_n 0.00760725f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_895 N_A_1107_21#_c_1125_n N_A_1400_21#_c_1517_n 0.0207118f $X=7.96 $Y=0.98
+ $X2=0 $Y2=0
cc_896 N_A_1107_21#_c_1126_n N_A_1400_21#_c_1517_n 0.00632961f $X=7.96 $Y=1.15
+ $X2=0 $Y2=0
cc_897 N_A_1107_21#_M1047_g N_A_1714_47#_c_1852_n 7.04843e-19 $X=7.785 $Y=2.065
+ $X2=0 $Y2=0
cc_898 N_A_1107_21#_M1036_g N_VPWR_c_2030_n 0.00326498f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_899 N_A_1107_21#_c_1130_n N_VPWR_c_2030_n 0.0124698f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_900 N_A_1107_21#_c_1179_p N_VPWR_c_2030_n 0.00820313f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_901 N_A_1107_21#_c_1132_n N_VPWR_c_2030_n 0.0125544f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_902 N_A_1107_21#_c_1133_n N_VPWR_c_2030_n 7.62241e-19 $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_903 N_A_1107_21#_M1047_g N_VPWR_c_2031_n 0.0163458f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_904 N_A_1107_21#_c_1143_n N_VPWR_c_2031_n 0.0048929f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_905 N_A_1107_21#_c_1130_n N_VPWR_c_2033_n 0.00474052f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_906 N_A_1107_21#_c_1179_p N_VPWR_c_2033_n 0.00725778f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_907 N_A_1107_21#_c_1143_n N_VPWR_c_2033_n 0.00598455f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_908 N_A_1107_21#_M1036_g N_VPWR_c_2040_n 0.00535335f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_909 N_A_1107_21#_c_1132_n N_VPWR_c_2040_n 0.00111392f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_910 N_A_1107_21#_M1047_g N_VPWR_c_2041_n 0.00585385f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_911 N_A_1107_21#_M1011_d N_VPWR_c_2026_n 0.0031612f $X=6.215 $Y=2.065 $X2=0
+ $Y2=0
cc_912 N_A_1107_21#_M1036_g N_VPWR_c_2026_n 0.00664368f $X=5.61 $Y=2.275 $X2=0
+ $Y2=0
cc_913 N_A_1107_21#_M1047_g N_VPWR_c_2026_n 0.00762825f $X=7.785 $Y=2.065 $X2=0
+ $Y2=0
cc_914 N_A_1107_21#_c_1130_n N_VPWR_c_2026_n 0.00386836f $X=6.385 $Y=1.91 $X2=0
+ $Y2=0
cc_915 N_A_1107_21#_c_1179_p N_VPWR_c_2026_n 0.0029026f $X=6.47 $Y=2.21 $X2=0
+ $Y2=0
cc_916 N_A_1107_21#_c_1143_n N_VPWR_c_2026_n 0.00505387f $X=6.815 $Y=1.91 $X2=0
+ $Y2=0
cc_917 N_A_1107_21#_c_1132_n N_VPWR_c_2026_n 0.00128163f $X=5.72 $Y=1.74 $X2=0
+ $Y2=0
cc_918 N_A_1107_21#_c_1143_n A_1351_329# 0.00339576f $X=6.815 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_919 N_A_1107_21#_c_1123_n A_1351_329# 0.00178287f $X=6.9 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_920 N_A_1107_21#_M1038_g N_VGND_c_2421_n 0.00361232f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_921 N_A_1107_21#_c_1121_n N_VGND_c_2422_n 0.0114734f $X=8.015 $Y=0.985 $X2=0
+ $Y2=0
cc_922 N_A_1107_21#_c_1124_n N_VGND_c_2422_n 0.0040026f $X=7.795 $Y=0.98 $X2=0
+ $Y2=0
cc_923 N_A_1107_21#_c_1125_n N_VGND_c_2422_n 0.00376516f $X=7.96 $Y=0.98 $X2=0
+ $Y2=0
cc_924 N_A_1107_21#_c_1126_n N_VGND_c_2422_n 8.2379e-19 $X=7.96 $Y=1.15 $X2=0
+ $Y2=0
cc_925 N_A_1107_21#_M1038_g N_VGND_c_2426_n 0.0035977f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_926 N_A_1107_21#_c_1121_n N_VGND_c_2430_n 0.00447018f $X=8.015 $Y=0.985 $X2=0
+ $Y2=0
cc_927 N_A_1107_21#_M1029_d N_VGND_c_2438_n 0.00178362f $X=6.73 $Y=0.235 $X2=0
+ $Y2=0
cc_928 N_A_1107_21#_M1038_g N_VGND_c_2438_n 0.00580574f $X=5.61 $Y=0.445 $X2=0
+ $Y2=0
cc_929 N_A_1107_21#_c_1121_n N_VGND_c_2438_n 0.0044523f $X=8.015 $Y=0.985 $X2=0
+ $Y2=0
cc_930 N_A_1107_21#_M1029_d N_A_1251_47#_c_2632_n 0.0030477f $X=6.73 $Y=0.235
+ $X2=0 $Y2=0
cc_931 N_A_1107_21#_c_1122_n N_A_1251_47#_c_2632_n 0.0147335f $X=6.9 $Y=1.065
+ $X2=0 $Y2=0
cc_932 N_A_1107_21#_c_1124_n N_A_1251_47#_c_2632_n 0.00259503f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_933 N_A_1107_21#_c_1121_n N_A_1251_47#_c_2635_n 0.00462428f $X=8.015 $Y=0.985
+ $X2=0 $Y2=0
cc_934 N_A_1107_21#_c_1124_n N_A_1251_47#_c_2635_n 0.0122543f $X=7.795 $Y=0.98
+ $X2=0 $Y2=0
cc_935 N_SET_B_c_1266_n N_A_931_47#_M1029_g 0.00629904f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_936 N_SET_B_M1044_g N_A_931_47#_M1029_g 0.0205543f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_937 SET_B N_A_931_47#_M1029_g 0.00184456f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_938 N_SET_B_c_1272_n N_A_931_47#_M1029_g 0.0049202f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_939 N_SET_B_c_1273_n N_A_931_47#_M1029_g 0.00134438f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_940 N_SET_B_M1011_g N_A_931_47#_M1037_g 0.0228864f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_941 N_SET_B_c_1266_n N_A_931_47#_c_1396_n 0.00216489f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_942 N_SET_B_M1011_g N_A_931_47#_c_1396_n 6.04572e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_943 N_SET_B_M1044_g N_A_931_47#_c_1396_n 0.00182721f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_944 SET_B N_A_931_47#_c_1396_n 0.0244028f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_945 N_SET_B_c_1273_n N_A_931_47#_c_1396_n 0.00111115f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1266_n N_A_931_47#_c_1397_n 0.00310411f $X=6.14 $Y=1.145 $X2=0
+ $Y2=0
cc_947 N_SET_B_M1011_g N_A_931_47#_c_1397_n 0.0131452f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_948 SET_B N_A_931_47#_c_1397_n 0.0245807f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_949 N_SET_B_c_1272_n N_A_931_47#_c_1397_n 0.00369274f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_950 N_SET_B_c_1273_n N_A_931_47#_c_1397_n 6.67689e-19 $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_951 N_SET_B_M1011_g N_A_931_47#_c_1398_n 5.20457e-19 $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_952 N_SET_B_M1011_g N_A_931_47#_c_1399_n 0.021088f $X=6.14 $Y=2.275 $X2=0
+ $Y2=0
cc_953 N_SET_B_c_1272_n N_A_1400_21#_c_1500_n 0.00317213f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_954 N_SET_B_c_1272_n N_A_1400_21#_c_1506_n 5.29205e-19 $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_955 N_SET_B_M1008_g N_A_1400_21#_c_1515_n 0.00584134f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_956 N_SET_B_c_1272_n N_A_1400_21#_c_1515_n 0.0486626f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_957 N_SET_B_c_1274_n N_A_1400_21#_c_1515_n 0.0135087f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_958 N_SET_B_M1004_g N_A_1887_21#_M1005_g 0.015714f $X=10.055 $Y=0.445 $X2=0
+ $Y2=0
cc_959 N_SET_B_M1008_g N_A_1887_21#_M1005_g 0.0134226f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1272_n N_A_1887_21#_M1005_g 0.00634101f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_961 N_SET_B_c_1274_n N_A_1887_21#_M1005_g 0.00139314f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_962 N_SET_B_c_1275_n N_A_1887_21#_M1005_g 0.00233878f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1276_n N_A_1887_21#_M1005_g 0.0208839f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_964 N_SET_B_M1008_g N_A_1887_21#_M1042_g 0.0109753f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_965 N_SET_B_M1008_g N_A_1887_21#_c_1676_n 0.00710111f $X=10.055 $Y=2.275
+ $X2=0 $Y2=0
cc_966 N_SET_B_M1008_g N_A_1887_21#_c_1677_n 0.0197396f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_967 N_SET_B_M1008_g N_A_1887_21#_c_1678_n 0.0136222f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1275_n N_A_1887_21#_c_1667_n 0.00715913f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_969 N_SET_B_M1004_g N_A_1887_21#_c_1699_n 6.60782e-19 $X=10.055 $Y=0.445
+ $X2=0 $Y2=0
cc_970 N_SET_B_c_1274_n N_A_1887_21#_c_1699_n 4.23354e-19 $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_971 N_SET_B_c_1275_n N_A_1887_21#_c_1699_n 0.00228797f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_972 N_SET_B_M1004_g N_A_1714_47#_M1018_g 0.0242751f $X=10.055 $Y=0.445 $X2=0
+ $Y2=0
cc_973 N_SET_B_c_1275_n N_A_1714_47#_M1018_g 0.00127662f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_974 N_SET_B_M1008_g N_A_1714_47#_M1024_g 0.0325064f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_975 N_SET_B_c_1272_n N_A_1714_47#_c_1855_n 0.00885264f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1272_n N_A_1714_47#_c_1841_n 0.017797f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_977 N_SET_B_c_1274_n N_A_1714_47#_c_1841_n 0.0022902f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_978 N_SET_B_c_1275_n N_A_1714_47#_c_1841_n 0.0118231f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_979 N_SET_B_M1008_g N_A_1714_47#_c_1842_n 0.0117551f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_980 N_SET_B_c_1272_n N_A_1714_47#_c_1842_n 0.00876649f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_981 N_SET_B_c_1274_n N_A_1714_47#_c_1842_n 0.00124273f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1275_n N_A_1714_47#_c_1842_n 0.0248097f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1276_n N_A_1714_47#_c_1842_n 0.00455716f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1276_n N_A_1714_47#_c_1844_n 0.00111157f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_985 N_SET_B_c_1276_n N_A_1714_47#_c_1845_n 0.0212871f $X=9.93 $Y=0.98 $X2=0
+ $Y2=0
cc_986 N_SET_B_M1011_g N_VPWR_c_2030_n 0.0094739f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_987 N_SET_B_M1011_g N_VPWR_c_2033_n 0.00373914f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_988 N_SET_B_M1008_g N_VPWR_c_2036_n 0.00368415f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_989 N_SET_B_M1011_g N_VPWR_c_2026_n 0.00439789f $X=6.14 $Y=2.275 $X2=0 $Y2=0
cc_990 N_SET_B_M1008_g N_VPWR_c_2026_n 0.00444663f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_991 N_SET_B_M1008_g N_VPWR_c_2050_n 0.00857728f $X=10.055 $Y=2.275 $X2=0
+ $Y2=0
cc_992 N_SET_B_c_1272_n N_VGND_M1003_s 0.00213358f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_993 N_SET_B_c_1266_n N_VGND_c_2421_n 8.58768e-19 $X=6.14 $Y=1.145 $X2=0 $Y2=0
cc_994 N_SET_B_M1044_g N_VGND_c_2421_n 0.00289978f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_995 SET_B N_VGND_c_2421_n 0.010979f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_996 N_SET_B_c_1272_n N_VGND_c_2422_n 0.00409691f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_997 N_SET_B_M1004_g N_VGND_c_2423_n 0.00602618f $X=10.055 $Y=0.445 $X2=0
+ $Y2=0
cc_998 N_SET_B_c_1272_n N_VGND_c_2423_n 0.00606882f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_999 N_SET_B_c_1274_n N_VGND_c_2423_n 7.41662e-19 $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1000 N_SET_B_c_1275_n N_VGND_c_2423_n 0.00367619f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1001 N_SET_B_M1044_g N_VGND_c_2428_n 0.00422832f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_1002 SET_B N_VGND_c_2428_n 0.00221313f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1003 N_SET_B_M1004_g N_VGND_c_2435_n 0.00412007f $X=10.055 $Y=0.445 $X2=0
+ $Y2=0
cc_1004 N_SET_B_c_1275_n N_VGND_c_2435_n 0.00372651f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1005 N_SET_B_M1044_g N_VGND_c_2438_n 0.00586703f $X=6.18 $Y=0.445 $X2=0 $Y2=0
cc_1006 N_SET_B_M1004_g N_VGND_c_2438_n 0.00609966f $X=10.055 $Y=0.445 $X2=0
+ $Y2=0
cc_1007 SET_B N_VGND_c_2438_n 0.00214749f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1008 N_SET_B_c_1272_n N_VGND_c_2438_n 0.165394f $X=9.745 $Y=0.85 $X2=0 $Y2=0
cc_1009 N_SET_B_c_1273_n N_VGND_c_2438_n 0.014741f $X=6.355 $Y=0.85 $X2=0 $Y2=0
cc_1010 N_SET_B_c_1274_n N_VGND_c_2438_n 0.0143955f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1011 N_SET_B_c_1275_n N_VGND_c_2438_n 0.00251752f $X=9.89 $Y=0.85 $X2=0 $Y2=0
cc_1012 N_SET_B_c_1272_n N_A_1251_47#_M1044_d 0.00182819f $X=9.745 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1013 N_SET_B_c_1273_n N_A_1251_47#_M1044_d 6.80926e-19 $X=6.355 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1014 N_SET_B_c_1272_n N_A_1251_47#_M1028_d 0.0019616f $X=9.745 $Y=0.85 $X2=0
+ $Y2=0
cc_1015 N_SET_B_c_1272_n N_A_1251_47#_c_2632_n 0.00543044f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1016 N_SET_B_c_1272_n N_A_1251_47#_c_2635_n 0.00269828f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1017 N_SET_B_M1044_g N_A_1251_47#_c_2642_n 0.00296999f $X=6.18 $Y=0.445 $X2=0
+ $Y2=0
cc_1018 SET_B N_A_1251_47#_c_2642_n 0.00198247f $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_1019 N_SET_B_c_1272_n N_A_1251_47#_c_2642_n 0.00537146f $X=9.745 $Y=0.85
+ $X2=0 $Y2=0
cc_1020 N_SET_B_c_1273_n N_A_1251_47#_c_2642_n 0.0020226f $X=6.355 $Y=0.85 $X2=0
+ $Y2=0
cc_1021 N_SET_B_c_1272_n A_1618_47# 0.00371138f $X=9.745 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_1022 N_SET_B_M1004_g N_A_2026_47#_c_2662_n 0.00423086f $X=10.055 $Y=0.445
+ $X2=0 $Y2=0
cc_1023 N_SET_B_c_1275_n N_A_2026_47#_c_2662_n 0.0022235f $X=9.89 $Y=0.85 $X2=0
+ $Y2=0
cc_1024 N_A_931_47#_M1029_g N_A_1400_21#_c_1500_n 0.0282065f $X=6.655 $Y=0.555
+ $X2=0 $Y2=0
cc_1025 N_A_931_47#_M1029_g N_A_1400_21#_c_1501_n 0.00228862f $X=6.655 $Y=0.555
+ $X2=0 $Y2=0
cc_1026 N_A_931_47#_c_1399_n N_A_1400_21#_c_1501_n 0.0322452f $X=6.56 $Y=1.32
+ $X2=0 $Y2=0
cc_1027 N_A_931_47#_M1037_g N_A_1400_21#_M1032_g 0.0322452f $X=6.68 $Y=2.065
+ $X2=0 $Y2=0
cc_1028 N_A_931_47#_M1037_g N_VPWR_c_2030_n 0.00136797f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1029 N_A_931_47#_M1037_g N_VPWR_c_2033_n 0.00432313f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1030 N_A_931_47#_c_1405_n N_VPWR_c_2040_n 0.0377433f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1031 N_A_931_47#_M1041_d N_VPWR_c_2026_n 0.00173085f $X=4.665 $Y=2.065 $X2=0
+ $Y2=0
cc_1032 N_A_931_47#_M1037_g N_VPWR_c_2026_n 0.00600471f $X=6.68 $Y=2.065 $X2=0
+ $Y2=0
cc_1033 N_A_931_47#_c_1405_n N_VPWR_c_2026_n 0.0132511f $X=5.295 $Y=2.335 $X2=0
+ $Y2=0
cc_1034 N_A_931_47#_c_1405_n N_A_453_363#_c_2245_n 0.0128808f $X=5.295 $Y=2.335
+ $X2=0 $Y2=0
cc_1035 N_A_931_47#_c_1405_n A_1017_413# 0.00858887f $X=5.295 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1036 N_A_931_47#_c_1401_n A_1017_413# 0.00579571f $X=5.38 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1037 N_A_931_47#_c_1411_n N_VGND_c_2426_n 0.055608f $X=5.545 $Y=0.365 $X2=0
+ $Y2=0
cc_1038 N_A_931_47#_M1029_g N_VGND_c_2428_n 0.00357877f $X=6.655 $Y=0.555 $X2=0
+ $Y2=0
cc_1039 N_A_931_47#_M1043_d N_VGND_c_2438_n 0.00275359f $X=4.655 $Y=0.235 $X2=0
+ $Y2=0
cc_1040 N_A_931_47#_M1029_g N_VGND_c_2438_n 0.00535752f $X=6.655 $Y=0.555 $X2=0
+ $Y2=0
cc_1041 N_A_931_47#_c_1411_n N_VGND_c_2438_n 0.0218827f $X=5.545 $Y=0.365 $X2=0
+ $Y2=0
cc_1042 N_A_931_47#_c_1411_n A_1041_47# 0.00568226f $X=5.545 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1043 N_A_931_47#_M1029_g N_A_1251_47#_c_2632_n 0.00821062f $X=6.655 $Y=0.555
+ $X2=0 $Y2=0
cc_1044 N_A_931_47#_c_1399_n N_A_1251_47#_c_2642_n 0.00126312f $X=6.56 $Y=1.32
+ $X2=0 $Y2=0
cc_1045 N_A_1400_21#_c_1515_n N_A_1887_21#_M1005_g 0.00413877f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1046 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1676_n 0.015309f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1047 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1677_n 0.0070058f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1048 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1678_n 0.010417f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1049 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1706_n 0.00964432f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1050 N_A_1400_21#_M1030_g N_A_1887_21#_c_1667_n 0.012752f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1051 N_A_1400_21#_M1031_g N_A_1887_21#_c_1667_n 0.0057985f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1052 N_A_1400_21#_c_1504_n N_A_1887_21#_c_1667_n 0.00591558f $X=11.355
+ $Y=0.84 $X2=0 $Y2=0
cc_1053 N_A_1400_21#_c_1512_n N_A_1887_21#_c_1667_n 0.0127165f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1054 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1667_n 0.0265111f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1055 N_A_1400_21#_c_1518_n N_A_1887_21#_c_1667_n 5.59542e-19 $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1056 N_A_1400_21#_c_1507_n N_A_1887_21#_c_1667_n 0.00911985f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1057 N_A_1400_21#_c_1508_n N_A_1887_21#_c_1667_n 0.044948f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1058 N_A_1400_21#_M1006_s N_A_1887_21#_c_1680_n 0.00479715f $X=11.555
+ $Y=1.505 $X2=0 $Y2=0
cc_1059 N_A_1400_21#_M1030_g N_A_1887_21#_c_1680_n 0.00741003f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1060 N_A_1400_21#_c_1512_n N_A_1887_21#_c_1680_n 0.0212381f $X=11.355 $Y=1.66
+ $X2=0 $Y2=0
cc_1061 N_A_1400_21#_c_1513_n N_A_1887_21#_c_1680_n 0.0321071f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1062 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1680_n 0.00664652f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1063 N_A_1400_21#_c_1518_n N_A_1887_21#_c_1680_n 0.00170504f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1064 N_A_1400_21#_c_1507_n N_A_1887_21#_c_1680_n 0.00265268f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1065 N_A_1400_21#_c_1513_n N_A_1887_21#_c_1681_n 0.00840283f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1066 N_A_1400_21#_c_1515_n N_A_1887_21#_c_1723_n 0.00453864f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1067 N_A_1400_21#_M1031_g N_A_1887_21#_c_1699_n 0.00365275f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1068 N_A_1400_21#_c_1505_n N_A_1887_21#_c_1699_n 0.00292314f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1069 N_A_1400_21#_M1030_g N_A_1887_21#_c_1726_n 0.00480312f $X=10.895
+ $Y=2.065 $X2=0 $Y2=0
cc_1070 N_A_1400_21#_M1031_g N_A_1714_47#_M1018_g 0.0294176f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1071 N_A_1400_21#_M1030_g N_A_1714_47#_M1024_g 0.039703f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1072 N_A_1400_21#_c_1515_n N_A_1714_47#_M1024_g 0.00711753f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1073 N_A_1400_21#_c_1515_n N_A_1714_47#_c_1847_n 0.0219541f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1074 N_A_1400_21#_c_1515_n N_A_1714_47#_c_1842_n 0.0228784f $X=11.125 $Y=1.53
+ $X2=0 $Y2=0
cc_1075 N_A_1400_21#_M1031_g N_A_1714_47#_c_1844_n 2.38141e-19 $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1076 N_A_1400_21#_c_1515_n N_A_1714_47#_c_1844_n 0.00714757f $X=11.125
+ $Y=1.53 $X2=0 $Y2=0
cc_1077 N_A_1400_21#_M1031_g N_A_1714_47#_c_1845_n 0.0117459f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1078 N_A_1400_21#_c_1507_n N_A_1714_47#_c_1845_n 0.039703f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1079 N_A_1400_21#_c_1503_n N_RESET_B_M1013_g 0.00680862f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1080 N_A_1400_21#_c_1505_n N_RESET_B_M1013_g 0.00288669f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1081 N_A_1400_21#_c_1508_n N_RESET_B_M1013_g 0.00237866f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1082 N_A_1400_21#_c_1513_n N_RESET_B_M1006_g 0.00360287f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1083 N_A_1400_21#_c_1518_n N_RESET_B_M1006_g 0.00264823f $X=11.27 $Y=1.53
+ $X2=0 $Y2=0
cc_1084 N_A_1400_21#_c_1507_n N_RESET_B_M1006_g 0.0025096f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1085 N_A_1400_21#_c_1508_n N_RESET_B_M1006_g 0.00309824f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1086 N_A_1400_21#_c_1503_n RESET_B 0.0186919f $X=11.565 $Y=0.84 $X2=0 $Y2=0
cc_1087 N_A_1400_21#_c_1513_n RESET_B 0.015564f $X=11.68 $Y=1.66 $X2=0 $Y2=0
cc_1088 N_A_1400_21#_c_1507_n RESET_B 5.50348e-19 $X=10.95 $Y=1.32 $X2=0 $Y2=0
cc_1089 N_A_1400_21#_c_1508_n RESET_B 0.0185145f $X=11.165 $Y=1.32 $X2=0 $Y2=0
cc_1090 N_A_1400_21#_M1031_g N_RESET_B_c_1940_n 0.00201274f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1091 N_A_1400_21#_c_1503_n N_RESET_B_c_1940_n 0.00512123f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1092 N_A_1400_21#_c_1513_n N_RESET_B_c_1940_n 0.00527649f $X=11.68 $Y=1.66
+ $X2=0 $Y2=0
cc_1093 N_A_1400_21#_c_1507_n N_RESET_B_c_1940_n 0.0092343f $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1094 N_A_1400_21#_c_1508_n N_RESET_B_c_1940_n 0.00327697f $X=11.165 $Y=1.32
+ $X2=0 $Y2=0
cc_1095 N_A_1400_21#_c_1506_n N_VPWR_M1032_d 0.00297048f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1096 N_A_1400_21#_c_1517_n N_VPWR_M1032_d 0.00221014f $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1097 N_A_1400_21#_c_1512_n N_VPWR_M1030_d 0.00314302f $X=11.355 $Y=1.66 $X2=0
+ $Y2=0
cc_1098 N_A_1400_21#_c_1501_n N_VPWR_c_2031_n 0.00111411f $X=7.1 $Y=1.485 $X2=0
+ $Y2=0
cc_1099 N_A_1400_21#_M1032_g N_VPWR_c_2031_n 0.00353361f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1100 N_A_1400_21#_c_1506_n N_VPWR_c_2031_n 0.011531f $X=7.32 $Y=1.32 $X2=0
+ $Y2=0
cc_1101 N_A_1400_21#_c_1517_n N_VPWR_c_2031_n 7.83548e-19 $X=8.05 $Y=1.53 $X2=0
+ $Y2=0
cc_1102 N_A_1400_21#_M1032_g N_VPWR_c_2033_n 0.00583607f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1103 N_A_1400_21#_M1030_g N_VPWR_c_2035_n 0.0111257f $X=10.895 $Y=2.065 $X2=0
+ $Y2=0
cc_1104 N_A_1400_21#_M1030_g N_VPWR_c_2036_n 0.00339283f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1105 N_A_1400_21#_M1032_g N_VPWR_c_2026_n 0.00670824f $X=7.1 $Y=2.065 $X2=0
+ $Y2=0
cc_1106 N_A_1400_21#_M1030_g N_VPWR_c_2026_n 0.00383548f $X=10.895 $Y=2.065
+ $X2=0 $Y2=0
cc_1107 N_A_1400_21#_c_1517_n A_1572_329# 0.00272182f $X=8.05 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1108 N_A_1400_21#_c_1500_n N_VGND_c_2422_n 0.00315399f $X=7.075 $Y=0.95 $X2=0
+ $Y2=0
cc_1109 N_A_1400_21#_c_1503_n N_VGND_c_2424_n 0.00352079f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1110 N_A_1400_21#_c_1505_n N_VGND_c_2424_n 0.00629548f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1111 N_A_1400_21#_c_1500_n N_VGND_c_2428_n 0.00357877f $X=7.075 $Y=0.95 $X2=0
+ $Y2=0
cc_1112 N_A_1400_21#_M1031_g N_VGND_c_2435_n 0.00357877f $X=10.95 $Y=0.555 $X2=0
+ $Y2=0
cc_1113 N_A_1400_21#_c_1503_n N_VGND_c_2435_n 0.00300947f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1114 N_A_1400_21#_c_1504_n N_VGND_c_2435_n 0.00167376f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1115 N_A_1400_21#_c_1505_n N_VGND_c_2435_n 0.0128605f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1116 N_A_1400_21#_M1013_s N_VGND_c_2438_n 0.00387761f $X=11.555 $Y=0.235
+ $X2=0 $Y2=0
cc_1117 N_A_1400_21#_c_1500_n N_VGND_c_2438_n 0.00661646f $X=7.075 $Y=0.95 $X2=0
+ $Y2=0
cc_1118 N_A_1400_21#_M1031_g N_VGND_c_2438_n 0.00657041f $X=10.95 $Y=0.555 $X2=0
+ $Y2=0
cc_1119 N_A_1400_21#_c_1503_n N_VGND_c_2438_n 0.00541125f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1120 N_A_1400_21#_c_1504_n N_VGND_c_2438_n 0.00326613f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1121 N_A_1400_21#_c_1505_n N_VGND_c_2438_n 0.0075831f $X=11.68 $Y=0.43 $X2=0
+ $Y2=0
cc_1122 N_A_1400_21#_c_1500_n N_A_1251_47#_c_2632_n 0.0105921f $X=7.075 $Y=0.95
+ $X2=0 $Y2=0
cc_1123 N_A_1400_21#_c_1504_n N_A_2026_47#_M1031_d 0.00388496f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1124 N_A_1400_21#_M1031_g N_A_2026_47#_c_2665_n 0.0112584f $X=10.95 $Y=0.555
+ $X2=0 $Y2=0
cc_1125 N_A_1400_21#_c_1504_n N_A_2026_47#_c_2665_n 0.0138009f $X=11.355 $Y=0.84
+ $X2=0 $Y2=0
cc_1126 N_A_1400_21#_c_1505_n N_A_2026_47#_c_2665_n 0.0149851f $X=11.68 $Y=0.43
+ $X2=0 $Y2=0
cc_1127 N_A_1400_21#_c_1507_n N_A_2026_47#_c_2665_n 5.45076e-19 $X=10.95 $Y=1.32
+ $X2=0 $Y2=0
cc_1128 N_A_1887_21#_c_1667_n N_A_1714_47#_M1018_g 0.00267624f $X=10.817
+ $Y=1.915 $X2=0 $Y2=0
cc_1129 N_A_1887_21#_c_1699_n N_A_1714_47#_M1018_g 0.00474602f $X=10.74 $Y=0.73
+ $X2=0 $Y2=0
cc_1130 N_A_1887_21#_c_1706_n N_A_1714_47#_M1024_g 0.0118664f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1131 N_A_1887_21#_M1042_g N_A_1714_47#_c_1852_n 0.00204127f $X=9.515 $Y=2.275
+ $X2=0 $Y2=0
cc_1132 N_A_1887_21#_M1005_g N_A_1714_47#_c_1841_n 0.0101965f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1133 N_A_1887_21#_M1005_g N_A_1714_47#_c_1847_n 0.00912509f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1134 N_A_1887_21#_M1042_g N_A_1714_47#_c_1847_n 0.0058046f $X=9.515 $Y=2.275
+ $X2=0 $Y2=0
cc_1135 N_A_1887_21#_c_1676_n N_A_1714_47#_c_1847_n 0.0248025f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1136 N_A_1887_21#_c_1735_p N_A_1714_47#_c_1847_n 0.0135579f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1137 N_A_1887_21#_M1005_g N_A_1714_47#_c_1842_n 0.0115262f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_1138 N_A_1887_21#_c_1676_n N_A_1714_47#_c_1842_n 0.0154989f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1139 N_A_1887_21#_c_1677_n N_A_1714_47#_c_1842_n 0.00130368f $X=9.635 $Y=1.74
+ $X2=0 $Y2=0
cc_1140 N_A_1887_21#_c_1678_n N_A_1714_47#_c_1842_n 0.00635717f $X=10.24 $Y=2
+ $X2=0 $Y2=0
cc_1141 N_A_1887_21#_c_1723_n N_A_1714_47#_c_1842_n 0.00162703f $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1142 N_A_1887_21#_c_1706_n N_A_1714_47#_c_1844_n 0.00158774f $X=10.73 $Y=2
+ $X2=0 $Y2=0
cc_1143 N_A_1887_21#_c_1667_n N_A_1714_47#_c_1844_n 0.0241086f $X=10.817
+ $Y=1.915 $X2=0 $Y2=0
cc_1144 N_A_1887_21#_c_1723_n N_A_1714_47#_c_1844_n 9.97507e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1145 N_A_1887_21#_c_1667_n N_A_1714_47#_c_1845_n 0.0123488f $X=10.817
+ $Y=1.915 $X2=0 $Y2=0
cc_1146 N_A_1887_21#_c_1723_n N_A_1714_47#_c_1845_n 4.0151e-19 $X=10.325 $Y=2
+ $X2=0 $Y2=0
cc_1147 N_A_1887_21#_c_1659_n N_RESET_B_M1013_g 0.0182169f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1148 N_A_1887_21#_c_1661_n N_RESET_B_M1013_g 0.0180063f $X=12.475 $Y=1.16
+ $X2=0 $Y2=0
cc_1149 N_A_1887_21#_c_1668_n N_RESET_B_M1013_g 0.00220565f $X=12.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1150 N_A_1887_21#_c_1680_n N_RESET_B_M1006_g 0.0142369f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1151 N_A_1887_21#_c_1661_n RESET_B 7.2676e-19 $X=12.475 $Y=1.16 $X2=0 $Y2=0
cc_1152 N_A_1887_21#_c_1680_n RESET_B 0.00314679f $X=12.16 $Y=2 $X2=0 $Y2=0
cc_1153 N_A_1887_21#_c_1668_n RESET_B 0.0193193f $X=12.34 $Y=1.16 $X2=0 $Y2=0
cc_1154 N_A_1887_21#_M1039_g N_RESET_B_c_1940_n 0.0294485f $X=12.375 $Y=1.985
+ $X2=0 $Y2=0
cc_1155 N_A_1887_21#_c_1681_n N_RESET_B_c_1940_n 0.00991514f $X=12.245 $Y=1.915
+ $X2=0 $Y2=0
cc_1156 N_A_1887_21#_c_1668_n N_RESET_B_c_1940_n 6.95467e-19 $X=12.34 $Y=1.16
+ $X2=0 $Y2=0
cc_1157 N_A_1887_21#_c_1663_n N_A_2596_47#_M1002_g 0.0046261f $X=13.19 $Y=1.535
+ $X2=0 $Y2=0
cc_1158 N_A_1887_21#_c_1675_n N_A_2596_47#_M1002_g 0.0111957f $X=13.315 $Y=1.61
+ $X2=0 $Y2=0
cc_1159 N_A_1887_21#_c_1659_n N_A_2596_47#_c_1974_n 0.00110305f $X=12.375
+ $Y=0.995 $X2=0 $Y2=0
cc_1160 N_A_1887_21#_c_1662_n N_A_2596_47#_c_1974_n 0.00388761f $X=13.19
+ $Y=1.025 $X2=0 $Y2=0
cc_1161 N_A_1887_21#_c_1664_n N_A_2596_47#_c_1974_n 0.00984702f $X=13.315
+ $Y=0.73 $X2=0 $Y2=0
cc_1162 N_A_1887_21#_c_1665_n N_A_2596_47#_c_1974_n 0.00979941f $X=13.315
+ $Y=0.805 $X2=0 $Y2=0
cc_1163 N_A_1887_21#_M1039_g N_A_2596_47#_c_1980_n 0.00166592f $X=12.375
+ $Y=1.985 $X2=0 $Y2=0
cc_1164 N_A_1887_21#_c_1663_n N_A_2596_47#_c_1980_n 0.00715595f $X=13.19
+ $Y=1.535 $X2=0 $Y2=0
cc_1165 N_A_1887_21#_c_1674_n N_A_2596_47#_c_1980_n 0.0107587f $X=13.315
+ $Y=1.685 $X2=0 $Y2=0
cc_1166 N_A_1887_21#_c_1675_n N_A_2596_47#_c_1980_n 0.0101477f $X=13.315 $Y=1.61
+ $X2=0 $Y2=0
cc_1167 N_A_1887_21#_c_1665_n N_A_2596_47#_c_1975_n 0.00368279f $X=13.315
+ $Y=0.805 $X2=0 $Y2=0
cc_1168 N_A_1887_21#_c_1675_n N_A_2596_47#_c_1975_n 0.00324612f $X=13.315
+ $Y=1.61 $X2=0 $Y2=0
cc_1169 N_A_1887_21#_c_1662_n N_A_2596_47#_c_1976_n 0.0131382f $X=13.19 $Y=1.025
+ $X2=0 $Y2=0
cc_1170 N_A_1887_21#_c_1660_n N_A_2596_47#_c_1977_n 0.0154274f $X=13.115 $Y=1.16
+ $X2=0 $Y2=0
cc_1171 N_A_1887_21#_c_1662_n N_A_2596_47#_c_1977_n 0.00115562f $X=13.19
+ $Y=1.025 $X2=0 $Y2=0
cc_1172 N_A_1887_21#_c_1663_n N_A_2596_47#_c_1977_n 0.00115562f $X=13.19
+ $Y=1.535 $X2=0 $Y2=0
cc_1173 N_A_1887_21#_c_1666_n N_A_2596_47#_c_1977_n 0.00732445f $X=13.19 $Y=1.16
+ $X2=0 $Y2=0
cc_1174 N_A_1887_21#_c_1662_n N_A_2596_47#_c_1978_n 0.0025256f $X=13.19 $Y=1.025
+ $X2=0 $Y2=0
cc_1175 N_A_1887_21#_c_1664_n N_A_2596_47#_c_1978_n 0.0159526f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1176 N_A_1887_21#_c_1678_n N_VPWR_M1042_d 0.00124767f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1177 N_A_1887_21#_c_1735_p N_VPWR_M1042_d 0.00160397f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1178 N_A_1887_21#_c_1680_n N_VPWR_M1030_d 0.0044189f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1179 N_A_1887_21#_c_1680_n N_VPWR_M1006_d 0.00750664f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1180 N_A_1887_21#_c_1681_n N_VPWR_M1006_d 0.00487804f $X=12.245 $Y=1.915
+ $X2=0 $Y2=0
cc_1181 N_A_1887_21#_c_1674_n N_VPWR_c_2032_n 0.00446435f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1182 N_A_1887_21#_c_1680_n N_VPWR_c_2035_n 0.0844105f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1183 N_A_1887_21#_c_1678_n N_VPWR_c_2036_n 0.00359839f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1184 N_A_1887_21#_c_1783_p N_VPWR_c_2036_n 0.00713694f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1185 N_A_1887_21#_c_1706_n N_VPWR_c_2036_n 0.00458994f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1186 N_A_1887_21#_c_1680_n N_VPWR_c_2036_n 5.56361e-19 $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1187 N_A_1887_21#_c_1726_n N_VPWR_c_2036_n 0.00270619f $X=10.817 $Y=2 $X2=0
+ $Y2=0
cc_1188 N_A_1887_21#_M1042_g N_VPWR_c_2041_n 0.00542601f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1189 N_A_1887_21#_c_1735_p N_VPWR_c_2041_n 9.91118e-19 $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1190 N_A_1887_21#_M1039_g N_VPWR_c_2043_n 0.0046653f $X=12.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1191 N_A_1887_21#_c_1674_n N_VPWR_c_2043_n 0.00464873f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1192 N_A_1887_21#_M1008_d N_VPWR_c_2026_n 0.00327257f $X=10.13 $Y=2.065 $X2=0
+ $Y2=0
cc_1193 N_A_1887_21#_M1042_g N_VPWR_c_2026_n 0.00997697f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1194 N_A_1887_21#_M1039_g N_VPWR_c_2026_n 0.00929621f $X=12.375 $Y=1.985
+ $X2=0 $Y2=0
cc_1195 N_A_1887_21#_c_1674_n N_VPWR_c_2026_n 0.00922843f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1196 N_A_1887_21#_c_1678_n N_VPWR_c_2026_n 0.00704318f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1197 N_A_1887_21#_c_1735_p N_VPWR_c_2026_n 0.00270501f $X=9.8 $Y=2 $X2=0
+ $Y2=0
cc_1198 N_A_1887_21#_c_1783_p N_VPWR_c_2026_n 0.00608739f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1199 N_A_1887_21#_c_1706_n N_VPWR_c_2026_n 0.00829558f $X=10.73 $Y=2 $X2=0
+ $Y2=0
cc_1200 N_A_1887_21#_c_1680_n N_VPWR_c_2026_n 0.00701098f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1201 N_A_1887_21#_c_1726_n N_VPWR_c_2026_n 0.00481592f $X=10.817 $Y=2 $X2=0
+ $Y2=0
cc_1202 N_A_1887_21#_M1042_g N_VPWR_c_2050_n 0.00321606f $X=9.515 $Y=2.275 $X2=0
+ $Y2=0
cc_1203 N_A_1887_21#_c_1677_n N_VPWR_c_2050_n 7.01948e-19 $X=9.635 $Y=1.74 $X2=0
+ $Y2=0
cc_1204 N_A_1887_21#_c_1678_n N_VPWR_c_2050_n 0.0106677f $X=10.24 $Y=2 $X2=0
+ $Y2=0
cc_1205 N_A_1887_21#_c_1735_p N_VPWR_c_2050_n 0.0126362f $X=9.8 $Y=2 $X2=0 $Y2=0
cc_1206 N_A_1887_21#_c_1783_p N_VPWR_c_2050_n 0.00687131f $X=10.325 $Y=2.21
+ $X2=0 $Y2=0
cc_1207 N_A_1887_21#_M1039_g N_VPWR_c_2051_n 0.0100464f $X=12.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1208 N_A_1887_21#_c_1680_n N_VPWR_c_2051_n 0.00915613f $X=12.16 $Y=2 $X2=0
+ $Y2=0
cc_1209 N_A_1887_21#_c_1706_n A_2122_329# 0.00202121f $X=10.73 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1210 N_A_1887_21#_c_1667_n A_2122_329# 0.0030402f $X=10.817 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1211 N_A_1887_21#_c_1726_n A_2122_329# 5.84995e-19 $X=10.817 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1212 N_A_1887_21#_c_1660_n N_Q_N_c_2374_n 0.00367611f $X=13.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1213 N_A_1887_21#_c_1674_n N_Q_N_c_2374_n 0.00131217f $X=13.315 $Y=1.685
+ $X2=0 $Y2=0
cc_1214 N_A_1887_21#_c_1675_n N_Q_N_c_2374_n 5.75727e-19 $X=13.315 $Y=1.61 $X2=0
+ $Y2=0
cc_1215 N_A_1887_21#_c_1659_n N_Q_N_c_2371_n 0.0051543f $X=12.375 $Y=0.995 $X2=0
+ $Y2=0
cc_1216 N_A_1887_21#_M1039_g N_Q_N_c_2371_n 0.00269981f $X=12.375 $Y=1.985 $X2=0
+ $Y2=0
cc_1217 N_A_1887_21#_c_1660_n N_Q_N_c_2371_n 0.0206846f $X=13.115 $Y=1.16 $X2=0
+ $Y2=0
cc_1218 N_A_1887_21#_c_1661_n N_Q_N_c_2371_n 6.7688e-19 $X=12.475 $Y=1.16 $X2=0
+ $Y2=0
cc_1219 N_A_1887_21#_c_1663_n N_Q_N_c_2371_n 5.75727e-19 $X=13.19 $Y=1.535 $X2=0
+ $Y2=0
cc_1220 N_A_1887_21#_c_1665_n N_Q_N_c_2371_n 8.62582e-19 $X=13.315 $Y=0.805
+ $X2=0 $Y2=0
cc_1221 N_A_1887_21#_c_1681_n N_Q_N_c_2371_n 0.0126467f $X=12.245 $Y=1.915 $X2=0
+ $Y2=0
cc_1222 N_A_1887_21#_c_1668_n N_Q_N_c_2371_n 0.0224114f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1223 N_A_1887_21#_c_1660_n Q_N 0.00357569f $X=13.115 $Y=1.16 $X2=0 $Y2=0
cc_1224 N_A_1887_21#_c_1674_n Q_N 8.69219e-19 $X=13.315 $Y=1.685 $X2=0 $Y2=0
cc_1225 N_A_1887_21#_c_1664_n N_Q_N_c_2373_n 0.00104845f $X=13.315 $Y=0.73 $X2=0
+ $Y2=0
cc_1226 N_A_1887_21#_M1005_g N_VGND_c_2423_n 0.00844839f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1227 N_A_1887_21#_c_1659_n N_VGND_c_2424_n 0.0127745f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1228 N_A_1887_21#_c_1661_n N_VGND_c_2424_n 0.00200592f $X=12.475 $Y=1.16
+ $X2=0 $Y2=0
cc_1229 N_A_1887_21#_c_1668_n N_VGND_c_2424_n 0.0105198f $X=12.34 $Y=1.16 $X2=0
+ $Y2=0
cc_1230 N_A_1887_21#_c_1664_n N_VGND_c_2425_n 0.00415965f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1231 N_A_1887_21#_M1005_g N_VGND_c_2430_n 0.00486043f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1232 N_A_1887_21#_c_1659_n N_VGND_c_2436_n 0.0046653f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1233 N_A_1887_21#_c_1664_n N_VGND_c_2436_n 0.00533769f $X=13.315 $Y=0.73
+ $X2=0 $Y2=0
cc_1234 N_A_1887_21#_c_1665_n N_VGND_c_2436_n 2.84936e-19 $X=13.315 $Y=0.805
+ $X2=0 $Y2=0
cc_1235 N_A_1887_21#_M1018_d N_VGND_c_2438_n 0.00216833f $X=10.605 $Y=0.235
+ $X2=0 $Y2=0
cc_1236 N_A_1887_21#_M1005_g N_VGND_c_2438_n 0.00476342f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_1237 N_A_1887_21#_c_1659_n N_VGND_c_2438_n 0.00934473f $X=12.375 $Y=0.995
+ $X2=0 $Y2=0
cc_1238 N_A_1887_21#_c_1664_n N_VGND_c_2438_n 0.0109269f $X=13.315 $Y=0.73 $X2=0
+ $Y2=0
cc_1239 N_A_1887_21#_M1018_d N_A_2026_47#_c_2665_n 0.00332514f $X=10.605
+ $Y=0.235 $X2=0 $Y2=0
cc_1240 N_A_1887_21#_c_1699_n N_A_2026_47#_c_2665_n 0.0115748f $X=10.74 $Y=0.73
+ $X2=0 $Y2=0
cc_1241 N_A_1714_47#_M1024_g N_VPWR_c_2035_n 0.00209073f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1242 N_A_1714_47#_M1024_g N_VPWR_c_2036_n 0.00425094f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1243 N_A_1714_47#_c_1852_n N_VPWR_c_2041_n 0.0377433f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1244 N_A_1714_47#_M1033_d N_VPWR_c_2026_n 0.00205544f $X=8.58 $Y=2.065 $X2=0
+ $Y2=0
cc_1245 N_A_1714_47#_M1024_g N_VPWR_c_2026_n 0.00591666f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1246 N_A_1714_47#_c_1852_n N_VPWR_c_2026_n 0.0272797f $X=9.21 $Y=2.335 $X2=0
+ $Y2=0
cc_1247 N_A_1714_47#_M1024_g N_VPWR_c_2050_n 0.00144209f $X=10.535 $Y=2.065
+ $X2=0 $Y2=0
cc_1248 N_A_1714_47#_c_1852_n A_1800_413# 0.0111731f $X=9.21 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1249 N_A_1714_47#_c_1847_n A_1800_413# 0.00577347f $X=9.295 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1250 N_A_1714_47#_c_1855_n N_VGND_c_2430_n 0.0433004f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1251 N_A_1714_47#_M1018_g N_VGND_c_2435_n 0.00357877f $X=10.53 $Y=0.555 $X2=0
+ $Y2=0
cc_1252 N_A_1714_47#_M1009_d N_VGND_c_2438_n 0.00269406f $X=8.57 $Y=0.235 $X2=0
+ $Y2=0
cc_1253 N_A_1714_47#_M1018_g N_VGND_c_2438_n 0.00541008f $X=10.53 $Y=0.555 $X2=0
+ $Y2=0
cc_1254 N_A_1714_47#_c_1855_n N_VGND_c_2438_n 0.0129075f $X=9.21 $Y=0.365 $X2=0
+ $Y2=0
cc_1255 N_A_1714_47#_c_1855_n A_1822_47# 0.00370882f $X=9.21 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1256 N_A_1714_47#_c_1841_n A_1822_47# 0.00307731f $X=9.295 $Y=1.235 $X2=-0.19
+ $Y2=-0.24
cc_1257 N_A_1714_47#_M1018_g N_A_2026_47#_c_2665_n 0.00964551f $X=10.53 $Y=0.555
+ $X2=0 $Y2=0
cc_1258 N_A_1714_47#_c_1844_n N_A_2026_47#_c_2665_n 0.00273006f $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1259 N_A_1714_47#_c_1844_n N_A_2026_47#_c_2662_n 0.001984f $X=10.475 $Y=1.24
+ $X2=0 $Y2=0
cc_1260 N_A_1714_47#_c_1845_n N_A_2026_47#_c_2662_n 3.56528e-19 $X=10.475
+ $Y=1.24 $X2=0 $Y2=0
cc_1261 N_RESET_B_M1006_g N_VPWR_c_2042_n 0.00655753f $X=11.89 $Y=1.825 $X2=0
+ $Y2=0
cc_1262 N_RESET_B_M1013_g N_VGND_c_2424_n 0.00665319f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1263 N_RESET_B_M1013_g N_VGND_c_2435_n 0.00585385f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1264 N_RESET_B_M1013_g N_VGND_c_2438_n 0.0120869f $X=11.89 $Y=0.445 $X2=0
+ $Y2=0
cc_1265 N_A_2596_47#_M1002_g N_VPWR_c_2032_n 0.0147323f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1266 N_A_2596_47#_c_1980_n N_VPWR_c_2032_n 0.048761f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1267 N_A_2596_47#_c_1975_n N_VPWR_c_2032_n 0.010763f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1268 N_A_2596_47#_c_1976_n N_VPWR_c_2032_n 0.00249491f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1269 N_A_2596_47#_c_1980_n N_VPWR_c_2043_n 0.0169293f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1270 N_A_2596_47#_M1002_g N_VPWR_c_2044_n 0.0046653f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1271 N_A_2596_47#_M1002_g N_VPWR_c_2026_n 0.00895857f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1272 N_A_2596_47#_c_1980_n N_VPWR_c_2026_n 0.0115924f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1273 N_A_2596_47#_c_1980_n N_Q_N_c_2371_n 0.0871059f $X=13.105 $Y=1.91 $X2=0
+ $Y2=0
cc_1274 N_A_2596_47#_c_1977_n N_Q_N_c_2371_n 0.0251545f $X=13.117 $Y=1.16 $X2=0
+ $Y2=0
cc_1275 N_A_2596_47#_c_1974_n N_Q_N_c_2373_n 0.0590331f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1276 N_A_2596_47#_M1002_g N_Q_c_2403_n 0.0105677f $X=13.79 $Y=1.985 $X2=0
+ $Y2=0
cc_1277 N_A_2596_47#_c_1975_n N_Q_c_2403_n 0.0266143f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1278 N_A_2596_47#_c_1976_n N_Q_c_2403_n 0.00804901f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1279 N_A_2596_47#_c_1978_n N_Q_c_2403_n 0.00640119f $X=13.725 $Y=0.995 $X2=0
+ $Y2=0
cc_1280 N_A_2596_47#_c_1974_n N_VGND_c_2425_n 0.0212529f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1281 N_A_2596_47#_c_1975_n N_VGND_c_2425_n 0.0103062f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1282 N_A_2596_47#_c_1976_n N_VGND_c_2425_n 0.00246314f $X=13.71 $Y=1.16 $X2=0
+ $Y2=0
cc_1283 N_A_2596_47#_c_1978_n N_VGND_c_2425_n 0.00939953f $X=13.725 $Y=0.995
+ $X2=0 $Y2=0
cc_1284 N_A_2596_47#_c_1974_n N_VGND_c_2436_n 0.0199778f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1285 N_A_2596_47#_c_1978_n N_VGND_c_2437_n 0.0046653f $X=13.725 $Y=0.995
+ $X2=0 $Y2=0
cc_1286 N_A_2596_47#_M1046_s N_VGND_c_2438_n 0.00210122f $X=12.98 $Y=0.235 $X2=0
+ $Y2=0
cc_1287 N_A_2596_47#_c_1974_n N_VGND_c_2438_n 0.0118987f $X=13.105 $Y=0.51 $X2=0
+ $Y2=0
cc_1288 N_A_2596_47#_c_1978_n N_VGND_c_2438_n 0.00895857f $X=13.725 $Y=0.995
+ $X2=0 $Y2=0
cc_1289 N_VPWR_c_2026_n N_A_453_363#_M1014_d 0.00306969f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1290 N_VPWR_c_2028_n N_A_453_363#_c_2246_n 0.0161853f $X=1.62 $Y=1.97 $X2=0
+ $Y2=0
cc_1291 N_VPWR_c_2039_n N_A_453_363#_c_2246_n 0.0138534f $X=3.31 $Y=2.72 $X2=0
+ $Y2=0
cc_1292 N_VPWR_c_2026_n N_A_453_363#_c_2246_n 0.00564495f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1293 N_VPWR_c_2040_n N_A_453_363#_c_2245_n 0.0154725f $X=5.705 $Y=2.72 $X2=0
+ $Y2=0
cc_1294 N_VPWR_c_2026_n N_A_453_363#_c_2245_n 0.00409094f $X=14.03 $Y=2.72 $X2=0
+ $Y2=0
cc_1295 N_VPWR_c_2026_n A_752_413# 0.00238611f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1296 N_VPWR_c_2026_n A_1017_413# 0.00355877f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1297 N_VPWR_c_2026_n A_1351_329# 0.0026811f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1298 N_VPWR_c_2026_n A_1572_329# 0.00777501f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1299 N_VPWR_c_2026_n A_1800_413# 0.00555699f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1300 N_VPWR_c_2026_n A_2122_329# 0.00245111f $X=14.03 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1301 N_VPWR_c_2026_n N_Q_N_M1039_d 0.00387172f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1302 N_VPWR_c_2032_n Q_N 0.00155557f $X=13.58 $Y=1.94 $X2=0 $Y2=0
cc_1303 N_VPWR_c_2043_n Q_N 0.0197934f $X=13.45 $Y=2.72 $X2=0 $Y2=0
cc_1304 N_VPWR_c_2026_n Q_N 0.0108988f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1305 N_VPWR_c_2026_n N_Q_M1002_d 0.00387172f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1306 N_VPWR_c_2044_n Q 0.018001f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1307 N_VPWR_c_2026_n Q 0.00993603f $X=14.03 $Y=2.72 $X2=0 $Y2=0
cc_1308 N_A_453_363#_c_2245_n N_VGND_c_2426_n 0.0115451f $X=4.315 $Y=0.47 $X2=0
+ $Y2=0
cc_1309 N_A_453_363#_c_2239_n N_VGND_c_2434_n 0.0254287f $X=2.67 $Y=0.43 $X2=0
+ $Y2=0
cc_1310 N_A_453_363#_M1022_d N_VGND_c_2438_n 0.00195871f $X=2.295 $Y=0.235 $X2=0
+ $Y2=0
cc_1311 N_A_453_363#_M1023_d N_VGND_c_2438_n 0.00295839f $X=4.18 $Y=0.235 $X2=0
+ $Y2=0
cc_1312 N_A_453_363#_c_2239_n N_VGND_c_2438_n 0.0070926f $X=2.67 $Y=0.43 $X2=0
+ $Y2=0
cc_1313 N_A_453_363#_c_2245_n N_VGND_c_2438_n 0.00398697f $X=4.315 $Y=0.47 $X2=0
+ $Y2=0
cc_1314 N_Q_N_c_2371_n N_VGND_c_2424_n 0.00205006f $X=12.642 $Y=1.63 $X2=0 $Y2=0
cc_1315 N_Q_N_c_2373_n N_VGND_c_2436_n 0.0196011f $X=12.642 $Y=0.573 $X2=0 $Y2=0
cc_1316 N_Q_N_M1001_d N_VGND_c_2438_n 0.00387172f $X=12.45 $Y=0.235 $X2=0 $Y2=0
cc_1317 N_Q_N_c_2373_n N_VGND_c_2438_n 0.010859f $X=12.642 $Y=0.573 $X2=0 $Y2=0
cc_1318 Q N_VGND_c_2437_n 0.0179623f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1319 N_Q_M1016_d N_VGND_c_2438_n 0.00387172f $X=13.865 $Y=0.235 $X2=0 $Y2=0
cc_1320 Q N_VGND_c_2438_n 0.00992739f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1321 N_VGND_c_2438_n A_381_47# 0.00204609f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1322 N_VGND_c_2438_n A_764_47# 0.00302076f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1323 N_VGND_c_2438_n A_1041_47# 0.0022723f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1324 N_VGND_c_2438_n N_A_1251_47#_M1044_d 0.00211076f $X=14.03 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1325 N_VGND_c_2438_n N_A_1251_47#_M1028_d 0.00184756f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1326 N_VGND_c_2422_n N_A_1251_47#_c_2632_n 0.0113334f $X=7.805 $Y=0.38 $X2=0
+ $Y2=0
cc_1327 N_VGND_c_2428_n N_A_1251_47#_c_2632_n 0.0131017f $X=7.64 $Y=0 $X2=0
+ $Y2=0
cc_1328 N_VGND_c_2438_n N_A_1251_47#_c_2632_n 0.00350344f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1329 N_VGND_c_2422_n N_A_1251_47#_c_2635_n 0.00239801f $X=7.805 $Y=0.38 $X2=0
+ $Y2=0
cc_1330 N_VGND_c_2428_n N_A_1251_47#_c_2642_n 0.0535339f $X=7.64 $Y=0 $X2=0
+ $Y2=0
cc_1331 N_VGND_c_2438_n N_A_1251_47#_c_2642_n 0.0158341f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1332 N_VGND_c_2438_n A_1618_47# 0.00474691f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1333 N_VGND_c_2438_n A_1822_47# 0.00257693f $X=14.03 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1334 N_VGND_c_2438_n N_A_2026_47#_M1004_d 0.00259397f $X=14.03 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1335 N_VGND_c_2438_n N_A_2026_47#_M1031_d 0.00224765f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1336 N_VGND_c_2435_n N_A_2026_47#_c_2665_n 0.0113648f $X=12 $Y=0 $X2=0 $Y2=0
cc_1337 N_VGND_c_2438_n N_A_2026_47#_c_2665_n 0.00654393f $X=14.03 $Y=0 $X2=0
+ $Y2=0
cc_1338 N_VGND_c_2423_n N_A_2026_47#_c_2662_n 0.0120194f $X=9.735 $Y=0.36 $X2=0
+ $Y2=0
cc_1339 N_VGND_c_2435_n N_A_2026_47#_c_2662_n 0.0547553f $X=12 $Y=0 $X2=0 $Y2=0
cc_1340 N_VGND_c_2438_n N_A_2026_47#_c_2662_n 0.0353125f $X=14.03 $Y=0 $X2=0
+ $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.075000 0.875000 1.275000 ;
        RECT 0.705000 1.275000 0.875000 1.445000 ;
        RECT 0.705000 1.445000 1.880000 1.615000 ;
        RECT 1.710000 1.075000 3.230000 1.275000 ;
        RECT 1.710000 1.275000 1.880000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.075000 1.540000 1.275000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.420000 1.075000 4.090000 1.275000 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.005000 1.075000 1.295000 1.120000 ;
        RECT 1.005000 1.120000 4.055000 1.260000 ;
        RECT 1.005000 1.260000 1.295000 1.305000 ;
        RECT 3.765000 1.075000 4.055000 1.120000 ;
        RECT 3.765000 1.260000 4.055000 1.305000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.656750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.625000 0.645000 3.955000 0.725000 ;
        RECT 3.625000 0.725000 5.895000 0.905000 ;
        RECT 4.985000 0.645000 5.315000 0.725000 ;
        RECT 5.025000 1.415000 5.895000 1.625000 ;
        RECT 5.025000 1.625000 5.275000 2.125000 ;
        RECT 5.485000 0.905000 5.895000 1.415000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.190000  0.085000 0.360000 0.555000 ;
        RECT 1.030000  0.085000 1.200000 0.555000 ;
        RECT 1.870000  0.085000 2.040000 0.555000 ;
        RECT 2.810000  0.085000 2.980000 0.555000 ;
        RECT 4.645000  0.085000 4.815000 0.555000 ;
        RECT 5.485000  0.085000 5.655000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.570000 2.135000 0.820000 2.635000 ;
        RECT 2.770000 2.135000 3.020000 2.635000 ;
        RECT 3.610000 2.135000 3.915000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.120000 0.725000 1.700000 0.905000 ;
      RECT 0.120000 0.905000 0.290000 1.785000 ;
      RECT 0.120000 1.785000 2.220000 1.955000 ;
      RECT 0.120000 2.135000 0.400000 2.465000 ;
      RECT 0.145000 2.125000 0.315000 2.135000 ;
      RECT 0.530000 0.255000 0.860000 0.725000 ;
      RECT 0.990000 2.135000 1.240000 2.295000 ;
      RECT 0.990000 2.295000 2.080000 2.465000 ;
      RECT 1.065000 2.125000 1.235000 2.135000 ;
      RECT 1.370000 0.255000 1.700000 0.725000 ;
      RECT 1.410000 1.955000 1.660000 2.125000 ;
      RECT 1.830000 2.135000 2.080000 2.295000 ;
      RECT 2.050000 1.445000 4.785000 1.615000 ;
      RECT 2.050000 1.615000 2.220000 1.785000 ;
      RECT 2.285000 2.125000 2.600000 2.465000 ;
      RECT 2.310000 0.255000 2.640000 0.725000 ;
      RECT 2.310000 0.725000 3.400000 0.905000 ;
      RECT 2.390000 1.785000 4.855000 1.955000 ;
      RECT 2.390000 1.955000 2.600000 2.125000 ;
      RECT 3.150000 0.255000 4.380000 0.475000 ;
      RECT 3.150000 0.475000 3.400000 0.725000 ;
      RECT 3.190000 1.955000 3.440000 2.465000 ;
      RECT 4.085000 1.955000 4.855000 2.295000 ;
      RECT 4.085000 2.295000 5.695000 2.465000 ;
      RECT 4.615000 1.075000 5.275000 1.245000 ;
      RECT 4.615000 1.245000 4.785000 1.445000 ;
      RECT 5.445000 1.795000 5.695000 2.295000 ;
    LAYER mcon ;
      RECT 0.145000 2.125000 0.315000 2.295000 ;
      RECT 1.065000 2.125000 1.235000 2.295000 ;
    LAYER met1 ;
      RECT 0.085000 2.095000 0.375000 2.140000 ;
      RECT 0.085000 2.140000 1.295000 2.280000 ;
      RECT 0.085000 2.280000 0.375000 2.325000 ;
      RECT 1.005000 2.095000 1.295000 2.140000 ;
      RECT 1.005000 2.280000 1.295000 2.325000 ;
  END
END sky130_fd_sc_hd__xor2_2
END LIBRARY

* File: sky130_fd_sc_hd__a221o_1.spice
* Created: Thu Aug 27 14:01:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a221o_1.pex.spice"
.subckt sky130_fd_sc_hd__a221o_1  VNB VPB C1 B2 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_C1_M1011_g N_A_27_47#_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1006 A_205_47# N_B2_M1006_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.10725 PD=0.86 PS=0.98 NRD=9.228 NRS=10.152 M=1 R=4.33333 SA=75000.7
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1007_d N_B1_M1007_g A_205_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.06825 PD=1.82 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_465_47# N_A1_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=20.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_465_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.102375 AS=0.10725 PD=0.965 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_A_27_47#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.102375 PD=1.82 PS=0.965 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_109_297#_M1008_d N_C1_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1001 N_A_193_297#_M1001_d N_B2_M1001_g N_A_109_297#_M1008_d VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_109_297#_M1000_d N_B1_M1000_g N_A_193_297#_M1001_d VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_193_297#_M1010_d N_A1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.26 PD=1.33 PS=2.52 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_193_297#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1575 AS=0.165 PD=1.315 PS=1.33 NRD=7.8603 NRS=5.8903 M=1 R=6.66667
+ SA=75000.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.1575 PD=2.52 PS=1.315 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a221o_1.pxi.spice"
*
.ends
*
*

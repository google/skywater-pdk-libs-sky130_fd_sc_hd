* File: sky130_fd_sc_hd__a21o_4.spice
* Created: Tue Sep  1 18:52:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21o_4.pex.spice"
.subckt sky130_fd_sc_hd__a21o_4  VNB VPB B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_84_21#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.091 PD=1.87 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_A_84_21#_M1003_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1003_d N_A_84_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_84_21#_M1014_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.264875 AS=0.091 PD=1.465 PS=0.93 NRD=20.304 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_84_21#_M1007_d N_B1_M1007_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.264875 PD=0.92 PS=1.465 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75002.5 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1010 N_A_84_21#_M1007_d N_B1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10075 PD=0.92 PS=0.96 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75002.9
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1009 A_901_47# N_A2_M1009_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65 AD=0.07475
+ AS=0.10075 PD=0.88 PS=0.96 NRD=11.076 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1006 N_A_84_21#_M1006_d N_A1_M1006_g A_901_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.07475 PD=0.92 PS=0.88 NRD=0 NRS=11.076 M=1 R=4.33333
+ SA=75003.7 SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_A_84_21#_M1006_d N_A1_M1008_g A_741_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75004.1
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 A_741_47# N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.169 PD=0.92 PS=1.82 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75004.6 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_84_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_X_M1002_d N_A_84_21#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1011 N_X_M1011_d N_A_84_21#_M1011_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1015 N_X_M1011_d N_A_84_21#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1017 N_A_483_297#_M1017_d N_B1_M1017_g N_A_84_21#_M1017_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1019 N_A_483_297#_M1019_d N_B1_M1019_g N_A_84_21#_M1017_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_483_297#_M1019_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_483_297#_M1000_d N_A1_M1000_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.2 A=0.15 P=2.3 MULT=1
MM1018 N_A_483_297#_M1000_d N_A1_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1018_s N_A2_M1013_g N_A_483_297#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.395 PD=1.27 PS=2.79 NRD=0 NRS=25.5903 M=1 R=6.66667 SA=75002.3
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=9.4695 P=15.01
*
.include "sky130_fd_sc_hd__a21o_4.pxi.spice"
*
.ends
*
*

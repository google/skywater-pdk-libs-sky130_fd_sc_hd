* File: sky130_fd_sc_hd__nand4b_2.spice.pex
* Created: Thu Aug 27 14:30:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND4B_2%A_N 3 7 9 10 17
r29 14 17 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.47 $Y2=1.16
r30 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.16 $X2=0.21
+ $Y2=1.53
r31 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r32 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r33 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r34 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r35 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%A_27_47# 1 2 7 9 12 14 16 19 23 27 30 32 35
+ 40 44 46 50
c88 14 0 1.05021e-19 $X=1.83 $Y=0.995
r89 49 50 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16
+ $X2=1.83 $Y2=1.16
r90 36 49 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.215 $Y=1.16
+ $X2=1.41 $Y2=1.16
r91 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r92 33 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.16
+ $X2=0.585 $Y2=1.16
r93 33 35 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.67 $Y=1.16
+ $X2=1.215 $Y2=1.16
r94 32 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=1.915
+ $X2=0.585 $Y2=2
r95 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=1.245
+ $X2=0.585 $Y2=1.16
r96 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.585 $Y=1.245
+ $X2=0.585 $Y2=1.915
r97 30 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=1.075
+ $X2=0.585 $Y2=1.16
r98 29 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=0.72
r99 29 30 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.585 $Y=0.805
+ $X2=0.585 $Y2=1.075
r100 25 44 24.0086 $w=1.68e-07 $l=3.68e-07 $layer=LI1_cond $X=0.217 $Y=2
+ $X2=0.585 $Y2=2
r101 25 27 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.217 $Y=2.085
+ $X2=0.217 $Y2=2.29
r102 21 40 24.0086 $w=1.68e-07 $l=3.68e-07 $layer=LI1_cond $X=0.217 $Y=0.72
+ $X2=0.585 $Y2=0.72
r103 21 23 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.43
r104 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.16
r105 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.325
+ $X2=1.83 $Y2=1.985
r106 14 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=1.16
r107 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.995
+ $X2=1.83 $Y2=0.56
r108 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r109 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.985
r110 7 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r111 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r112 2 27 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.29
r113 1 23 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%B 1 3 6 8 10 13 15 16 17 25
c49 1 0 1.51188e-19 $X=2.25 $Y=0.995
r50 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.865
+ $Y=1.16 $X2=2.865 $Y2=1.16
r51 23 25 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.865 $Y2=1.16
r52 21 23 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.67 $Y2=1.16
r53 17 26 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=2.865 $Y2=1.175
r54 16 26 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=2.555 $Y=1.175
+ $X2=2.865 $Y2=1.175
r55 15 16 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.095 $Y=1.175
+ $X2=2.555 $Y2=1.175
r56 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.16
r57 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.985
r58 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r59 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=0.56
r60 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.325
+ $X2=2.25 $Y2=1.16
r61 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.25 $Y=1.325 $X2=2.25
+ $Y2=1.985
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.995
+ $X2=2.25 $Y2=1.16
r63 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.25 $Y=0.995 $X2=2.25
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%C 3 5 7 10 12 14 15 16 17 28
c47 28 0 1.17704e-19 $X=4.03 $Y=1.16
r48 26 28 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.02 $Y=1.16 $X2=4.03
+ $Y2=1.16
r49 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.02
+ $Y=1.16 $X2=4.02 $Y2=1.16
r50 24 26 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.98 $Y=1.16 $X2=4.02
+ $Y2=1.16
r51 23 24 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=3.61 $Y=1.16
+ $X2=3.98 $Y2=1.16
r52 21 23 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.56 $Y=1.16 $X2=3.61
+ $Y2=1.16
r53 17 27 19.1318 $w=1.98e-07 $l=3.45e-07 $layer=LI1_cond $X=4.365 $Y=1.175
+ $X2=4.02 $Y2=1.175
r54 16 27 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=4.02 $Y2=1.175
r55 15 16 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.445 $Y=1.175
+ $X2=3.905 $Y2=1.175
r56 12 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=1.16
r57 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.03 $Y=0.995
+ $X2=4.03 $Y2=0.56
r58 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.98 $Y=1.325
+ $X2=3.98 $Y2=1.16
r59 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.98 $Y=1.325
+ $X2=3.98 $Y2=1.985
r60 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.61 $Y=0.995
+ $X2=3.61 $Y2=1.16
r61 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.61 $Y=0.995 $X2=3.61
+ $Y2=0.56
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.325
+ $X2=3.56 $Y2=1.16
r63 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.56 $Y=1.325 $X2=3.56
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%D 3 5 7 10 12 14 15 16 22
c40 16 0 1.17704e-19 $X=5.285 $Y=1.19
r41 22 24 42.3981 $w=3.24e-07 $l=2.85e-07 $layer=POLY_cond $X=4.96 $Y=1.16
+ $X2=5.245 $Y2=1.16
r42 21 22 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=4.91 $Y=1.16 $X2=4.96
+ $Y2=1.16
r43 20 21 55.0432 $w=3.24e-07 $l=3.7e-07 $layer=POLY_cond $X=4.54 $Y=1.16
+ $X2=4.91 $Y2=1.16
r44 19 20 7.43827 $w=3.24e-07 $l=5e-08 $layer=POLY_cond $X=4.49 $Y=1.16 $X2=4.54
+ $Y2=1.16
r45 16 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.245
+ $Y=1.16 $X2=5.245 $Y2=1.16
r46 15 16 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=4.825 $Y=1.175
+ $X2=5.245 $Y2=1.175
r47 12 22 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=0.995
+ $X2=4.96 $Y2=1.16
r48 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.96 $Y=0.995
+ $X2=4.96 $Y2=0.56
r49 8 21 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=1.325
+ $X2=4.91 $Y2=1.16
r50 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.91 $Y=1.325
+ $X2=4.91 $Y2=1.985
r51 5 20 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=0.995
+ $X2=4.54 $Y2=1.16
r52 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.54 $Y=0.995 $X2=4.54
+ $Y2=0.56
r53 1 19 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.49 $Y=1.325
+ $X2=4.49 $Y2=1.16
r54 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.49 $Y=1.325 $X2=4.49
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%VPWR 1 2 3 4 5 6 21 25 29 33 35 37 42 43 45
+ 46 47 58 66 72 78 80 84
r78 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 77 78 8.96211 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.16 $Y=2.53
+ $X2=1.285 $Y2=2.53
r81 74 77 0.217469 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=1.15 $Y=2.53 $X2=1.16
+ $Y2=2.53
r82 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 71 74 10.221 $w=5.48e-07 $l=4.7e-07 $layer=LI1_cond $X=0.68 $Y=2.53 $X2=1.15
+ $Y2=2.53
r84 71 72 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=2.53
+ $X2=0.515 $Y2=2.53
r85 69 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r86 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r87 66 83 5.41725 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=5.277 $Y2=2.72
r88 66 68 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=4.83 $Y2=2.72
r89 65 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 65 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r91 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r92 62 80 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=3.435 $Y=2.72
+ $X2=3.115 $Y2=2.72
r93 62 64 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.435 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 61 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r95 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r96 58 80 13.0174 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.115 $Y2=2.72
r97 58 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 57 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r99 57 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r100 56 78 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.285 $Y2=2.72
r101 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r102 51 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r103 47 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r104 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r105 45 64 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 45 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.235 $Y2=2.72
r107 44 68 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.365 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 44 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.365 $Y=2.72
+ $X2=4.235 $Y2=2.72
r109 42 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r110 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.04 $Y2=2.72
r111 41 60 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.53 $Y2=2.72
r112 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.04 $Y2=2.72
r113 37 40 19.8395 $w=3.93e-07 $l=6.8e-07 $layer=LI1_cond $X=5.232 $Y=1.66
+ $X2=5.232 $Y2=2.34
r114 35 83 2.91009 $w=3.95e-07 $l=1.05119e-07 $layer=LI1_cond $X=5.232 $Y=2.635
+ $X2=5.277 $Y2=2.72
r115 35 40 8.60685 $w=3.93e-07 $l=2.95e-07 $layer=LI1_cond $X=5.232 $Y=2.635
+ $X2=5.232 $Y2=2.34
r116 31 46 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.235 $Y=2.635
+ $X2=4.235 $Y2=2.72
r117 31 33 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=4.235 $Y=2.635
+ $X2=4.235 $Y2=2
r118 27 80 2.66764 $w=6.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=2.635
+ $X2=3.115 $Y2=2.72
r119 27 29 11.8673 $w=6.38e-07 $l=6.35e-07 $layer=LI1_cond $X=3.115 $Y=2.635
+ $X2=3.115 $Y2=2
r120 23 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r121 23 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2
r122 19 77 5.37178 $w=2.5e-07 $l=2.75e-07 $layer=LI1_cond $X=1.16 $Y=2.255
+ $X2=1.16 $Y2=2.53
r123 19 21 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.16 $Y=2.255
+ $X2=1.16 $Y2=1.66
r124 6 40 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.485 $X2=5.2 $Y2=2.34
r125 6 37 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.485 $X2=5.2 $Y2=1.66
r126 5 33 300 $w=1.7e-07 $l=5.93949e-07 $layer=licon1_PDIFF $count=2 $X=4.055
+ $Y=1.485 $X2=4.225 $Y2=2
r127 4 29 150 $w=1.7e-07 $l=7.38918e-07 $layer=licon1_PDIFF $count=4 $X=2.745
+ $Y=1.485 $X2=3.27 $Y2=2
r128 3 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
r129 2 77 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.34
r130 2 21 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.66
r131 1 71 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%Y 1 2 3 4 5 18 20 24 26 30 32 36 39 41 42
+ 43 44 53
c83 42 0 1.51188e-19 $X=1.55 $Y=0.765
c84 32 0 1.59237e-19 $X=4.535 $Y=1.555
r85 53 61 1.226 $w=2.33e-07 $l=2.5e-08 $layer=LI1_cond $X=1.667 $Y=0.85
+ $X2=1.667 $Y2=0.825
r86 43 44 9.2696 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=1.667 $Y=1.19
+ $X2=1.667 $Y2=1.445
r87 42 61 4.63843 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.62 $Y=0.72
+ $X2=1.62 $Y2=0.825
r88 42 43 15.2024 $w=2.33e-07 $l=3.1e-07 $layer=LI1_cond $X=1.667 $Y=0.88
+ $X2=1.667 $Y2=1.19
r89 42 53 1.4712 $w=2.33e-07 $l=3e-08 $layer=LI1_cond $X=1.667 $Y=0.88 $X2=1.667
+ $Y2=0.85
r90 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.7 $Y=1.665 $X2=4.7
+ $Y2=2
r91 33 41 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=1.555
+ $X2=3.77 $Y2=1.555
r92 32 34 7.17723 $w=2.2e-07 $l=2.13014e-07 $layer=LI1_cond $X=4.535 $Y=1.555
+ $X2=4.7 $Y2=1.665
r93 32 33 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=4.535 $Y=1.555
+ $X2=3.935 $Y2=1.555
r94 28 41 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.77 $Y=1.665
+ $X2=3.77 $Y2=1.555
r95 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.77 $Y=1.665
+ $X2=3.77 $Y2=2.34
r96 27 39 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=1.555
+ $X2=2.46 $Y2=1.555
r97 26 41 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=1.555
+ $X2=3.77 $Y2=1.555
r98 26 27 51.3361 $w=2.18e-07 $l=9.8e-07 $layer=LI1_cond $X=3.605 $Y=1.555
+ $X2=2.625 $Y2=1.555
r99 22 39 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.46 $Y=1.665
+ $X2=2.46 $Y2=1.555
r100 22 24 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.46 $Y=1.665
+ $X2=2.46 $Y2=2.34
r101 21 44 2.25663 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.555
+ $X2=1.62 $Y2=1.555
r102 20 39 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=2.46 $Y2=1.555
r103 20 21 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=1.785 $Y2=1.555
r104 16 44 4.1757 $w=2.82e-07 $l=1.1e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.555
r105 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2.34
r106 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.565
+ $Y=1.485 $X2=4.7 $Y2=2
r107 4 41 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.485 $X2=3.77 $Y2=1.66
r108 4 30 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.485 $X2=3.77 $Y2=2.34
r109 3 39 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.66
r110 3 24 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.34
r111 2 44 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.66
r112 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2.34
r113 1 42 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%VGND 1 2 9 13 16 17 18 20 33 34 37
r68 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r70 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r71 30 31 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r72 28 31 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.37
+ $Y2=0
r73 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r74 27 30 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.37
+ $Y2=0
r75 27 28 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r76 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r77 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r78 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r79 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r80 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r81 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r82 16 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.37
+ $Y2=0
r83 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.75
+ $Y2=0
r84 15 33 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5.29
+ $Y2=0
r85 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.75
+ $Y2=0
r86 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0
r87 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0.38
r88 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r89 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r90 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.235 $X2=4.75 $Y2=0.38
r91 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%A_215_47# 1 2 3 10 12 14 20 22
r40 20 22 32.2257 $w=2.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.125 $Y=0.77
+ $X2=2.88 $Y2=0.77
r41 17 20 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.125 $Y2=0.77
r42 17 19 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.55
r43 16 19 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.465
+ $X2=2.04 $Y2=0.55
r44 15 25 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=1.16 $Y2=0.36
r45 14 16 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.955 $Y=0.36
+ $X2=2.04 $Y2=0.465
r46 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=0.36
+ $X2=1.285 $Y2=0.36
r47 10 25 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.36
r48 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.72
r49 3 22 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.72
r50 2 19 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.55
r51 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
r52 1 12 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%A_465_47# 1 2 11
c16 11 0 1.05021e-19 $X=3.82 $Y=0.38
r17 8 11 71.8268 $w=2.08e-07 $l=1.36e-06 $layer=LI1_cond $X=2.46 $Y=0.36
+ $X2=3.82 $Y2=0.36
r18 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.235 $X2=3.82 $Y2=0.38
r19 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND4B_2%A_655_47# 1 2 3 10 16 18 22 25
c39 25 0 1.59237e-19 $X=4.285 $Y=0.76
r40 20 22 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=5.172 $Y=0.715
+ $X2=5.172 $Y2=0.38
r41 19 25 5.71385 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=4.455 $Y=0.81
+ $X2=4.305 $Y2=0.76
r42 18 20 7.51555 $w=1.9e-07 $l=2.09175e-07 $layer=LI1_cond $X=5.005 $Y=0.81
+ $X2=5.172 $Y2=0.715
r43 18 19 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=5.005 $Y=0.81
+ $X2=4.455 $Y2=0.81
r44 14 25 0.905018 $w=2.6e-07 $l=1.54677e-07 $layer=LI1_cond $X=4.285 $Y=0.615
+ $X2=4.305 $Y2=0.76
r45 14 16 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.285 $Y=0.615
+ $X2=4.285 $Y2=0.42
r46 10 25 5.71385 $w=2.3e-07 $l=1.54919e-07 $layer=LI1_cond $X=4.155 $Y=0.77
+ $X2=4.305 $Y2=0.76
r47 10 12 32.2257 $w=2.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.155 $Y=0.77
+ $X2=3.4 $Y2=0.77
r48 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.035
+ $Y=0.235 $X2=5.17 $Y2=0.38
r49 2 25 182 $w=1.7e-07 $l=6.08379e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.285 $Y2=0.76
r50 2 16 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.285 $Y2=0.42
r51 1 12 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.235 $X2=3.4 $Y2=0.72
.ends


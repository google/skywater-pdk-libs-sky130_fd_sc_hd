* File: sky130_fd_sc_hd__and4_2.spice.SKY130_FD_SC_HD__AND4_2.pxi
* Created: Thu Aug 27 14:08:27 2020
* 
x_PM_SKY130_FD_SC_HD__AND4_2%A N_A_M1010_g N_A_M1005_g A A A A N_A_c_67_n
+ PM_SKY130_FD_SC_HD__AND4_2%A
x_PM_SKY130_FD_SC_HD__AND4_2%B N_B_M1000_g N_B_M1004_g B B N_B_c_98_n
+ PM_SKY130_FD_SC_HD__AND4_2%B
x_PM_SKY130_FD_SC_HD__AND4_2%C N_C_M1009_g N_C_M1001_g C C C N_C_c_134_n C
+ PM_SKY130_FD_SC_HD__AND4_2%C
x_PM_SKY130_FD_SC_HD__AND4_2%D N_D_M1011_g N_D_M1007_g D D D N_D_c_171_n
+ PM_SKY130_FD_SC_HD__AND4_2%D
x_PM_SKY130_FD_SC_HD__AND4_2%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1005_d
+ N_A_27_47#_M1001_d N_A_27_47#_c_207_n N_A_27_47#_M1002_g N_A_27_47#_M1003_g
+ N_A_27_47#_c_208_n N_A_27_47#_M1006_g N_A_27_47#_M1008_g N_A_27_47#_c_209_n
+ N_A_27_47#_c_215_n N_A_27_47#_c_216_n N_A_27_47#_c_217_n N_A_27_47#_c_218_n
+ N_A_27_47#_c_219_n N_A_27_47#_c_230_n N_A_27_47#_c_220_n N_A_27_47#_c_221_n
+ N_A_27_47#_c_210_n N_A_27_47#_c_211_n PM_SKY130_FD_SC_HD__AND4_2%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4_2%VPWR N_VPWR_M1005_s N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_M1008_s N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n
+ VPWR N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_311_n
+ PM_SKY130_FD_SC_HD__AND4_2%VPWR
x_PM_SKY130_FD_SC_HD__AND4_2%X N_X_M1002_d N_X_M1003_d X X X X X X N_X_c_367_n X
+ X PM_SKY130_FD_SC_HD__AND4_2%X
x_PM_SKY130_FD_SC_HD__AND4_2%VGND N_VGND_M1011_d N_VGND_M1006_s N_VGND_c_393_n
+ N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n VGND
+ N_VGND_c_398_n N_VGND_c_399_n PM_SKY130_FD_SC_HD__AND4_2%VGND
cc_1 VNB N_A_M1010_g 0.0333566f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.0123275f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_A_c_67_n 0.0434142f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_M1000_g 0.0290309f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB B 0.00433576f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_6 VNB N_B_c_98_n 0.0223143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_C_M1009_g 0.0295632f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_8 VNB C 0.00314205f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_9 VNB N_C_c_134_n 0.0211728f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_10 VNB C 9.08932e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_M1011_g 0.0322687f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_12 VNB D 0.00302038f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_13 VNB N_D_c_171_n 0.0264732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_207_n 0.0192267f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_15 VNB N_A_27_47#_c_208_n 0.0225075f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_16 VNB N_A_27_47#_c_209_n 0.00423441f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_17 VNB N_A_27_47#_c_210_n 0.00227932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_211_n 0.0583948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_311_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB X 0.00201168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_393_n 0.00689263f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_22 VNB N_VGND_c_394_n 0.0115788f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_23 VNB N_VGND_c_395_n 0.0293542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_396_n 0.0650884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_397_n 0.00452017f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_26 VNB N_VGND_c_398_n 0.0189827f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.53
cc_27 VNB N_VGND_c_399_n 0.200677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_A_M1005_g 0.0543554f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_29 VPB A 0.0352093f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_30 VPB N_A_c_67_n 0.0122403f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_31 VPB N_B_M1004_g 0.0536847f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_32 VPB B 0.00202659f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_33 VPB N_B_c_98_n 0.0045253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_C_M1001_g 0.0514578f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_35 VPB N_C_c_134_n 0.00434406f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_36 VPB C 9.67007e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_D_M1007_g 0.057054f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_38 VPB D 0.00149309f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_39 VPB N_D_c_171_n 0.00617182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_M1003_g 0.0222598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_M1008_g 0.0265747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_209_n 0.00182681f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_43 VPB N_A_27_47#_c_215_n 0.00802897f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.87
cc_44 VPB N_A_27_47#_c_216_n 0.0140507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_217_n 0.00865494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_218_n 0.00479524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_219_n 0.00340454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_220_n 0.00927739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_221_n 0.00581074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_210_n 3.22892e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_211_n 0.0137597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_312_n 0.010303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_313_n 0.0128048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_314_n 0.0170817f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_55 VPB N_VPWR_c_315_n 0.0121186f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_56 VPB N_VPWR_c_316_n 0.0055866f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_57 VPB N_VPWR_c_317_n 0.0118719f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.53
cc_58 VPB N_VPWR_c_318_n 0.0316095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_319_n 0.0241746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_320_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_321_n 0.0183167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_322_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_311_n 0.0434836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB X 0.00240359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 N_A_M1010_g N_B_M1000_g 0.0241025f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_B_M1004_g 0.0264512f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_67 N_A_M1010_g B 8.86104e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_c_67_n N_B_c_98_n 0.0241025f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1010_g N_A_27_47#_c_209_n 0.0132083f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_27_47#_c_209_n 0.003442f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_71 A N_A_27_47#_c_209_n 0.0523589f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_c_67_n N_A_27_47#_c_209_n 0.00822859f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_A_27_47#_c_215_n 0.00410577f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_215_n 0.0229715f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_M1010_g N_A_27_47#_c_230_n 0.0133769f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_76 A N_A_27_47#_c_230_n 0.0129122f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_77 N_A_c_67_n N_A_27_47#_c_230_n 0.0018399f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_A_27_47#_c_220_n 0.00674131f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_79 A N_A_27_47#_c_220_n 0.0137695f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_80 A N_VPWR_M1005_s 0.00232353f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_81 N_A_M1005_g N_VPWR_c_313_n 0.00912703f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_82 A N_VPWR_c_313_n 0.0163288f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A_M1005_g N_VPWR_c_314_n 0.0046653f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_VPWR_c_311_n 0.0081138f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_85 A N_VPWR_c_311_n 0.00103325f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_M1010_g N_VGND_c_396_n 0.00357877f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_87 A N_VGND_c_396_n 7.89669e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_M1010_g N_VGND_c_399_n 0.0062704f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_89 A N_VGND_c_399_n 0.00167133f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_90 N_B_M1000_g N_C_M1009_g 0.0261617f $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_91 B N_C_M1009_g 0.00666548f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_92 N_B_M1004_g N_C_M1001_g 0.0295302f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_93 N_B_M1000_g C 5.04318e-19 $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_94 B C 0.0564166f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_95 N_B_c_98_n N_C_c_134_n 0.0153179f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_96 B C 0.0131522f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_97 N_B_M1000_g N_A_27_47#_c_209_n 0.00480689f $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_98 N_B_M1004_g N_A_27_47#_c_209_n 0.00336799f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_99 B N_A_27_47#_c_209_n 0.0459638f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_100 N_B_M1004_g N_A_27_47#_c_215_n 0.00825436f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_101 N_B_M1004_g N_A_27_47#_c_216_n 0.0158535f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_102 B N_A_27_47#_c_216_n 0.0282582f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_103 N_B_c_98_n N_A_27_47#_c_216_n 0.00216998f $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_M1000_g N_A_27_47#_c_230_n 0.00537407f $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_105 B N_A_27_47#_c_230_n 0.010879f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_106 N_B_c_98_n N_A_27_47#_c_220_n 4.83855e-19 $X=0.975 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VPWR_c_313_n 5.01889e-19 $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VPWR_c_314_n 0.00585385f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_VPWR_c_315_n 0.00378136f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_VPWR_c_311_n 0.0109372f $X=0.975 $Y=2.275 $X2=0 $Y2=0
cc_111 B A_198_47# 0.00558091f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_112 N_B_M1000_g N_VGND_c_396_n 0.00456292f $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_113 B N_VGND_c_396_n 0.0108559f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_114 N_B_M1000_g N_VGND_c_399_n 0.00762877f $X=0.915 $Y=0.445 $X2=0 $Y2=0
cc_115 B N_VGND_c_399_n 0.0118708f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_116 N_C_M1009_g N_D_M1011_g 0.0319714f $X=1.445 $Y=0.445 $X2=0 $Y2=0
cc_117 C N_D_M1011_g 0.00505898f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_118 N_C_M1001_g N_D_M1007_g 0.0381082f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_119 N_C_M1009_g D 5.1265e-19 $X=1.445 $Y=0.445 $X2=0 $Y2=0
cc_120 C D 0.0542882f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_121 N_C_c_134_n D 3.74081e-19 $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_122 C D 0.0120144f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_123 N_C_c_134_n N_D_c_171_n 0.0204248f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_124 C N_D_c_171_n 9.92458e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_125 N_C_M1001_g N_A_27_47#_c_216_n 0.0154498f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_126 N_C_c_134_n N_A_27_47#_c_216_n 0.00217887f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_127 C N_A_27_47#_c_216_n 0.0125872f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_128 N_C_M1001_g N_A_27_47#_c_217_n 0.00813665f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_129 N_C_c_134_n N_A_27_47#_c_221_n 0.00122005f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_130 C N_A_27_47#_c_221_n 0.0114677f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_131 N_C_M1001_g N_VPWR_c_315_n 0.0050897f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_132 N_C_M1001_g N_VPWR_c_319_n 0.00585385f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_133 N_C_M1001_g N_VPWR_c_311_n 0.0107669f $X=1.495 $Y=2.275 $X2=0 $Y2=0
cc_134 C A_304_47# 0.00421027f $X=1.53 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_135 N_C_M1009_g N_VGND_c_396_n 0.00455696f $X=1.445 $Y=0.445 $X2=0 $Y2=0
cc_136 C N_VGND_c_396_n 0.00914931f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_137 N_C_M1009_g N_VGND_c_399_n 0.00770669f $X=1.445 $Y=0.445 $X2=0 $Y2=0
cc_138 C N_VGND_c_399_n 0.00998001f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_139 N_D_M1011_g N_A_27_47#_c_207_n 0.00793557f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_140 D N_A_27_47#_c_207_n 0.00257271f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_141 N_D_M1007_g N_A_27_47#_M1003_g 0.0173658f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_142 N_D_M1007_g N_A_27_47#_c_217_n 0.00740742f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_143 N_D_M1007_g N_A_27_47#_c_218_n 0.0177483f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_144 D N_A_27_47#_c_218_n 0.0201637f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_145 N_D_c_171_n N_A_27_47#_c_218_n 0.0015341f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_146 N_D_M1007_g N_A_27_47#_c_219_n 0.00345909f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_147 D N_A_27_47#_c_219_n 7.54467e-19 $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_148 D N_A_27_47#_c_210_n 0.0188787f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_149 N_D_c_171_n N_A_27_47#_c_210_n 0.00153285f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_150 D N_A_27_47#_c_211_n 8.54683e-19 $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_151 N_D_c_171_n N_A_27_47#_c_211_n 0.0168563f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_152 N_D_M1007_g N_VPWR_c_316_n 0.00942361f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_153 N_D_M1007_g N_VPWR_c_319_n 0.00585385f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_154 N_D_M1007_g N_VPWR_c_311_n 0.0114739f $X=1.925 $Y=2.275 $X2=0 $Y2=0
cc_155 D N_VGND_M1011_d 0.0036301f $X=1.99 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_156 N_D_M1011_g N_VGND_c_393_n 0.00687546f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_157 D N_VGND_c_393_n 0.0368405f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_158 N_D_M1011_g N_VGND_c_396_n 0.00455696f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_159 D N_VGND_c_396_n 0.00777742f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_160 N_D_M1011_g N_VGND_c_399_n 0.00810877f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_161 D N_VGND_c_399_n 0.00857482f $X=1.99 $Y=0.425 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_218_n N_VPWR_M1007_d 0.0202922f $X=2.33 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_219_n N_VPWR_M1007_d 2.254e-19 $X=2.442 $Y=1.495 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_215_n N_VPWR_c_314_n 0.0171956f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_215_n N_VPWR_c_315_n 0.0101331f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_216_n N_VPWR_c_315_n 0.0211463f $X=1.585 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_217_n N_VPWR_c_315_n 0.0114393f $X=1.71 $Y=2.3 $X2=0 $Y2=0
cc_168 N_A_27_47#_M1003_g N_VPWR_c_316_n 0.00860349f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_217_n N_VPWR_c_316_n 0.0184784f $X=1.71 $Y=2.3 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_218_n N_VPWR_c_316_n 0.0268644f $X=2.33 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_210_n N_VPWR_c_316_n 2.20379e-19 $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_211_n N_VPWR_c_316_n 6.55132e-19 $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1008_g N_VPWR_c_318_n 0.00495855f $X=3.17 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_217_n N_VPWR_c_319_n 0.0145827f $X=1.71 $Y=2.3 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1003_g N_VPWR_c_321_n 0.00541359f $X=2.69 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1008_g N_VPWR_c_321_n 0.00583607f $X=3.17 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1005_d N_VPWR_c_311_n 0.0064797f $X=0.545 $Y=2.065 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1001_d N_VPWR_c_311_n 0.00327378f $X=1.57 $Y=2.065 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1003_g N_VPWR_c_311_n 0.0104145f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1008_g N_VPWR_c_311_n 0.0115395f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_215_n N_VPWR_c_311_n 0.00954569f $X=0.725 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_217_n N_VPWR_c_311_n 0.00955092f $X=1.71 $Y=2.3 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1003_g X 0.0146211f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_207_n N_X_c_367_n 0.00738638f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_211_n N_X_c_367_n 0.00166806f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_207_n X 0.00252118f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_47#_M1003_g X 0.00103112f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_208_n X 0.00279269f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_27_47#_M1008_g X 0.00438042f $X=3.17 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_219_n X 0.00610696f $X=2.442 $Y=1.495 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_210_n X 0.0173706f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_211_n X 0.0302953f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1003_g X 0.00332862f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_218_n X 0.0134082f $X=2.33 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_211_n X 0.00177765f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_209_n A_109_47# 8.40128e-19 $X=0.585 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_197 N_A_27_47#_c_230_n A_109_47# 0.00457961f $X=0.585 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_198 N_A_27_47#_c_207_n N_VGND_c_393_n 0.00329057f $X=2.69 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_210_n N_VGND_c_393_n 0.0184228f $X=2.56 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_211_n N_VGND_c_393_n 0.00354291f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_208_n N_VGND_c_395_n 0.00491123f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_230_n N_VGND_c_396_n 0.0289623f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_207_n N_VGND_c_398_n 0.00541489f $X=2.69 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_27_47#_c_208_n N_VGND_c_398_n 0.00585385f $X=3.17 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_M1010_s N_VGND_c_399_n 0.00230958f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_207_n N_VGND_c_399_n 0.0102793f $X=2.69 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_208_n N_VGND_c_399_n 0.0115781f $X=3.17 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_230_n N_VGND_c_399_n 0.0179555f $X=0.585 $Y=0.42 $X2=0 $Y2=0
cc_209 N_VPWR_c_311_n N_X_M1003_d 0.0035017f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_321_n X 0.0202561f $X=3.245 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_311_n X 0.0126193f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_212 X N_VGND_c_393_n 8.90272e-19 $X=2.985 $Y=0.85 $X2=0 $Y2=0
cc_213 N_X_c_367_n N_VGND_c_398_n 0.0159697f $X=2.982 $Y=0.805 $X2=0 $Y2=0
cc_214 N_X_M1002_d N_VGND_c_399_n 0.00349438f $X=2.765 $Y=0.235 $X2=0 $Y2=0
cc_215 N_X_c_367_n N_VGND_c_399_n 0.0123804f $X=2.982 $Y=0.805 $X2=0 $Y2=0
cc_216 A_109_47# N_VGND_c_399_n 0.00826258f $X=0.545 $Y=0.235 $X2=1.71 $Y2=2.3
cc_217 A_198_47# N_VGND_c_399_n 0.00766156f $X=0.99 $Y=0.235 $X2=0 $Y2=0
cc_218 A_304_47# N_VGND_c_399_n 0.00737302f $X=1.52 $Y=0.235 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__xor2_2.pxi.spice
* Created: Tue Sep  1 19:33:28 2020
* 
x_PM_SKY130_FD_SC_HD__XOR2_2%A N_A_c_103_n N_A_M1011_g N_A_M1004_g N_A_c_104_n
+ N_A_M1016_g N_A_M1019_g N_A_c_105_n N_A_M1005_g N_A_M1000_g N_A_c_106_n
+ N_A_M1012_g N_A_M1002_g N_A_c_116_n N_A_c_107_n N_A_c_108_n N_A_c_109_n
+ N_A_c_139_p N_A_c_118_n N_A_c_119_n A N_A_c_110_n N_A_c_111_n
+ PM_SKY130_FD_SC_HD__XOR2_2%A
x_PM_SKY130_FD_SC_HD__XOR2_2%B N_B_c_234_n N_B_M1009_g N_B_M1013_g N_B_c_235_n
+ N_B_M1015_g N_B_M1014_g N_B_c_236_n N_B_M1001_g N_B_M1003_g N_B_c_237_n
+ N_B_M1018_g N_B_M1006_g B N_B_c_239_n N_B_c_240_n N_B_c_271_n N_B_c_241_n
+ N_B_c_242_n N_B_c_243_n PM_SKY130_FD_SC_HD__XOR2_2%B
x_PM_SKY130_FD_SC_HD__XOR2_2%A_112_47# N_A_112_47#_M1011_s N_A_112_47#_M1009_d
+ N_A_112_47#_M1013_s N_A_112_47#_c_354_n N_A_112_47#_M1007_g
+ N_A_112_47#_M1010_g N_A_112_47#_c_355_n N_A_112_47#_M1008_g
+ N_A_112_47#_M1017_g N_A_112_47#_c_356_n N_A_112_47#_c_357_n
+ N_A_112_47#_c_358_n N_A_112_47#_c_381_n N_A_112_47#_c_368_n
+ N_A_112_47#_c_387_n N_A_112_47#_c_359_n N_A_112_47#_c_392_n
+ N_A_112_47#_c_369_n N_A_112_47#_c_370_n N_A_112_47#_c_371_n
+ N_A_112_47#_c_372_n N_A_112_47#_c_360_n N_A_112_47#_c_361_n
+ N_A_112_47#_c_362_n N_A_112_47#_c_363_n N_A_112_47#_c_406_n
+ N_A_112_47#_c_364_n PM_SKY130_FD_SC_HD__XOR2_2%A_112_47#
x_PM_SKY130_FD_SC_HD__XOR2_2%A_27_297# N_A_27_297#_M1004_s N_A_27_297#_M1019_s
+ N_A_27_297#_M1014_d N_A_27_297#_c_531_n N_A_27_297#_c_546_n
+ N_A_27_297#_c_527_n N_A_27_297#_c_523_n N_A_27_297#_c_524_n
+ N_A_27_297#_c_530_n N_A_27_297#_c_554_n PM_SKY130_FD_SC_HD__XOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HD__XOR2_2%VPWR N_VPWR_M1004_d N_VPWR_M1000_s N_VPWR_M1003_s
+ N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n
+ VPWR N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_579_n
+ N_VPWR_c_589_n N_VPWR_c_590_n PM_SKY130_FD_SC_HD__XOR2_2%VPWR
x_PM_SKY130_FD_SC_HD__XOR2_2%A_470_297# N_A_470_297#_M1000_d
+ N_A_470_297#_M1002_d N_A_470_297#_M1006_d N_A_470_297#_M1010_d
+ N_A_470_297#_M1017_d N_A_470_297#_c_672_n N_A_470_297#_c_670_n
+ N_A_470_297#_c_673_n N_A_470_297#_c_699_n N_A_470_297#_c_683_n
+ N_A_470_297#_c_713_p N_A_470_297#_c_668_n N_A_470_297#_c_686_n
+ N_A_470_297#_c_674_n N_A_470_297#_c_669_n
+ PM_SKY130_FD_SC_HD__XOR2_2%A_470_297#
x_PM_SKY130_FD_SC_HD__XOR2_2%X N_X_M1001_d N_X_M1007_d N_X_M1010_s N_X_c_715_n
+ N_X_c_716_n N_X_c_717_n N_X_c_718_n X N_X_c_748_n PM_SKY130_FD_SC_HD__XOR2_2%X
x_PM_SKY130_FD_SC_HD__XOR2_2%VGND N_VGND_M1011_d N_VGND_M1016_d N_VGND_M1015_s
+ N_VGND_M1005_d N_VGND_M1007_s N_VGND_M1008_s N_VGND_c_766_n N_VGND_c_767_n
+ N_VGND_c_768_n N_VGND_c_769_n N_VGND_c_770_n N_VGND_c_771_n N_VGND_c_772_n
+ N_VGND_c_773_n N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n N_VGND_c_777_n
+ N_VGND_c_778_n N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ VGND N_VGND_c_783_n N_VGND_c_784_n PM_SKY130_FD_SC_HD__XOR2_2%VGND
x_PM_SKY130_FD_SC_HD__XOR2_2%A_470_47# N_A_470_47#_M1005_s N_A_470_47#_M1012_s
+ N_A_470_47#_M1018_s N_A_470_47#_c_865_n N_A_470_47#_c_866_n
+ N_A_470_47#_c_867_n N_A_470_47#_c_878_n N_A_470_47#_c_880_n
+ N_A_470_47#_c_868_n PM_SKY130_FD_SC_HD__XOR2_2%A_470_47#
cc_1 VNB N_A_c_103_n 0.0191865f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_c_104_n 0.0160105f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_3 VNB N_A_c_105_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=0.995
cc_4 VNB N_A_c_106_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=0.995
cc_5 VNB N_A_c_107_n 9.96253e-19 $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=1.445
cc_6 VNB N_A_c_108_n 0.00215578f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.175
cc_7 VNB N_A_c_109_n 0.0263018f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=1.16
cc_8 VNB N_A_c_110_n 0.0344148f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_9 VNB N_A_c_111_n 0.0392959f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.16
cc_10 VNB N_B_c_234_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_11 VNB N_B_c_235_n 0.0215f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.995
cc_12 VNB N_B_c_236_n 0.0167643f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=0.995
cc_13 VNB N_B_c_237_n 0.022021f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=0.995
cc_14 VNB B 0.00495909f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.275
cc_15 VNB N_B_c_239_n 0.00325917f $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=1.275
cc_16 VNB N_B_c_240_n 0.00336897f $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=1.445
cc_17 VNB N_B_c_241_n 0.00203829f $X=-0.19 $Y=-0.24 $X2=1.71 $Y2=1.53
cc_18 VNB N_B_c_242_n 0.0366805f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.445
cc_19 VNB N_B_c_243_n 0.0395261f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=1.16
cc_20 VNB N_A_112_47#_c_354_n 0.0214858f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_21 VNB N_A_112_47#_c_355_n 0.0191719f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=0.56
cc_22 VNB N_A_112_47#_c_356_n 0.0189501f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.325
cc_23 VNB N_A_112_47#_c_357_n 0.00411695f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.985
cc_24 VNB N_A_112_47#_c_358_n 0.0077223f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.985
cc_25 VNB N_A_112_47#_c_359_n 0.00462689f $X=-0.19 $Y=-0.24 $X2=3.065 $Y2=1.175
cc_26 VNB N_A_112_47#_c_360_n 0.00117487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_112_47#_c_361_n 0.0037828f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_28 VNB N_A_112_47#_c_362_n 0.00210839f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_29 VNB N_A_112_47#_c_363_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=1.16
cc_30 VNB N_A_112_47#_c_364_n 0.0390403f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_579_n 0.250759f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.445
cc_32 VNB N_X_c_715_n 0.0158993f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.56
cc_33 VNB N_X_c_716_n 0.0234946f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=0.995
cc_34 VNB N_X_c_717_n 0.00203744f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=1.985
cc_35 VNB N_X_c_718_n 0.0145224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_766_n 0.0112403f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=1.985
cc_37 VNB N_VGND_c_767_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_768_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.325
cc_39 VNB N_VGND_c_769_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.275
cc_40 VNB N_VGND_c_770_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.175
cc_41 VNB N_VGND_c_771_n 0.00420911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_772_n 0.00420911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_773_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.53
cc_44 VNB N_VGND_c_774_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=1.71 $Y2=1.53
cc_45 VNB N_VGND_c_775_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_776_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=1.16
cc_47 VNB N_VGND_c_777_n 0.0205874f $X=-0.19 $Y=-0.24 $X2=0.71 $Y2=1.16
cc_48 VNB N_VGND_c_778_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.16
cc_49 VNB N_VGND_c_779_n 0.0393681f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=1.16
cc_50 VNB N_VGND_c_780_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_781_n 0.0185607f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=1.16
cc_52 VNB N_VGND_c_782_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_783_n 0.0115962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_784_n 0.3108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_470_47#_c_865_n 0.00547724f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=1.985
cc_56 VNB N_A_470_47#_c_866_n 0.00429401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_470_47#_c_867_n 0.0047325f $X=-0.19 $Y=-0.24 $X2=2.685 $Y2=0.995
cc_58 VNB N_A_470_47#_c_868_n 0.00300719f $X=-0.19 $Y=-0.24 $X2=3.105 $Y2=0.995
cc_59 VPB N_A_M1004_g 0.0219153f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_60 VPB N_A_M1019_g 0.0178886f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_61 VPB N_A_M1000_g 0.025044f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=1.985
cc_62 VPB N_A_M1002_g 0.0184042f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=1.985
cc_63 VPB N_A_c_116_n 9.67218e-19 $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.445
cc_64 VPB N_A_c_107_n 0.00477515f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.445
cc_65 VPB N_A_c_118_n 3.34033e-19 $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.53
cc_66 VPB N_A_c_119_n 0.0048839f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.53
cc_67 VPB N_A_c_110_n 0.00472787f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.16
cc_68 VPB N_A_c_111_n 0.00581932f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=1.16
cc_69 VPB N_B_M1013_g 0.0183437f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.985
cc_70 VPB N_B_M1014_g 0.0228017f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_71 VPB N_B_M1003_g 0.0190422f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=1.985
cc_72 VPB N_B_M1006_g 0.0234854f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=1.985
cc_73 VPB N_B_c_240_n 0.00164129f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.445
cc_74 VPB N_B_c_242_n 0.00453888f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.445
cc_75 VPB N_B_c_243_n 0.00578959f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=1.16
cc_76 VPB N_A_112_47#_M1010_g 0.0218603f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=0.995
cc_77 VPB N_A_112_47#_M1017_g 0.0220154f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=0.995
cc_78 VPB N_A_112_47#_c_356_n 0.019177f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=1.325
cc_79 VPB N_A_112_47#_c_368_n 0.00712491f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.275
cc_80 VPB N_A_112_47#_c_369_n 0.00462339f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.16
cc_81 VPB N_A_112_47#_c_370_n 0.00281079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_112_47#_c_371_n 0.0262927f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.53
cc_83 VPB N_A_112_47#_c_372_n 0.00246874f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.53
cc_84 VPB N_A_112_47#_c_360_n 0.00347332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_112_47#_c_364_n 0.00428376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_27_297#_c_523_n 0.0106541f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=1.325
cc_87 VPB N_A_27_297#_c_524_n 0.0078945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_580_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.985
cc_89 VPB N_VPWR_c_581_n 0.00454762f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=0.56
cc_90 VPB N_VPWR_c_582_n 0.00485375f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=1.985
cc_91 VPB N_VPWR_c_583_n 0.0485326f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=0.56
cc_92 VPB N_VPWR_c_584_n 0.00478242f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=0.56
cc_93 VPB N_VPWR_c_585_n 0.0176443f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=1.985
cc_94 VPB N_VPWR_c_586_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.16
cc_95 VPB N_VPWR_c_587_n 0.0524598f $X=-0.19 $Y=1.305 $X2=1.71 $Y2=1.53
cc_96 VPB N_VPWR_c_579_n 0.058756f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.445
cc_97 VPB N_VPWR_c_589_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_590_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_470_297#_c_668_n 0.00483491f $X=-0.19 $Y=1.305 $X2=3.065 $Y2=1.16
cc_100 VPB N_A_470_297#_c_669_n 0.0112805f $X=-0.19 $Y=1.305 $X2=0.875 $Y2=1.53
cc_101 VPB N_X_c_716_n 0.00762153f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=0.995
cc_102 VPB X 0.0209804f $X=-0.19 $Y=1.305 $X2=3.105 $Y2=0.56
cc_103 N_A_c_104_n N_B_c_234_n 0.0258694f $X=0.905 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_104 N_A_M1019_g N_B_M1013_g 0.044538f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_c_116_n N_B_M1013_g 6.08253e-19 $X=0.79 $Y=1.445 $X2=0 $Y2=0
cc_106 N_A_c_107_n N_B_M1013_g 6.92959e-19 $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_107 N_A_c_119_n N_B_M1013_g 0.010197f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A_c_107_n N_B_M1014_g 0.00457937f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_109 N_A_c_119_n N_B_M1014_g 0.00986014f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_110 N_A_c_106_n N_B_c_236_n 0.0238362f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_M1002_g N_B_M1003_g 0.028954f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_c_109_n B 0.0141425f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_c_111_n B 5.8921e-19 $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_108_n N_B_c_239_n 0.0140423f $X=1.88 $Y=1.175 $X2=0 $Y2=0
cc_115 N_A_c_109_n N_B_c_239_n 0.0628729f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_119_n N_B_c_239_n 0.00627342f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_117 N_A_c_116_n N_B_c_240_n 0.00141189f $X=0.79 $Y=1.445 $X2=0 $Y2=0
cc_118 N_A_c_107_n N_B_c_240_n 9.2125e-19 $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_119 N_A_c_108_n N_B_c_240_n 2.63318e-19 $X=1.88 $Y=1.175 $X2=0 $Y2=0
cc_120 N_A_c_139_p N_B_c_240_n 0.0065861f $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_121 N_A_c_119_n N_B_c_240_n 0.00822356f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_122 N_A_c_110_n N_B_c_240_n 0.00479793f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_c_109_n N_B_c_271_n 2.48533e-19 $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_108_n N_B_c_241_n 0.0138658f $X=1.88 $Y=1.175 $X2=0 $Y2=0
cc_125 N_A_c_139_p N_B_c_241_n 0.0133176f $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_126 N_A_c_119_n N_B_c_241_n 0.0318166f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_127 N_A_c_110_n N_B_c_241_n 0.00155395f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_116_n N_B_c_242_n 2.62013e-19 $X=0.79 $Y=1.445 $X2=0 $Y2=0
cc_129 N_A_c_107_n N_B_c_242_n 0.0026345f $X=1.795 $Y=1.445 $X2=0 $Y2=0
cc_130 N_A_c_108_n N_B_c_242_n 0.0144999f $X=1.88 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A_c_119_n N_B_c_242_n 0.00254515f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_132 N_A_c_110_n N_B_c_242_n 0.0180897f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_c_109_n N_B_c_243_n 5.94456e-19 $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_111_n N_B_c_243_n 0.0195749f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_119_n N_A_112_47#_M1013_s 0.00165831f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_136 N_A_c_103_n N_A_112_47#_c_356_n 0.0264874f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_116_n N_A_112_47#_c_356_n 0.00666755f $X=0.79 $Y=1.445 $X2=0 $Y2=0
cc_138 N_A_c_139_p N_A_112_47#_c_356_n 0.0110237f $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_139 N_A_c_118_n N_A_112_47#_c_356_n 0.0072664f $X=0.875 $Y=1.53 $X2=0 $Y2=0
cc_140 N_A_c_103_n N_A_112_47#_c_357_n 0.0138637f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_M1004_g N_A_112_47#_c_381_n 0.0163198f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1019_g N_A_112_47#_c_381_n 0.010512f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_c_139_p N_A_112_47#_c_381_n 0.00391811f $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_144 N_A_c_118_n N_A_112_47#_c_381_n 0.00815634f $X=0.875 $Y=1.53 $X2=0 $Y2=0
cc_145 N_A_c_119_n N_A_112_47#_c_381_n 0.0269978f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A_c_110_n N_A_112_47#_c_381_n 0.00115169f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_103_n N_A_112_47#_c_387_n 0.0109314f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_104_n N_A_112_47#_c_387_n 0.00630972f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_104_n N_A_112_47#_c_359_n 0.00991999f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_139_p N_A_112_47#_c_359_n 9.99879e-19 $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_151 N_A_c_119_n N_A_112_47#_c_359_n 0.00659421f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_152 N_A_c_104_n N_A_112_47#_c_392_n 5.22228e-19 $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_109_n N_A_112_47#_c_369_n 0.00468456f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_c_119_n N_A_112_47#_c_369_n 0.0107313f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_155 N_A_M1000_g N_A_112_47#_c_370_n 0.0043148f $X=2.685 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1000_g N_A_112_47#_c_371_n 0.0122132f $X=2.685 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_A_112_47#_c_371_n 0.0102491f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_c_109_n N_A_112_47#_c_371_n 0.0667248f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_c_111_n N_A_112_47#_c_371_n 0.00309155f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_109_n N_A_112_47#_c_372_n 0.0127997f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_c_119_n N_A_112_47#_c_372_n 0.0154683f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_162 N_A_c_103_n N_A_112_47#_c_363_n 0.00165338f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_104_n N_A_112_47#_c_363_n 0.00112787f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_139_p N_A_112_47#_c_363_n 0.025389f $X=0.79 $Y=1.175 $X2=0 $Y2=0
cc_165 N_A_c_110_n N_A_112_47#_c_363_n 0.00230339f $X=0.905 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_c_119_n N_A_112_47#_c_406_n 0.0116047f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_c_119_n N_A_27_297#_M1019_s 0.00162081f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_168 N_A_c_119_n N_A_27_297#_M1014_d 0.00143861f $X=1.71 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_M1004_g N_A_27_297#_c_527_n 0.00237973f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_M1019_g N_A_27_297#_c_527_n 0.00237973f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_M1004_g N_A_27_297#_c_523_n 6.70354e-19 $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_M1019_g N_A_27_297#_c_530_n 5.83285e-19 $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_c_118_n N_VPWR_M1004_d 0.00234844f $X=0.875 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_M1004_g N_VPWR_c_580_n 0.00321647f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_M1019_g N_VPWR_c_580_n 0.00321647f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_M1000_g N_VPWR_c_581_n 0.00302074f $X=2.685 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_M1002_g N_VPWR_c_581_n 0.00157837f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A_M1019_g N_VPWR_c_583_n 0.00585385f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_M1000_g N_VPWR_c_583_n 0.00585385f $X=2.685 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_M1004_g N_VPWR_c_585_n 0.00585385f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_M1002_g N_VPWR_c_586_n 0.00585385f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_M1004_g N_VPWR_c_579_n 0.00577127f $X=0.485 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1019_g N_VPWR_c_579_n 0.00483015f $X=0.905 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1000_g N_VPWR_c_579_n 0.0072109f $X=2.685 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_M1002_g N_VPWR_c_579_n 0.00591203f $X=3.105 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_M1000_g N_A_470_297#_c_670_n 0.00959653f $X=2.685 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_M1002_g N_A_470_297#_c_670_n 0.00955237f $X=3.105 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_c_103_n N_VGND_c_767_n 0.00316354f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_104_n N_VGND_c_768_n 0.00146448f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_105_n N_VGND_c_769_n 0.00194637f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_108_n N_VGND_c_769_n 2.22494e-19 $X=1.88 $Y=1.175 $X2=0 $Y2=0
cc_192 N_A_c_109_n N_VGND_c_769_n 0.00470501f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_105_n N_VGND_c_770_n 0.00268723f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_106_n N_VGND_c_770_n 0.00268723f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_103_n N_VGND_c_773_n 0.00423334f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_104_n N_VGND_c_773_n 0.00423334f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_105_n N_VGND_c_777_n 0.00423334f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_c_106_n N_VGND_c_779_n 0.00421816f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_c_103_n N_VGND_c_784_n 0.00668462f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_104_n N_VGND_c_784_n 0.0057435f $X=0.905 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_105_n N_VGND_c_784_n 0.00704237f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_106_n N_VGND_c_784_n 0.00579251f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_105_n N_A_470_47#_c_865_n 0.00630972f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_106_n N_A_470_47#_c_865_n 5.22228e-19 $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_c_105_n N_A_470_47#_c_866_n 0.00860496f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A_c_106_n N_A_470_47#_c_866_n 0.011056f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_c_109_n N_A_470_47#_c_866_n 0.0388239f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_c_111_n N_A_470_47#_c_866_n 0.0027332f $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_105_n N_A_470_47#_c_867_n 0.00128204f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_109_n N_A_470_47#_c_867_n 0.0251706f $X=3.065 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_c_111_n N_A_470_47#_c_867_n 5.11864e-19 $X=3.105 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_c_105_n N_A_470_47#_c_878_n 4.58193e-19 $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_106_n N_A_470_47#_c_878_n 0.00376498f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_106_n N_A_470_47#_c_880_n 0.00358777f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_M1013_g N_A_112_47#_c_381_n 0.00917601f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B_c_234_n N_A_112_47#_c_387_n 5.22228e-19 $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_234_n N_A_112_47#_c_359_n 0.00972036f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_235_n N_A_112_47#_c_359_n 0.00482542f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B_c_239_n N_A_112_47#_c_359_n 0.00610524f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_220 N_B_c_240_n N_A_112_47#_c_359_n 0.00795571f $X=1.295 $Y=1.19 $X2=0 $Y2=0
cc_221 N_B_c_241_n N_A_112_47#_c_359_n 0.0333186f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_c_242_n N_A_112_47#_c_359_n 0.00279167f $X=1.745 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_c_234_n N_A_112_47#_c_392_n 0.00630972f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_235_n N_A_112_47#_c_392_n 0.00717381f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B_M1014_g N_A_112_47#_c_369_n 0.0109232f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_226 N_B_c_239_n N_A_112_47#_c_369_n 0.00169022f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_227 N_B_M1014_g N_A_112_47#_c_370_n 0.00542416f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_228 N_B_M1003_g N_A_112_47#_c_371_n 0.0105728f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B_M1006_g N_A_112_47#_c_371_n 0.0126757f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_230 B N_A_112_47#_c_371_n 0.0425285f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_231 N_B_c_239_n N_A_112_47#_c_371_n 0.0158942f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_232 N_B_c_271_n N_A_112_47#_c_371_n 0.00706515f $X=3.91 $Y=1.19 $X2=0 $Y2=0
cc_233 N_B_c_243_n N_A_112_47#_c_371_n 0.00344827f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B_M1014_g N_A_112_47#_c_372_n 0.00116202f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B_c_239_n N_A_112_47#_c_372_n 0.00139134f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_236 B N_A_112_47#_c_360_n 9.10568e-19 $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_237 N_B_c_271_n N_A_112_47#_c_360_n 0.00110457f $X=3.91 $Y=1.19 $X2=0 $Y2=0
cc_238 N_B_c_243_n N_A_112_47#_c_360_n 0.00432723f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_239 B N_A_112_47#_c_361_n 0.00578167f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_240 N_B_c_271_n N_A_112_47#_c_361_n 0.00123012f $X=3.91 $Y=1.19 $X2=0 $Y2=0
cc_241 N_B_c_243_n N_A_112_47#_c_361_n 0.00106738f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B_M1013_g N_A_27_297#_c_531_n 0.00825038f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_243 N_B_M1014_g N_A_27_297#_c_531_n 0.00851673f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_244 N_B_M1013_g N_A_27_297#_c_530_n 0.00298436f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_245 N_B_M1014_g N_A_27_297#_c_530_n 7.71958e-19 $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_246 N_B_M1003_g N_VPWR_c_582_n 0.00169496f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_247 N_B_M1006_g N_VPWR_c_582_n 0.00317329f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_248 N_B_M1013_g N_VPWR_c_583_n 0.00357877f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B_M1014_g N_VPWR_c_583_n 0.00357877f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_250 N_B_M1003_g N_VPWR_c_586_n 0.00585385f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_251 N_B_M1006_g N_VPWR_c_587_n 0.00585385f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_252 N_B_M1013_g N_VPWR_c_579_n 0.00508422f $X=1.325 $Y=1.985 $X2=0 $Y2=0
cc_253 N_B_M1014_g N_VPWR_c_579_n 0.00655123f $X=1.745 $Y=1.985 $X2=0 $Y2=0
cc_254 N_B_M1003_g N_VPWR_c_579_n 0.00605104f $X=3.525 $Y=1.985 $X2=0 $Y2=0
cc_255 N_B_M1006_g N_VPWR_c_579_n 0.00734991f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_256 N_B_M1014_g N_A_470_297#_c_672_n 0.00368782f $X=1.745 $Y=1.985 $X2=0
+ $Y2=0
cc_257 N_B_M1014_g N_A_470_297#_c_673_n 5.93156e-19 $X=1.745 $Y=1.985 $X2=0
+ $Y2=0
cc_258 N_B_M1003_g N_A_470_297#_c_674_n 0.00992019f $X=3.525 $Y=1.985 $X2=0
+ $Y2=0
cc_259 N_B_M1006_g N_A_470_297#_c_674_n 0.00991827f $X=4 $Y=1.985 $X2=0 $Y2=0
cc_260 N_B_c_237_n N_X_c_715_n 0.00985078f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_261 N_B_c_237_n N_X_c_717_n 0.00496301f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_262 B N_X_c_717_n 0.0303013f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_263 N_B_c_239_n N_X_c_717_n 9.93721e-19 $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_264 N_B_c_271_n N_X_c_717_n 0.00684958f $X=3.91 $Y=1.19 $X2=0 $Y2=0
cc_265 N_B_c_243_n N_X_c_717_n 0.00361233f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B_c_234_n N_VGND_c_768_n 0.00146448f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_c_235_n N_VGND_c_769_n 0.00316354f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B_c_239_n N_VGND_c_769_n 0.00123192f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_269 N_B_c_237_n N_VGND_c_771_n 0.0019578f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_234_n N_VGND_c_775_n 0.00423334f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B_c_235_n N_VGND_c_775_n 0.00541359f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B_c_236_n N_VGND_c_779_n 0.00357877f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_273 N_B_c_237_n N_VGND_c_779_n 0.00357877f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B_c_234_n N_VGND_c_784_n 0.0057435f $X=1.325 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B_c_235_n N_VGND_c_784_n 0.0108276f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_276 N_B_c_236_n N_VGND_c_784_n 0.00543665f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B_c_237_n N_VGND_c_784_n 0.00669559f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B_c_235_n N_A_470_47#_c_865_n 0.0030909f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B_c_236_n N_A_470_47#_c_866_n 8.19387e-19 $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B_c_239_n N_A_470_47#_c_866_n 0.00928666f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_281 N_B_c_235_n N_A_470_47#_c_867_n 0.00312932f $X=1.745 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_239_n N_A_470_47#_c_867_n 0.00252741f $X=3.765 $Y=1.19 $X2=0 $Y2=0
cc_283 N_B_c_236_n N_A_470_47#_c_868_n 0.0124238f $X=3.525 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_237_n N_A_470_47#_c_868_n 0.00971555f $X=4 $Y=0.995 $X2=0 $Y2=0
cc_285 B N_A_470_47#_c_868_n 0.00447603f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_286 N_A_112_47#_c_356_n N_A_27_297#_M1004_s 0.00542017f $X=0.205 $Y=1.785
+ $X2=-0.19 $Y2=-0.24
cc_287 N_A_112_47#_c_381_n N_A_27_297#_M1004_s 0.00296717f $X=1.41 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_288 N_A_112_47#_c_368_n N_A_27_297#_M1004_s 0.00243062f $X=0.29 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_289 N_A_112_47#_c_381_n N_A_27_297#_M1019_s 0.00311999f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_290 N_A_112_47#_c_369_n N_A_27_297#_M1014_d 0.00580203f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_291 N_A_112_47#_c_370_n N_A_27_297#_M1014_d 0.00230597f $X=2.135 $Y=1.785
+ $X2=0 $Y2=0
cc_292 N_A_112_47#_c_372_n N_A_27_297#_M1014_d 0.0013619f $X=2.22 $Y=1.53 $X2=0
+ $Y2=0
cc_293 N_A_112_47#_M1013_s N_A_27_297#_c_531_n 0.00312348f $X=1.4 $Y=1.485 $X2=0
+ $Y2=0
cc_294 N_A_112_47#_c_381_n N_A_27_297#_c_531_n 0.00477489f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_295 N_A_112_47#_c_369_n N_A_27_297#_c_531_n 0.00506389f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_296 N_A_112_47#_c_406_n N_A_27_297#_c_531_n 0.0112811f $X=1.535 $Y=1.87 $X2=0
+ $Y2=0
cc_297 N_A_112_47#_c_369_n N_A_27_297#_c_546_n 0.0144865f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_298 N_A_112_47#_c_381_n N_A_27_297#_c_527_n 0.014974f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_299 N_A_112_47#_c_381_n N_A_27_297#_c_523_n 0.00242129f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_300 N_A_112_47#_c_368_n N_A_27_297#_c_523_n 0.00499157f $X=0.29 $Y=1.87 $X2=0
+ $Y2=0
cc_301 N_A_112_47#_c_381_n N_A_27_297#_c_524_n 0.0042519f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_302 N_A_112_47#_c_368_n N_A_27_297#_c_524_n 0.0120194f $X=0.29 $Y=1.87 $X2=0
+ $Y2=0
cc_303 N_A_112_47#_c_381_n N_A_27_297#_c_530_n 0.00818191f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_304 N_A_112_47#_c_406_n N_A_27_297#_c_530_n 0.00148888f $X=1.535 $Y=1.87
+ $X2=0 $Y2=0
cc_305 N_A_112_47#_c_381_n N_A_27_297#_c_554_n 0.0112383f $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_306 N_A_112_47#_c_381_n N_VPWR_M1004_d 0.00364797f $X=1.41 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_307 N_A_112_47#_c_371_n N_VPWR_M1000_s 0.00166235f $X=4.615 $Y=1.53 $X2=0
+ $Y2=0
cc_308 N_A_112_47#_c_371_n N_VPWR_M1003_s 0.00224844f $X=4.615 $Y=1.53 $X2=0
+ $Y2=0
cc_309 N_A_112_47#_c_381_n N_VPWR_c_580_n 0.011057f $X=1.41 $Y=1.87 $X2=0 $Y2=0
cc_310 N_A_112_47#_M1010_g N_VPWR_c_587_n 0.00357877f $X=4.94 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_112_47#_M1017_g N_VPWR_c_587_n 0.00357877f $X=5.36 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_112_47#_M1013_s N_VPWR_c_579_n 0.00215227f $X=1.4 $Y=1.485 $X2=0
+ $Y2=0
cc_313 N_A_112_47#_M1010_g N_VPWR_c_579_n 0.00655123f $X=4.94 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_112_47#_M1017_g N_VPWR_c_579_n 0.00629538f $X=5.36 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_112_47#_c_381_n N_VPWR_c_579_n 5.77144e-19 $X=1.41 $Y=1.87 $X2=0
+ $Y2=0
cc_316 N_A_112_47#_c_369_n N_VPWR_c_579_n 0.00660225f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_112_47#_c_371_n N_A_470_297#_M1000_d 0.00303335f $X=4.615 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_318 N_A_112_47#_c_371_n N_A_470_297#_M1002_d 0.00165831f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_319 N_A_112_47#_c_371_n N_A_470_297#_M1006_d 0.0027344f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_320 N_A_112_47#_c_371_n N_A_470_297#_M1010_d 0.0045218f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_321 N_A_112_47#_c_371_n N_A_470_297#_c_670_n 0.0305785f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_322 N_A_112_47#_c_369_n N_A_470_297#_c_673_n 0.0154012f $X=2.05 $Y=1.87 $X2=0
+ $Y2=0
cc_323 N_A_112_47#_c_371_n N_A_470_297#_c_673_n 0.0127945f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_324 N_A_112_47#_M1010_g N_A_470_297#_c_683_n 0.0121306f $X=4.94 $Y=1.985
+ $X2=0 $Y2=0
cc_325 N_A_112_47#_M1017_g N_A_470_297#_c_683_n 0.00988743f $X=5.36 $Y=1.985
+ $X2=0 $Y2=0
cc_326 N_A_112_47#_c_371_n N_A_470_297#_c_668_n 0.0037422f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_327 N_A_112_47#_c_371_n N_A_470_297#_c_686_n 0.0122451f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_328 N_A_112_47#_c_371_n N_A_470_297#_c_674_n 0.0743095f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_329 N_A_112_47#_c_371_n N_A_470_297#_c_669_n 0.0150001f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_330 N_A_112_47#_c_362_n N_A_470_297#_c_669_n 0.00160143f $X=5.11 $Y=1.16
+ $X2=0 $Y2=0
cc_331 N_A_112_47#_c_354_n N_X_c_715_n 0.0109318f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_112_47#_c_371_n N_X_c_715_n 0.0178076f $X=4.615 $Y=1.53 $X2=0 $Y2=0
cc_333 N_A_112_47#_c_361_n N_X_c_715_n 0.0141442f $X=4.785 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_112_47#_c_362_n N_X_c_715_n 0.0141481f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_112_47#_c_355_n N_X_c_716_n 0.020996f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A_112_47#_c_362_n N_X_c_716_n 0.0121906f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_112_47#_c_354_n N_X_c_718_n 0.00531018f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_112_47#_c_355_n N_X_c_718_n 0.0175841f $X=5.36 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_112_47#_c_362_n N_X_c_718_n 0.0214614f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_112_47#_c_364_n N_X_c_718_n 0.00224391f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_112_47#_M1010_g X 7.03718e-19 $X=4.94 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_112_47#_M1017_g X 0.0161546f $X=5.36 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A_112_47#_c_371_n X 0.00742871f $X=4.615 $Y=1.53 $X2=0 $Y2=0
cc_344 N_A_112_47#_c_360_n X 0.00189058f $X=4.7 $Y=1.445 $X2=0 $Y2=0
cc_345 N_A_112_47#_c_362_n X 0.0181901f $X=5.11 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_112_47#_c_364_n X 0.00222985f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_112_47#_c_357_n N_VGND_M1011_d 6.44201e-19 $X=0.53 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_348 N_A_112_47#_c_358_n N_VGND_M1011_d 0.00301785f $X=0.29 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_349 N_A_112_47#_c_359_n N_VGND_M1016_d 0.00162089f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_350 N_A_112_47#_c_358_n N_VGND_c_766_n 0.00114168f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_351 N_A_112_47#_c_357_n N_VGND_c_767_n 0.00491543f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_352 N_A_112_47#_c_358_n N_VGND_c_767_n 0.00856149f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_353 N_A_112_47#_c_359_n N_VGND_c_768_n 0.0118049f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_354 N_A_112_47#_c_354_n N_VGND_c_771_n 0.00316354f $X=4.94 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A_112_47#_c_355_n N_VGND_c_772_n 0.00316354f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_356 N_A_112_47#_c_357_n N_VGND_c_773_n 0.00198695f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_357 N_A_112_47#_c_387_n N_VGND_c_773_n 0.0188551f $X=0.695 $Y=0.39 $X2=0
+ $Y2=0
cc_358 N_A_112_47#_c_359_n N_VGND_c_773_n 0.00198695f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_359 N_A_112_47#_c_359_n N_VGND_c_775_n 0.00198695f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_360 N_A_112_47#_c_392_n N_VGND_c_775_n 0.0188551f $X=1.535 $Y=0.39 $X2=0
+ $Y2=0
cc_361 N_A_112_47#_c_354_n N_VGND_c_781_n 0.00435566f $X=4.94 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A_112_47#_c_355_n N_VGND_c_781_n 0.00435457f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_112_47#_M1011_s N_VGND_c_784_n 0.00215201f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_364 N_A_112_47#_M1009_d N_VGND_c_784_n 0.00215201f $X=1.4 $Y=0.235 $X2=0
+ $Y2=0
cc_365 N_A_112_47#_c_354_n N_VGND_c_784_n 0.0072173f $X=4.94 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_112_47#_c_355_n N_VGND_c_784_n 0.00695947f $X=5.36 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_112_47#_c_357_n N_VGND_c_784_n 0.00412013f $X=0.53 $Y=0.815 $X2=0
+ $Y2=0
cc_368 N_A_112_47#_c_358_n N_VGND_c_784_n 0.0024413f $X=0.29 $Y=0.815 $X2=0
+ $Y2=0
cc_369 N_A_112_47#_c_387_n N_VGND_c_784_n 0.0122069f $X=0.695 $Y=0.39 $X2=0
+ $Y2=0
cc_370 N_A_112_47#_c_359_n N_VGND_c_784_n 0.00835832f $X=1.37 $Y=0.815 $X2=0
+ $Y2=0
cc_371 N_A_112_47#_c_392_n N_VGND_c_784_n 0.0122069f $X=1.535 $Y=0.39 $X2=0
+ $Y2=0
cc_372 N_A_112_47#_c_392_n N_A_470_47#_c_865_n 0.00508738f $X=1.535 $Y=0.39
+ $X2=0 $Y2=0
cc_373 N_A_112_47#_c_371_n N_A_470_47#_c_866_n 0.0027094f $X=4.615 $Y=1.53 $X2=0
+ $Y2=0
cc_374 N_A_112_47#_c_359_n N_A_470_47#_c_867_n 0.00606598f $X=1.37 $Y=0.815
+ $X2=0 $Y2=0
cc_375 N_A_27_297#_c_527_n N_VPWR_M1004_d 2.19468e-19 $X=1.005 $Y=2.21 $X2=-0.19
+ $Y2=1.305
cc_376 N_A_27_297#_c_527_n N_VPWR_c_580_n 0.0132731f $X=1.005 $Y=2.21 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_523_n N_VPWR_c_580_n 3.62989e-19 $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_524_n N_VPWR_c_580_n 0.00503766f $X=0.23 $Y=2.21 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_530_n N_VPWR_c_580_n 3.7344e-19 $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_554_n N_VPWR_c_580_n 0.00502875f $X=1.15 $Y=2.21 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_531_n N_VPWR_c_583_n 0.0330174f $X=1.83 $Y=2.38 $X2=0 $Y2=0
cc_382 N_A_27_297#_c_546_n N_VPWR_c_583_n 0.0151213f $X=1.955 $Y=2.3 $X2=0 $Y2=0
cc_383 N_A_27_297#_c_527_n N_VPWR_c_583_n 8.18583e-19 $X=1.005 $Y=2.21 $X2=0
+ $Y2=0
cc_384 N_A_27_297#_c_554_n N_VPWR_c_583_n 0.0137704f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_527_n N_VPWR_c_585_n 8.25414e-19 $X=1.005 $Y=2.21 $X2=0
+ $Y2=0
cc_386 N_A_27_297#_c_523_n N_VPWR_c_585_n 3.6232e-19 $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_387 N_A_27_297#_c_524_n N_VPWR_c_585_n 0.0172358f $X=0.23 $Y=2.21 $X2=0 $Y2=0
cc_388 N_A_27_297#_M1004_s N_VPWR_c_579_n 0.00119537f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_389 N_A_27_297#_M1019_s N_VPWR_c_579_n 0.00115087f $X=0.98 $Y=1.485 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_M1014_d N_VPWR_c_579_n 0.00207714f $X=1.82 $Y=1.485 $X2=0
+ $Y2=0
cc_391 N_A_27_297#_c_531_n N_VPWR_c_579_n 0.0190921f $X=1.83 $Y=2.38 $X2=0 $Y2=0
cc_392 N_A_27_297#_c_546_n N_VPWR_c_579_n 0.00938089f $X=1.955 $Y=2.3 $X2=0
+ $Y2=0
cc_393 N_A_27_297#_c_527_n N_VPWR_c_579_n 0.0519284f $X=1.005 $Y=2.21 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_523_n N_VPWR_c_579_n 0.0285979f $X=0.375 $Y=2.21 $X2=0
+ $Y2=0
cc_395 N_A_27_297#_c_524_n N_VPWR_c_579_n 0.00254937f $X=0.23 $Y=2.21 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_530_n N_VPWR_c_579_n 0.0281673f $X=1.15 $Y=2.21 $X2=0 $Y2=0
cc_397 N_A_27_297#_c_554_n N_VPWR_c_579_n 0.00227213f $X=1.15 $Y=2.21 $X2=0
+ $Y2=0
cc_398 N_A_27_297#_c_546_n N_A_470_297#_c_668_n 0.0230175f $X=1.955 $Y=2.3 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_579_n N_A_470_297#_M1000_d 0.00213528f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_400 N_VPWR_c_579_n N_A_470_297#_M1002_d 0.00223619f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_579_n N_A_470_297#_M1006_d 0.00214355f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_579_n N_A_470_297#_M1010_d 0.00209344f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_579_n N_A_470_297#_M1017_d 0.00295147f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_M1000_s N_A_470_297#_c_670_n 0.00317795f $X=2.76 $Y=1.485 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_581_n N_A_470_297#_c_670_n 0.0117423f $X=2.895 $Y=2.3 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_579_n N_A_470_297#_c_670_n 0.0109496f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_586_n N_A_470_297#_c_699_n 0.0142343f $X=3.61 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_579_n N_A_470_297#_c_699_n 0.00955092f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_587_n N_A_470_297#_c_683_n 0.0159273f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_579_n N_A_470_297#_c_683_n 0.00962421f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_583_n N_A_470_297#_c_668_n 0.0201302f $X=2.77 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_579_n N_A_470_297#_c_668_n 0.0119856f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_M1003_s N_A_470_297#_c_674_n 0.00426328f $X=3.6 $Y=1.485 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_582_n N_A_470_297#_c_674_n 0.0158823f $X=3.79 $Y=2.3 $X2=0 $Y2=0
cc_415 N_VPWR_c_579_n N_A_470_297#_c_674_n 0.0111506f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_587_n N_A_470_297#_c_669_n 0.0839273f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_579_n N_A_470_297#_c_669_n 0.0501007f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_579_n N_X_M1010_s 0.00216833f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_419 N_A_470_297#_c_683_n N_X_M1010_s 0.00312348f $X=5.445 $Y=2.38 $X2=0 $Y2=0
cc_420 N_A_470_297#_M1017_d X 0.00375273f $X=5.435 $Y=1.485 $X2=0 $Y2=0
cc_421 N_A_470_297#_c_683_n X 0.00326218f $X=5.445 $Y=2.38 $X2=0 $Y2=0
cc_422 N_A_470_297#_c_713_p X 0.0166517f $X=5.57 $Y=1.96 $X2=0 $Y2=0
cc_423 N_A_470_297#_c_683_n N_X_c_748_n 0.0116103f $X=5.445 $Y=2.38 $X2=0 $Y2=0
cc_424 N_X_c_715_n N_VGND_M1007_s 0.00315681f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_425 N_X_c_718_n N_VGND_M1008_s 0.00326492f $X=5.15 $Y=0.73 $X2=0 $Y2=0
cc_426 N_X_c_715_n N_VGND_c_771_n 0.0127273f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_427 N_X_c_718_n N_VGND_c_772_n 0.0140244f $X=5.15 $Y=0.73 $X2=0 $Y2=0
cc_428 N_X_c_715_n N_VGND_c_779_n 0.00401766f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_429 N_X_c_715_n N_VGND_c_781_n 0.00198695f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_430 N_X_c_718_n N_VGND_c_781_n 0.00681853f $X=5.15 $Y=0.73 $X2=0 $Y2=0
cc_431 N_X_c_718_n N_VGND_c_783_n 0.00404417f $X=5.15 $Y=0.73 $X2=0 $Y2=0
cc_432 N_X_M1001_d N_VGND_c_784_n 0.00261003f $X=3.6 $Y=0.235 $X2=0 $Y2=0
cc_433 N_X_M1007_d N_VGND_c_784_n 0.0031882f $X=5.015 $Y=0.235 $X2=0 $Y2=0
cc_434 N_X_c_715_n N_VGND_c_784_n 0.0125287f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_435 N_X_c_718_n N_VGND_c_784_n 0.0205273f $X=5.15 $Y=0.73 $X2=0 $Y2=0
cc_436 N_X_c_715_n N_A_470_47#_M1018_s 0.00319929f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_437 N_X_c_717_n N_A_470_47#_c_866_n 0.00138158f $X=3.955 $Y=0.775 $X2=0 $Y2=0
cc_438 N_X_M1001_d N_A_470_47#_c_868_n 0.00408566f $X=3.6 $Y=0.235 $X2=0 $Y2=0
cc_439 N_X_c_715_n N_A_470_47#_c_868_n 0.0180755f $X=4.985 $Y=0.815 $X2=0 $Y2=0
cc_440 N_X_c_717_n N_A_470_47#_c_868_n 0.0170874f $X=3.955 $Y=0.775 $X2=0 $Y2=0
cc_441 N_VGND_c_784_n N_A_470_47#_M1005_s 0.00209319f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_442 N_VGND_c_784_n N_A_470_47#_M1012_s 0.00216812f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_784_n N_A_470_47#_M1018_s 0.00209344f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_769_n N_A_470_47#_c_865_n 0.0168055f $X=1.955 $Y=0.39 $X2=0
+ $Y2=0
cc_445 N_VGND_c_777_n N_A_470_47#_c_865_n 0.0209752f $X=2.81 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_784_n N_A_470_47#_c_865_n 0.0124119f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_M1005_d N_A_470_47#_c_866_n 0.00162089f $X=2.76 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_VGND_c_770_n N_A_470_47#_c_866_n 0.0118745f $X=2.895 $Y=0.39 $X2=0
+ $Y2=0
cc_449 N_VGND_c_777_n N_A_470_47#_c_866_n 0.00198695f $X=2.81 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_779_n N_A_470_47#_c_866_n 0.00198695f $X=4.645 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_784_n N_A_470_47#_c_866_n 0.00835832f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_779_n N_A_470_47#_c_880_n 0.0152433f $X=4.645 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_784_n N_A_470_47#_c_880_n 0.00947934f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_771_n N_A_470_47#_c_868_n 0.0131818f $X=4.73 $Y=0.39 $X2=0 $Y2=0
cc_455 N_VGND_c_779_n N_A_470_47#_c_868_n 0.0561952f $X=4.645 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_784_n N_A_470_47#_c_868_n 0.035263f $X=5.75 $Y=0 $X2=0 $Y2=0

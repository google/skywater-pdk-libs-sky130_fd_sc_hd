* File: sky130_fd_sc_hd__a21oi_1.spice
* Created: Tue Sep  1 18:52:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a21oi_1.pex.spice"
.subckt sky130_fd_sc_hd__a21oi_1  VNB VPB B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_B1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1005 A_199_47# N_A1_M1005_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65 AD=0.095875
+ AS=0.091 PD=0.945 PS=0.93 NRD=17.076 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_199_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.095875 PD=1.83 PS=0.945 NRD=0 NRS=17.076 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_113_297#_M1002_d N_B1_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_113_297#_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.1475 AS=0.14 PD=1.295 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_A_113_297#_M1000_d N_A2_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.1475 PD=2.53 PS=1.295 NRD=0 NRS=2.9353 M=1 R=6.66667 SA=75001.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.5631 P=7.65
*
.include "sky130_fd_sc_hd__a21oi_1.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_hd__sdfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=2.5698e+12p ps=2.353e+07u
M1001 a_1888_21# a_1714_47# a_2004_47# VNB nshort w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=4.158e+11p ps=3.99e+06u
M1002 Q_N a_1888_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1003 a_1823_47# a_193_47# a_1714_47# VNB nshort w=360000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=1.422e+11p ps=1.51e+06u
M1004 a_2004_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.5604e+12p ps=1.671e+07u
M1005 VPWR a_2696_47# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 a_381_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_1888_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.457e+11p pd=2.34e+06u as=0p ps=0u
M1008 a_1714_47# a_27_47# a_1619_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1009 VGND RESET_B a_1401_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1010 a_1017_413# a_193_47# a_931_47# VPB phighvt w=420000u l=150000u
+  ad=1.89e+11p pd=1.74e+06u as=1.134e+11p ps=1.38e+06u
M1011 a_1107_21# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.94e+11p pd=2.46e+06u as=0p ps=0u
M1012 a_453_47# SCE a_381_47# VNB nshort w=420000u l=150000u
+  ad=2.412e+11p pd=2.85e+06u as=0p ps=0u
M1013 VGND SCE a_423_315# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1014 a_1251_47# a_1401_21# a_1107_21# VNB nshort w=640000u l=150000u
+  ad=3.6e+11p pd=3.74e+06u as=1.728e+11p ps=1.82e+06u
M1015 Q a_2696_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1016 a_1107_21# a_931_47# a_1251_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_2004_47# a_1401_21# a_1888_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_2696_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_453_47# D a_752_413# VPB phighvt w=420000u l=150000u
+  ad=3.071e+11p pd=3.31e+06u as=1.134e+11p ps=1.38e+06u
M1020 a_1041_47# a_27_47# a_931_47# VNB nshort w=360000u l=150000u
+  ad=1.341e+11p pd=1.5e+06u as=1.44e+11p ps=1.52e+06u
M1021 a_1800_413# a_27_47# a_1714_47# VPB phighvt w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=1.134e+11p ps=1.38e+06u
M1022 a_752_413# SCE VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_764_47# a_423_315# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1024 a_453_47# D a_764_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_2122_329# a_1714_47# a_1888_21# VPB phighvt w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1026 VGND a_2696_47# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR CLK_N a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1028 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1029 VPWR a_1401_21# a_2122_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR RESET_B a_1401_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1031 VPWR a_1401_21# a_1351_329# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1032 a_1714_47# a_193_47# a_1572_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.486e+11p ps=2.82e+06u
M1033 VPWR a_1888_21# a_2696_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1034 a_381_363# SCD VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1035 VPWR SCE a_423_315# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1036 VPWR a_1107_21# a_1017_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1351_329# a_931_47# a_1107_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VGND a_1107_21# a_1041_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_453_47# a_423_315# a_381_363# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_931_47# a_27_47# a_453_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1619_47# a_1107_21# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VGND a_1888_21# a_1823_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_1888_21# a_1800_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VGND a_1888_21# a_2696_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1045 a_931_47# a_193_47# a_453_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_1888_21# Q_N VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1251_47# SET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 VGND CLK_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1049 VGND a_1888_21# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1050 a_1572_329# a_1107_21# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 Q_N a_1888_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__mux4_1.pex.spice
* Created: Thu Aug 27 14:28:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX4_1%A1 3 7 9 10 14 15
c30 14 0 1.84785e-19 $X=0.41 $Y=1.16
r31 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r32 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r33 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r34 9 10 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.322 $Y=1.19
+ $X2=0.322 $Y2=1.53
r35 9 15 1.00212 $w=3.43e-07 $l=3e-08 $layer=LI1_cond $X=0.322 $Y=1.19 $X2=0.322
+ $Y2=1.16
r36 7 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r37 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A0 3 7 9 10 14 15
c38 14 0 9.32549e-20 $X=0.89 $Y=1.16
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r40 9 10 9.0076 $w=4.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.022 $Y=1.19
+ $X2=1.022 $Y2=1.53
r41 9 15 0.794788 $w=4.33e-07 $l=3e-08 $layer=LI1_cond $X=1.022 $Y=1.19
+ $X2=1.022 $Y2=1.16
r42 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r43 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=2.275
r44 1 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r45 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_247_21# 1 2 9 11 12 15 19 21 24 26 29 33 35
+ 36 39 42 46 48 52 53
c162 53 0 1.11083e-19 $X=4.24 $Y=1.18
c163 46 0 3.23144e-19 $X=2.245 $Y=1.2
c164 35 0 1.82348e-19 $X=4.23 $Y=1.19
r165 52 54 61.7949 $w=2.34e-07 $l=3e-07 $layer=POLY_cond $X=4.24 $Y=1.185
+ $X2=4.54 $Y2=1.185
r166 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.24
+ $Y=1.18 $X2=4.24 $Y2=1.18
r167 50 52 29.8675 $w=2.34e-07 $l=1.45e-07 $layer=POLY_cond $X=4.095 $Y=1.185
+ $X2=4.24 $Y2=1.185
r168 47 56 7.29755 $w=3.26e-07 $l=2.64953e-07 $layer=LI1_cond $X=2.245 $Y=1.2
+ $X2=2.44 $Y2=1.365
r169 46 48 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.2
+ $X2=2.08 $Y2=1.2
r170 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.245
+ $Y=1.2 $X2=2.245 $Y2=1.2
r171 42 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.375 $Y=1.19
+ $X2=4.375 $Y2=1.19
r172 39 56 3.55521 $w=3.26e-07 $l=9.5e-08 $layer=LI1_cond $X=2.535 $Y=1.365
+ $X2=2.44 $Y2=1.365
r173 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.19
+ $X2=2.535 $Y2=1.19
r174 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.19
+ $X2=2.535 $Y2=1.19
r175 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.23 $Y=1.19
+ $X2=4.375 $Y2=1.19
r176 35 36 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=4.23 $Y=1.19
+ $X2=2.68 $Y2=1.19
r177 31 39 13.2853 $w=3.26e-07 $l=4.67253e-07 $layer=LI1_cond $X=2.89 $Y=1.625
+ $X2=2.535 $Y2=1.365
r178 31 33 22.2257 $w=3.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.89 $Y=1.625
+ $X2=2.89 $Y2=2.3
r179 27 56 0.102097 $w=3.6e-07 $l=2.6e-07 $layer=LI1_cond $X=2.44 $Y=1.105
+ $X2=2.44 $Y2=1.365
r180 27 29 16.3263 $w=3.58e-07 $l=5.1e-07 $layer=LI1_cond $X=2.44 $Y=1.105
+ $X2=2.44 $Y2=0.595
r181 22 54 13.1928 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.54 $Y=1.325
+ $X2=4.54 $Y2=1.185
r182 22 24 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.54 $Y=1.325
+ $X2=4.54 $Y2=2.025
r183 19 50 13.1928 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.095 $Y=1.045
+ $X2=4.095 $Y2=1.185
r184 19 21 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.095 $Y=1.045
+ $X2=4.095 $Y2=0.695
r185 18 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.26
+ $X2=1.83 $Y2=1.26
r186 18 48 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.905 $Y=1.26
+ $X2=2.08 $Y2=1.26
r187 13 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=1.26
r188 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.335
+ $X2=1.83 $Y2=2.025
r189 11 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=1.26
+ $X2=1.83 $Y2=1.26
r190 11 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.755 $Y=1.26
+ $X2=1.385 $Y2=1.26
r191 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.31 $Y=1.185
+ $X2=1.385 $Y2=1.26
r192 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.31 $Y=1.185
+ $X2=1.31 $Y2=0.445
r193 2 33 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=2.155 $X2=2.98 $Y2=2.3
r194 1 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.45 $X2=2.525 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%S0 3 5 6 7 9 10 11 15 16 18 20 22 24 25 27 31
+ 32 33 38
c107 38 0 1.80869e-19 $X=3.415 $Y=1.18
c108 20 0 1.30364e-19 $X=4.045 $Y=1.665
c109 16 0 1.57897e-19 $X=3.19 $Y=1.74
r110 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.18 $X2=3.415 $Y2=1.18
r111 32 33 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=3.415 $Y2=1.87
r112 32 38 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=3.415 $Y2=1.18
r113 31 37 28.8521 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.6 $Y=1.18
+ $X2=3.415 $Y2=1.18
r114 29 37 29.6319 $w=3.7e-07 $l=1.9e-07 $layer=POLY_cond $X=3.225 $Y=1.18
+ $X2=3.415 $Y2=1.18
r115 29 30 40.7976 $w=5.73e-07 $l=4.85e-07 $layer=POLY_cond $X=2.962 $Y=1.18
+ $X2=2.962 $Y2=1.665
r116 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.12 $Y=1.74
+ $X2=4.12 $Y2=2.025
r117 22 31 33.737 $w=3.7e-07 $l=2.19317e-07 $layer=POLY_cond $X=3.675 $Y=0.995
+ $X2=3.6 $Y2=1.18
r118 22 24 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.675 $Y=0.995 $X2=3.675
+ $Y2=0.695
r119 21 30 34.8849 $w=1.5e-07 $l=3.03e-07 $layer=POLY_cond $X=3.265 $Y=1.665
+ $X2=2.962 $Y2=1.665
r120 20 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.045 $Y=1.665
+ $X2=4.12 $Y2=1.74
r121 20 21 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=4.045 $Y=1.665
+ $X2=3.265 $Y2=1.665
r122 16 30 36.2869 $w=5.73e-07 $l=2.62838e-07 $layer=POLY_cond $X=3.19 $Y=1.74
+ $X2=2.962 $Y2=1.665
r123 16 18 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.19 $Y=1.74
+ $X2=3.19 $Y2=2.275
r124 13 29 45.54 $w=5.73e-07 $l=3.05817e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.962 $Y2=1.18
r125 13 15 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.735 $Y=0.995
+ $X2=2.735 $Y2=0.66
r126 12 15 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.735 $Y=0.255
+ $X2=2.735 $Y2=0.66
r127 10 30 34.8849 $w=1.5e-07 $l=3.02e-07 $layer=POLY_cond $X=2.66 $Y=1.665
+ $X2=2.962 $Y2=1.665
r128 10 11 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.66 $Y=1.665
+ $X2=2.325 $Y2=1.665
r129 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.25 $Y=1.74
+ $X2=2.325 $Y2=1.665
r130 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.25 $Y=1.74 $X2=2.25
+ $Y2=2.025
r131 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.66 $Y=0.18
+ $X2=2.735 $Y2=0.255
r132 5 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.66 $Y=0.18 $X2=1.87
+ $Y2=0.18
r133 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.795 $Y=0.255
+ $X2=1.87 $Y2=0.18
r134 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.795 $Y=0.255
+ $X2=1.795 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A3 3 7 9 10 14
c48 14 0 3.26131e-20 $X=4.96 $Y=1.22
c49 3 0 1.52475e-19 $X=5.015 $Y=2.275
r50 14 17 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.987 $Y=1.22
+ $X2=4.987 $Y2=1.385
r51 14 16 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.987 $Y=1.22
+ $X2=4.987 $Y2=1.055
r52 9 10 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=4.922 $Y=1.19
+ $X2=4.922 $Y2=1.53
r53 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.96
+ $Y=1.22 $X2=4.96 $Y2=1.22
r54 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.025 $Y=0.445
+ $X2=5.025 $Y2=1.055
r55 3 17 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.015 $Y=2.275
+ $X2=5.015 $Y2=1.385
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A2 3 7 9 12 13
r42 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.495 $Y=1.22
+ $X2=5.495 $Y2=1.385
r43 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.495 $Y=1.22
+ $X2=5.495 $Y2=1.055
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.22 $X2=5.495 $Y2=1.22
r45 9 13 2.41145 $w=6.18e-07 $l=1.25e-07 $layer=LI1_cond $X=5.37 $Y=1.365
+ $X2=5.495 $Y2=1.365
r46 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.445 $Y=0.445
+ $X2=5.445 $Y2=1.055
r47 3 15 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.435 $Y=2.275
+ $X2=5.435 $Y2=1.385
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%S1 3 7 9 13 17 19 20 28
c80 20 0 3.25148e-20 $X=6.26 $Y=1.19
r81 27 28 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.385 $Y=1.16
+ $X2=6.46 $Y2=1.16
r82 26 27 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.375 $Y=1.16
+ $X2=6.385 $Y2=1.16
r83 23 26 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.14 $Y=1.16
+ $X2=6.375 $Y2=1.16
r84 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.14
+ $Y=1.16 $X2=6.14 $Y2=1.16
r85 20 24 2.11073 $w=6.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.26 $Y=1.335
+ $X2=6.14 $Y2=1.335
r86 15 19 36.6911 $w=1.5e-07 $l=1.64481e-07 $layer=POLY_cond $X=7.325 $Y=1
+ $X2=7.32 $Y2=1.162
r87 15 17 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=7.325 $Y=1
+ $X2=7.325 $Y2=0.445
r88 11 19 36.6911 $w=1.5e-07 $l=1.65481e-07 $layer=POLY_cond $X=7.315 $Y=1.325
+ $X2=7.32 $Y2=1.162
r89 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.315 $Y=1.325
+ $X2=7.315 $Y2=2.275
r90 9 19 4.85217 $w=3.25e-07 $l=8e-08 $layer=POLY_cond $X=7.24 $Y=1.162 $X2=7.32
+ $Y2=1.162
r91 9 28 138.49 $w=3.25e-07 $l=7.8e-07 $layer=POLY_cond $X=7.24 $Y=1.162
+ $X2=6.46 $Y2=1.162
r92 5 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.385 $Y=0.995
+ $X2=6.385 $Y2=1.16
r93 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.385 $Y=0.995
+ $X2=6.385 $Y2=0.445
r94 1 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.375 $Y=1.325
+ $X2=6.375 $Y2=1.16
r95 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.375 $Y=1.325
+ $X2=6.375 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_1290_413# 1 2 9 11 13 14 18 22 23 26 29 30
+ 33 36 37 40
c100 37 0 5.58442e-20 $X=8.56 $Y=1.19
r101 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.355
+ $Y=1.19 $X2=8.355 $Y2=1.19
r102 37 41 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.56 $Y=1.19
+ $X2=8.355 $Y2=1.19
r103 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.56 $Y=1.19
+ $X2=8.56 $Y2=1.19
r104 33 47 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.72 $Y=1.19
+ $X2=6.6 $Y2=1.19
r105 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.72 $Y=1.19
+ $X2=6.72 $Y2=1.19
r106 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.865 $Y=1.19
+ $X2=6.72 $Y2=1.19
r107 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.415 $Y=1.19
+ $X2=8.56 $Y2=1.19
r108 29 30 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=8.415 $Y=1.19
+ $X2=6.865 $Y2=1.19
r109 26 28 10.4571 $w=1.73e-07 $l=1.65e-07 $layer=LI1_cond $X=6.597 $Y=0.49
+ $X2=6.597 $Y2=0.655
r110 22 23 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=6.592 $Y=2.3
+ $X2=6.592 $Y2=2.135
r111 19 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=1.275
+ $X2=6.6 $Y2=1.19
r112 19 23 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=6.6 $Y=1.275 $X2=6.6
+ $Y2=2.135
r113 18 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=1.105
+ $X2=6.6 $Y2=1.19
r114 18 28 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.6 $Y=1.105
+ $X2=6.6 $Y2=0.655
r115 15 16 73.5684 $w=1.9e-07 $l=2.9e-07 $layer=POLY_cond $X=7.8 $Y=1.19
+ $X2=8.09 $Y2=1.19
r116 14 40 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=8.165 $Y=1.19
+ $X2=8.355 $Y2=1.19
r117 14 16 17.6794 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=8.165 $Y=1.19
+ $X2=8.09 $Y2=1.19
r118 11 16 8.39207 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.09 $Y=1.055
+ $X2=8.09 $Y2=1.19
r119 11 13 115.68 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.09 $Y=1.055
+ $X2=8.09 $Y2=0.695
r120 7 15 8.39207 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.8 $Y=1.325
+ $X2=7.8 $Y2=1.19
r121 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=7.8 $Y=1.325 $X2=7.8
+ $Y2=2.04
r122 2 22 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=6.45
+ $Y=2.065 $X2=6.585 $Y2=2.3
r123 1 26 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=6.46
+ $Y=0.235 $X2=6.595 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_1478_413# 1 2 9 12 14 16 19 21 22 23 24 25
+ 29 30 34 37 40
c95 23 0 6.48099e-20 $X=8.645 $Y=1.75
r96 32 34 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=7.525 $Y=2.36
+ $X2=7.69 $Y2=2.36
r97 30 41 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.16
+ $X2=9.08 $Y2=1.325
r98 30 40 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.16
+ $X2=9.08 $Y2=0.995
r99 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.04
+ $Y=1.16 $X2=9.04 $Y2=1.16
r100 27 29 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=9.04 $Y=1.665
+ $X2=9.04 $Y2=1.16
r101 26 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.04 $Y=0.885
+ $X2=9.04 $Y2=1.16
r102 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.955 $Y=0.8
+ $X2=9.04 $Y2=0.885
r103 24 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.955 $Y=0.8
+ $X2=8.725 $Y2=0.8
r104 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.955 $Y=1.75
+ $X2=9.04 $Y2=1.665
r105 22 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.955 $Y=1.75
+ $X2=8.645 $Y2=1.75
r106 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.64 $Y=0.715
+ $X2=8.725 $Y2=0.8
r107 20 21 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.64 $Y=0.425
+ $X2=8.64 $Y2=0.715
r108 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.56 $Y=1.835
+ $X2=8.645 $Y2=1.75
r109 18 19 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.56 $Y=1.835
+ $X2=8.56 $Y2=2.295
r110 17 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=0.34
+ $X2=7.815 $Y2=0.34
r111 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.555 $Y=0.34
+ $X2=8.64 $Y2=0.425
r112 16 17 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.555 $Y=0.34
+ $X2=7.9 $Y2=0.34
r113 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=2.38
+ $X2=8.56 $Y2=2.295
r114 14 34 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.475 $Y=2.38
+ $X2=7.69 $Y2=2.38
r115 12 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.19 $Y=1.985
+ $X2=9.19 $Y2=1.325
r116 9 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.19 $Y=0.56
+ $X2=9.19 $Y2=0.995
r117 2 32 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.39
+ $Y=2.065 $X2=7.525 $Y2=2.34
r118 1 37 182 $w=1.7e-07 $l=4.98999e-07 $layer=licon1_NDIFF $count=1 $X=7.4
+ $Y=0.235 $X2=7.815 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_27_413# 1 2 9 11 12 15
c31 11 0 1.84785e-19 $X=1.535 $Y=1.88
r32 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=1.88
+ $X2=1.62 $Y2=1.88
r33 11 12 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=1.535 $Y=1.88
+ $X2=0.345 $Y2=1.88
r34 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.965
+ $X2=0.345 $Y2=1.88
r35 7 9 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=1.965
+ $X2=0.26 $Y2=2.3
r36 2 15 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.815 $X2=1.62 $Y2=1.96
r37 1 9 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%VPWR 1 2 3 4 5 18 22 26 30 34 36 38 43 51 59
+ 64 74 75 78 81 84 87 90
r115 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r116 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r117 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 75 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r121 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r122 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=8.98 $Y2=2.72
r123 72 74 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.145 $Y=2.72
+ $X2=9.43 $Y2=2.72
r124 71 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r125 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r126 68 71 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r127 68 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r128 67 70 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r129 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r130 65 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=6.155 $Y2=2.72
r131 65 67 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.33 $Y=2.72
+ $X2=6.67 $Y2=2.72
r132 64 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.815 $Y=2.72
+ $X2=8.98 $Y2=2.72
r133 64 70 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.815 $Y=2.72
+ $X2=8.51 $Y2=2.72
r134 63 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r135 63 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r136 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.39 $Y=2.72
+ $X2=5.225 $Y2=2.72
r138 60 62 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.39 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 59 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.98 $Y=2.72
+ $X2=6.155 $Y2=2.72
r140 59 62 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.98 $Y=2.72
+ $X2=5.75 $Y2=2.72
r141 58 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r142 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r143 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 55 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r145 54 57 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=2.72
+ $X2=3.4 $Y2=2.72
r148 52 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.565 $Y=2.72
+ $X2=3.91 $Y2=2.72
r149 51 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=5.225 $Y2=2.72
r150 51 57 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 50 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r152 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r153 47 50 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r154 47 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 46 49 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r156 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r157 44 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r158 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r159 43 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=2.72
+ $X2=3.4 $Y2=2.72
r160 43 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.235 $Y=2.72
+ $X2=2.99 $Y2=2.72
r161 38 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r162 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r163 36 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r164 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r165 32 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=8.98 $Y2=2.72
r166 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=2.635
+ $X2=8.98 $Y2=2.34
r167 28 87 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=2.635
+ $X2=6.155 $Y2=2.72
r168 28 30 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.155 $Y=2.635
+ $X2=6.155 $Y2=2.34
r169 24 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=2.635
+ $X2=5.225 $Y2=2.72
r170 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=2.635
+ $X2=5.225 $Y2=2.34
r171 20 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=2.635 $X2=3.4
+ $Y2=2.72
r172 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.4 $Y=2.635
+ $X2=3.4 $Y2=2.34
r173 16 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r174 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r175 5 34 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=8.855
+ $Y=1.485 $X2=8.98 $Y2=2.34
r176 4 30 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=2.065 $X2=6.165 $Y2=2.34
r177 3 26 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=2.065 $X2=5.225 $Y2=2.34
r178 2 22 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=2.065 $X2=3.4 $Y2=2.34
r179 1 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_193_413# 1 2 7 11 14
c23 11 0 7.11638e-20 $X=2.46 $Y=1.96
c24 7 0 3.23044e-20 $X=2.375 $Y=2.38
r25 9 11 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.46 $Y=2.295
+ $X2=2.46 $Y2=1.96
r26 8 14 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.185 $Y=2.38
+ $X2=1.1 $Y2=2.3
r27 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=2.46 $Y2=2.295
r28 7 8 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=1.185 $Y2=2.38
r29 2 11 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.815 $X2=2.46 $Y2=1.96
r30 1 14 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=2.065 $X2=1.1 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_277_47# 1 2 3 4 13 14 15 16 18 23 26 27 29
+ 30 31 32 39 41 42
c166 41 0 5.58442e-20 $X=8.055 $Y=0.85
c167 27 0 3.25148e-20 $X=7.085 $Y=2.135
c168 23 0 6.41913e-20 $X=2.04 $Y=2.04
c169 16 0 3.23044e-20 $X=1.58 $Y=1.54
c170 15 0 1.57897e-19 $X=1.875 $Y=1.54
c171 14 0 9.32549e-20 $X=1.495 $Y=1.455
r172 42 51 12.4025 $w=2.41e-07 $l=2.45e-07 $layer=LI1_cond $X=8.055 $Y=0.765
+ $X2=8.3 $Y2=0.765
r173 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.055 $Y=0.85
+ $X2=8.055 $Y2=0.85
r174 39 48 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=7.1 $Y=0.85 $X2=7.1
+ $Y2=0.935
r175 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.135 $Y=0.85
+ $X2=7.135 $Y2=0.85
r176 34 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=0.85
+ $X2=1.615 $Y2=0.85
r177 32 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.28 $Y=0.85
+ $X2=7.135 $Y2=0.85
r178 31 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.91 $Y=0.85
+ $X2=8.055 $Y2=0.85
r179 31 32 0.779701 $w=1.4e-07 $l=6.3e-07 $layer=MET1_cond $X=7.91 $Y=0.85
+ $X2=7.28 $Y2=0.85
r180 30 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=0.85
+ $X2=1.615 $Y2=0.85
r181 29 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.99 $Y=0.85
+ $X2=7.135 $Y2=0.85
r182 29 30 6.47276 $w=1.4e-07 $l=5.23e-06 $layer=MET1_cond $X=6.99 $Y=0.85
+ $X2=1.76 $Y2=0.85
r183 27 48 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=7.065 $Y=2.135
+ $X2=7.065 $Y2=0.935
r184 26 27 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=2.3
+ $X2=7.085 $Y2=2.135
r185 18 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=1.955
+ $X2=1.96 $Y2=2.04
r186 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.96 $Y=1.625
+ $X2=1.96 $Y2=1.955
r187 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.875 $Y=1.54
+ $X2=1.96 $Y2=1.625
r188 15 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.875 $Y=1.54
+ $X2=1.58 $Y2=1.54
r189 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.455
+ $X2=1.58 $Y2=1.54
r190 13 45 12.4444 $w=3.15e-07 $l=2.94449e-07 $layer=LI1_cond $X=1.495 $Y=0.935
+ $X2=1.58 $Y2=0.68
r191 13 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.495 $Y=0.935
+ $X2=1.495 $Y2=1.455
r192 4 26 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.065 $X2=7.105 $Y2=2.3
r193 3 23 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.815 $X2=2.04 $Y2=2.04
r194 2 51 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=8.165
+ $Y=0.485 $X2=8.3 $Y2=0.76
r195 1 45 182 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.585 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_757_363# 1 2 9 11 12 14 15 16 19
c57 16 0 3.26131e-20 $X=4.835 $Y=2
r58 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.645 $Y=2.085
+ $X2=5.645 $Y2=2.3
r59 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.56 $Y=2
+ $X2=5.645 $Y2=2.085
r60 15 16 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.56 $Y=2 $X2=4.835
+ $Y2=2
r61 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.75 $Y=2.085
+ $X2=4.835 $Y2=2
r62 13 14 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.75 $Y=2.085
+ $X2=4.75 $Y2=2.295
r63 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.665 $Y=2.38
+ $X2=4.75 $Y2=2.295
r64 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.665 $Y=2.38
+ $X2=3.995 $Y2=2.38
r65 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.91 $Y=2.295
+ $X2=3.995 $Y2=2.38
r66 7 9 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.91 $Y=2.295
+ $X2=3.91 $Y2=1.96
r67 2 19 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=5.51
+ $Y=2.065 $X2=5.645 $Y2=2.3
r68 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.815 $X2=3.91 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_750_97# 1 2 3 4 13 14 15 16 17 20 25 28 29
+ 30 35 36 39 42
c138 15 0 1.52475e-19 $X=4.165 $Y=1.53
c139 13 0 1.29552e-19 $X=3.82 $Y=0.92
c140 4 0 6.48099e-20 $X=7.875 $Y=1.83
r141 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.64 $Y=1.87
+ $X2=7.64 $Y2=1.87
r142 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.41 $Y=1.87
+ $X2=4.41 $Y2=1.87
r143 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.555 $Y=1.87
+ $X2=4.41 $Y2=1.87
r144 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.495 $Y=1.87
+ $X2=7.64 $Y2=1.87
r145 35 36 3.63861 $w=1.4e-07 $l=2.94e-06 $layer=MET1_cond $X=7.495 $Y=1.87
+ $X2=4.555 $Y2=1.87
r146 30 43 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=7.845 $Y=1.87
+ $X2=7.64 $Y2=1.87
r147 29 33 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.01 $Y=1.87
+ $X2=8.01 $Y2=2.04
r148 29 30 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.01 $Y=1.87
+ $X2=7.845 $Y2=1.87
r149 28 43 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=7.56 $Y=1.87 $X2=7.64
+ $Y2=1.87
r150 23 39 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.33 $Y=1.615
+ $X2=4.33 $Y2=1.87
r151 20 28 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.475 $Y=1.755
+ $X2=7.56 $Y2=1.87
r152 19 20 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=7.475 $Y=0.585
+ $X2=7.475 $Y2=1.755
r153 18 25 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.2 $Y=0.5
+ $X2=7.115 $Y2=0.42
r154 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=0.5
+ $X2=7.475 $Y2=0.585
r155 17 18 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.39 $Y=0.5 $X2=7.2
+ $Y2=0.5
r156 15 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.165 $Y=1.53
+ $X2=4.33 $Y2=1.615
r157 15 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.165 $Y=1.53
+ $X2=3.905 $Y2=1.53
r158 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.82 $Y=1.445
+ $X2=3.905 $Y2=1.53
r159 13 22 8.76925 $w=3.26e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.82 $Y=0.92
+ $X2=3.885 $Y2=0.76
r160 13 14 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.82 $Y=0.92
+ $X2=3.82 $Y2=1.445
r161 4 33 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.83 $X2=8.01 $Y2=2.04
r162 3 39 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.815 $X2=4.33 $Y2=2.04
r163 2 25 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.235 $X2=7.115 $Y2=0.42
r164 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.485 $X2=3.885 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%X 1 2 7 8 9 10 16
r10 10 27 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=9.445 $Y=1.87
+ $X2=9.445 $Y2=2.3
r11 9 10 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=9.445 $Y=1.53
+ $X2=9.445 $Y2=1.87
r12 8 9 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=9.445 $Y=1.19
+ $X2=9.445 $Y2=1.53
r13 7 8 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=9.445 $Y=0.85
+ $X2=9.445 $Y2=1.19
r14 7 16 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=9.445 $Y=0.85
+ $X2=9.445 $Y2=0.42
r15 2 27 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.485 $X2=9.4 $Y2=2.3
r16 1 16 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.265
+ $Y=0.235 $X2=9.4 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_27_47# 1 2 9 11 12 15 16 19
c43 19 0 1.87789e-19 $X=2.005 $Y=0.55
c44 14 0 1.06273e-19 $X=1.1 $Y=0.635
c45 11 0 3.65312e-20 $X=1.015 $Y=0.72
r46 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.005 $Y=0.425
+ $X2=2.005 $Y2=0.55
r47 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.92 $Y=0.34
+ $X2=2.005 $Y2=0.425
r48 15 16 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.92 $Y=0.34
+ $X2=1.185 $Y2=0.34
r49 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=0.425
+ $X2=1.185 $Y2=0.34
r50 13 14 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.1 $Y=0.425 $X2=1.1
+ $Y2=0.635
r51 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=1.1 $Y2=0.635
r52 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.72
+ $X2=0.345 $Y2=0.72
r53 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r54 7 9 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=0.635 $X2=0.26
+ $Y2=0.425
r55 2 19 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.405 $X2=2.005 $Y2=0.55
r56 1 9 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 61 65 72 73 76 79 82 85 88
c123 22 0 1.29552e-19 $X=2.945 $Y=0.64
r124 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r125 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r126 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r127 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r128 73 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.97
+ $Y2=0
r129 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r130 70 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.065 $Y=0 $X2=8.98
+ $Y2=0
r131 70 72 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.065 $Y=0
+ $X2=9.43 $Y2=0
r132 69 86 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.67 $Y=0 $X2=8.97
+ $Y2=0
r133 69 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r134 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r135 66 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6.175
+ $Y2=0
r136 66 68 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=0 $X2=6.67
+ $Y2=0
r137 65 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=0 $X2=8.98
+ $Y2=0
r138 65 68 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=8.895 $Y=0
+ $X2=6.67 $Y2=0
r139 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r140 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r141 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.01 $Y=0 $X2=6.175
+ $Y2=0
r142 61 63 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.01 $Y=0 $X2=5.75
+ $Y2=0
r143 60 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r144 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r145 57 60 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.83 $Y2=0
r146 57 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r147 56 59 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r148 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r149 54 79 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=2.945
+ $Y2=0
r150 54 56 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.45
+ $Y2=0
r151 53 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r152 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r153 50 53 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r154 50 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r155 49 52 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r156 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r157 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r158 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r159 46 79 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.945
+ $Y2=0
r160 46 52 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.53
+ $Y2=0
r161 41 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r162 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r163 39 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r164 39 88 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.225 $Y2=0
r165 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r166 37 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.83
+ $Y2=0
r167 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.235
+ $Y2=0
r168 36 63 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.75
+ $Y2=0
r169 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.235
+ $Y2=0
r170 32 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0
r171 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.98 $Y=0.085
+ $X2=8.98 $Y2=0.38
r172 28 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=0.085
+ $X2=6.175 $Y2=0
r173 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.175 $Y=0.085
+ $X2=6.175 $Y2=0.38
r174 24 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0
r175 24 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0.38
r176 20 79 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r177 20 22 22.0554 $w=2.88e-07 $l=5.55e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.64
r178 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r179 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r180 5 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.855
+ $Y=0.235 $X2=8.98 $Y2=0.38
r181 4 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.05
+ $Y=0.235 $X2=6.175 $Y2=0.38
r182 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.1
+ $Y=0.235 $X2=5.235 $Y2=0.38
r183 2 22 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.45 $X2=2.945 $Y2=0.64
r184 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_668_97# 1 2 9 12 14 15
c31 15 0 1.80869e-19 $X=4.625 $Y=0.36
c32 9 0 1.29575e-19 $X=3.465 $Y=0.63
r33 14 15 10.4695 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=4.815 $Y=0.36
+ $X2=4.625 $Y2=0.36
r34 12 15 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=3.55 $Y=0.34
+ $X2=4.625 $Y2=0.34
r35 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.465 $Y=0.425
+ $X2=3.55 $Y2=0.34
r36 7 9 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.465 $Y=0.425
+ $X2=3.465 $Y2=0.63
r37 2 14 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.69
+ $Y=0.235 $X2=4.815 $Y2=0.38
r38 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.34
+ $Y=0.485 $X2=3.465 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_1%A_834_97# 1 2 7 11 14
c38 14 0 3.34925e-20 $X=4.305 $Y=0.76
r39 9 11 11.9948 $w=2.43e-07 $l=2.55e-07 $layer=LI1_cond $X=5.617 $Y=0.715
+ $X2=5.617 $Y2=0.46
r40 8 14 0.716491 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.39 $Y=0.8
+ $X2=4.305 $Y2=0.76
r41 7 9 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=5.495 $Y=0.8
+ $X2=5.617 $Y2=0.715
r42 7 8 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=5.495 $Y=0.8
+ $X2=4.39 $Y2=0.8
r43 2 11 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=5.52
+ $Y=0.235 $X2=5.655 $Y2=0.46
r44 1 14 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=4.17
+ $Y=0.485 $X2=4.305 $Y2=0.76
.ends


* File: sky130_fd_sc_hd__or2_4.spice
* Created: Tue Sep  1 19:27:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or2_4.pex.spice"
.subckt sky130_fd_sc_hd__or2_4  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1011 N_A_35_297#_M1011_d N_B_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_35_297#_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.08775 PD=1.005 PS=0.92 NRD=7.38 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_35_297#_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.115375 PD=0.92 PS=1.005 NRD=0 NRS=6.456 M=1 R=4.33333
+ SA=75001.1 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1001_d N_A_35_297#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_35_297#_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1005_d N_A_35_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 A_121_297# N_B_M1006_g N_A_35_297#_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.28 PD=1.21 PS=2.56 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_121_297# VPB PHIGHVT L=0.15 W=1 AD=0.1775
+ AS=0.105 PD=1.355 PS=1.21 NRD=7.8603 NRS=9.8303 M=1 R=6.66667 SA=75000.6
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_35_297#_M1000_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.1775 PD=1.27 PS=1.355 NRD=0 NRS=6.8753 M=1 R=6.66667 SA=75001.1
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1000_d N_A_35_297#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_35_297#_M1007_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1007_d N_A_35_297#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_251 A_121_297# 0 1.02064e-19 $X=0.605 $Y=1.485
*
.include "sky130_fd_sc_hd__or2_4.pxi.spice"
*
.ends
*
*

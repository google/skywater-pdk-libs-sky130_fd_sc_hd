* NGSPICE file created from sky130_fd_sc_hd__a41oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VPWR A4 a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=8.35e+11p pd=5.67e+06u as=1.105e+12p ps=8.21e+06u
M1001 a_428_47# A2 a_336_47# VNB nshort w=650000u l=150000u
+  ad=2.7625e+11p pd=2.15e+06u as=2.015e+11p ps=1.92e+06u
M1002 VPWR A2 a_109_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_109_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A1 a_428_47# VNB nshort w=650000u l=150000u
+  ad=4.095e+11p pd=3.86e+06u as=0p ps=0u
M1005 a_109_297# A3 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_109_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1007 a_336_47# A3 a_236_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.275e+11p ps=2e+06u
M1008 VGND B1 Y VNB nshort w=650000u l=150000u
+  ad=3.2685e+11p pd=2.35e+06u as=0p ps=0u
M1009 a_236_47# A4 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__or4bb_1.spice.SKY130_FD_SC_HD__OR4BB_1.pxi
* Created: Thu Aug 27 14:44:42 2020
* 
x_PM_SKY130_FD_SC_HD__OR4BB_1%C_N N_C_N_M1011_g N_C_N_M1008_g C_N C_N
+ N_C_N_c_93_n N_C_N_c_94_n N_C_N_c_95_n PM_SKY130_FD_SC_HD__OR4BB_1%C_N
x_PM_SKY130_FD_SC_HD__OR4BB_1%D_N N_D_N_M1009_g N_D_N_M1013_g D_N N_D_N_c_126_n
+ N_D_N_c_127_n PM_SKY130_FD_SC_HD__OR4BB_1%D_N
x_PM_SKY130_FD_SC_HD__OR4BB_1%A_205_93# N_A_205_93#_M1009_d N_A_205_93#_M1013_d
+ N_A_205_93#_M1003_g N_A_205_93#_M1005_g N_A_205_93#_c_169_n
+ N_A_205_93#_c_163_n N_A_205_93#_c_164_n N_A_205_93#_c_165_n
+ N_A_205_93#_c_166_n N_A_205_93#_c_167_n PM_SKY130_FD_SC_HD__OR4BB_1%A_205_93#
x_PM_SKY130_FD_SC_HD__OR4BB_1%A_27_410# N_A_27_410#_M1008_s N_A_27_410#_M1011_s
+ N_A_27_410#_M1006_g N_A_27_410#_M1004_g N_A_27_410#_c_234_n
+ N_A_27_410#_c_240_n N_A_27_410#_c_241_n N_A_27_410#_c_242_n
+ N_A_27_410#_c_243_n N_A_27_410#_c_244_n N_A_27_410#_c_235_n
+ N_A_27_410#_c_236_n N_A_27_410#_c_237_n N_A_27_410#_c_247_n
+ PM_SKY130_FD_SC_HD__OR4BB_1%A_27_410#
x_PM_SKY130_FD_SC_HD__OR4BB_1%B N_B_M1001_g N_B_M1007_g N_B_c_323_n N_B_c_324_n
+ B N_B_c_327_n PM_SKY130_FD_SC_HD__OR4BB_1%B
x_PM_SKY130_FD_SC_HD__OR4BB_1%A N_A_M1010_g N_A_M1012_g A N_A_c_366_n
+ N_A_c_367_n PM_SKY130_FD_SC_HD__OR4BB_1%A
x_PM_SKY130_FD_SC_HD__OR4BB_1%A_311_413# N_A_311_413#_M1003_d
+ N_A_311_413#_M1007_d N_A_311_413#_M1005_s N_A_311_413#_M1000_g
+ N_A_311_413#_M1002_g N_A_311_413#_c_416_n N_A_311_413#_c_502_p
+ N_A_311_413#_c_417_n N_A_311_413#_c_407_n N_A_311_413#_c_408_n
+ N_A_311_413#_c_418_n N_A_311_413#_c_426_n N_A_311_413#_c_510_p
+ N_A_311_413#_c_409_n N_A_311_413#_c_461_n N_A_311_413#_c_419_n
+ N_A_311_413#_c_410_n N_A_311_413#_c_420_n N_A_311_413#_c_411_n
+ N_A_311_413#_c_412_n N_A_311_413#_c_413_n N_A_311_413#_c_414_n
+ PM_SKY130_FD_SC_HD__OR4BB_1%A_311_413#
x_PM_SKY130_FD_SC_HD__OR4BB_1%VPWR N_VPWR_M1011_d N_VPWR_M1012_d N_VPWR_c_522_n
+ N_VPWR_c_523_n VPWR N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n
+ N_VPWR_c_521_n N_VPWR_c_528_n N_VPWR_c_529_n PM_SKY130_FD_SC_HD__OR4BB_1%VPWR
x_PM_SKY130_FD_SC_HD__OR4BB_1%X N_X_M1000_d N_X_M1002_d N_X_c_581_n N_X_c_583_n
+ N_X_c_582_n X PM_SKY130_FD_SC_HD__OR4BB_1%X
x_PM_SKY130_FD_SC_HD__OR4BB_1%VGND N_VGND_M1008_d N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_M1010_d N_VGND_c_599_n N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n
+ VGND N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n N_VGND_c_606_n
+ N_VGND_c_607_n N_VGND_c_608_n N_VGND_c_609_n N_VGND_c_610_n N_VGND_c_611_n
+ PM_SKY130_FD_SC_HD__OR4BB_1%VGND
cc_1 VNB N_C_N_c_93_n 0.023245f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_2 VNB N_C_N_c_94_n 0.00602296f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_C_N_c_95_n 0.0208027f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_4 VNB D_N 0.00232937f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_5 VNB N_D_N_c_126_n 0.0266058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_D_N_c_127_n 0.0188611f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_7 VNB N_A_205_93#_M1003_g 0.0322926f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_8 VNB N_A_205_93#_c_163_n 0.00443081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_205_93#_c_164_n 6.63735e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_205_93#_c_165_n 0.0125002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_205_93#_c_166_n 0.00163498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_205_93#_c_167_n 0.0339165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_M1006_g 0.0266413f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_14 VNB N_A_27_410#_c_234_n 0.0222773f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.325
cc_15 VNB N_A_27_410#_c_235_n 2.24825e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_410#_c_236_n 0.0221852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_237_n 0.0186165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_M1001_g 0.0157284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_c_323_n 0.0147133f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_20 VNB N_B_c_324_n 0.00821622f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_21 VNB N_A_M1010_g 0.0277171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.26
cc_22 VNB N_A_c_366_n 0.0200358f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_23 VNB N_A_c_367_n 0.00432763f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_24 VNB N_A_311_413#_c_407_n 0.0113346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_311_413#_c_408_n 0.00438927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_311_413#_c_409_n 0.00233469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_311_413#_c_410_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_311_413#_c_411_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_311_413#_c_412_n 0.0234012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_311_413#_c_413_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_311_413#_c_414_n 0.0193297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_521_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_581_n 0.0137601f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_34 VNB N_X_c_582_n 0.0241563f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_35 VNB N_VGND_c_599_n 0.0126166f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_36 VNB N_VGND_c_600_n 0.00680485f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.53
cc_37 VNB N_VGND_c_601_n 3.0452e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_602_n 3.95722e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_603_n 0.0184121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_604_n 0.0123176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_605_n 0.0111699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_606_n 0.0166241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_607_n 0.238487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_608_n 0.0242387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_609_n 0.00593763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_610_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_611_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_C_N_M1011_g 0.0562995f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.26
cc_49 VPB N_C_N_c_93_n 0.00472379f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_50 VPB N_C_N_c_94_n 0.0023481f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_51 VPB N_D_N_M1013_g 0.0229391f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.675
cc_52 VPB D_N 5.14684e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_53 VPB N_D_N_c_126_n 0.00586379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_205_93#_M1005_g 0.0635781f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_55 VPB N_A_205_93#_c_169_n 0.00837676f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_56 VPB N_A_205_93#_c_164_n 0.0040018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_205_93#_c_167_n 0.0104025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_410#_M1004_g 0.0190829f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_59 VPB N_A_27_410#_c_234_n 0.026212f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.325
cc_60 VPB N_A_27_410#_c_240_n 0.016454f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.19
cc_61 VPB N_A_27_410#_c_241_n 0.0198572f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.53
cc_62 VPB N_A_27_410#_c_242_n 0.00680513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_410#_c_243_n 0.00589342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_410#_c_244_n 0.00201079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_410#_c_235_n 9.16196e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_410#_c_236_n 0.00435359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_410#_c_247_n 0.0113037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_B_M1001_g 0.0267766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB B 0.0122602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B_c_327_n 0.0353878f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_71 VPB N_A_M1012_g 0.0209374f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=0.675
cc_72 VPB N_A_c_366_n 0.00399502f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_73 VPB N_A_c_367_n 0.0033301f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_74 VPB N_A_311_413#_M1002_g 0.0244726f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_75 VPB N_A_311_413#_c_416_n 0.00575913f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_76 VPB N_A_311_413#_c_417_n 0.00241773f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_311_413#_c_418_n 0.003558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_311_413#_c_419_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_311_413#_c_420_n 0.00130727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_311_413#_c_412_n 0.00544454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_522_n 0.0106806f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_82 VPB N_VPWR_c_523_n 0.0108954f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_83 VPB N_VPWR_c_524_n 0.0145108f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_84 VPB N_VPWR_c_525_n 0.0633094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_526_n 0.0177135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_521_n 0.0671796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_528_n 0.00519112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_529_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_X_c_583_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_90 VPB N_X_c_582_n 0.00880472f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_91 VPB X 0.032187f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.325
cc_92 N_C_N_M1011_g N_D_N_M1013_g 0.0243394f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_93 N_C_N_c_94_n N_D_N_M1013_g 0.00410692f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_94 N_C_N_c_93_n D_N 2.85663e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_95 N_C_N_c_94_n D_N 0.0259635f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C_N_c_93_n N_D_N_c_126_n 0.019221f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_97 N_C_N_c_94_n N_D_N_c_126_n 0.00225922f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_98 N_C_N_c_95_n N_D_N_c_127_n 0.0104665f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_99 N_C_N_c_94_n N_A_205_93#_c_169_n 0.0114587f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_N_c_94_n N_A_205_93#_c_164_n 0.00627776f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_101 N_C_N_M1011_g N_A_27_410#_c_234_n 0.0132977f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_102 N_C_N_c_93_n N_A_27_410#_c_234_n 0.00753248f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_103 N_C_N_c_94_n N_A_27_410#_c_234_n 0.0528067f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_104 N_C_N_c_95_n N_A_27_410#_c_234_n 0.0052679f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C_N_M1011_g N_A_27_410#_c_240_n 0.00143901f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_106 N_C_N_M1011_g N_A_27_410#_c_241_n 0.0143338f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_107 N_C_N_c_93_n N_A_27_410#_c_241_n 8.32653e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_108 N_C_N_c_94_n N_A_27_410#_c_241_n 0.0279958f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_109 N_C_N_c_95_n N_A_27_410#_c_237_n 3.39179e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_110 N_C_N_c_94_n N_VPWR_M1011_d 0.00432228f $X=0.51 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_111 N_C_N_M1011_g N_VPWR_c_522_n 0.0100087f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_112 N_C_N_M1011_g N_VPWR_c_524_n 0.00334979f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_113 N_C_N_M1011_g N_VPWR_c_521_n 0.0048928f $X=0.47 $Y=2.26 $X2=0 $Y2=0
cc_114 N_C_N_c_94_n N_VGND_c_599_n 0.0108718f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_N_c_95_n N_VGND_c_599_n 0.00422719f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C_N_c_95_n N_VGND_c_607_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_N_c_95_n N_VGND_c_608_n 0.00510437f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_118 N_D_N_M1013_g N_A_205_93#_c_169_n 0.00312367f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_119 D_N N_A_205_93#_c_169_n 0.0141649f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_120 N_D_N_c_126_n N_A_205_93#_c_169_n 0.00349053f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_121 D_N N_A_205_93#_c_163_n 0.00622755f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_122 N_D_N_c_126_n N_A_205_93#_c_163_n 2.31143e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_123 N_D_N_c_127_n N_A_205_93#_c_163_n 0.00422498f $X=1.03 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_D_N_M1013_g N_A_205_93#_c_164_n 0.00310263f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_125 D_N N_A_205_93#_c_164_n 0.00622755f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_126 N_D_N_c_126_n N_A_205_93#_c_164_n 2.31143e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_127 D_N N_A_205_93#_c_165_n 0.012483f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_128 N_D_N_c_126_n N_A_205_93#_c_165_n 0.00272654f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_129 N_D_N_c_127_n N_A_205_93#_c_165_n 3.44947e-19 $X=1.03 $Y=0.995 $X2=0
+ $Y2=0
cc_130 D_N N_A_205_93#_c_166_n 0.014254f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_131 N_D_N_c_126_n N_A_205_93#_c_166_n 5.70522e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_132 D_N N_A_205_93#_c_167_n 8.91535e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_133 N_D_N_c_126_n N_A_205_93#_c_167_n 0.012914f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_134 N_D_N_M1013_g N_A_27_410#_c_241_n 0.0154775f $X=0.955 $Y=1.695 $X2=0
+ $Y2=0
cc_135 D_N N_A_27_410#_c_241_n 0.00124584f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_136 N_D_N_M1013_g N_VPWR_c_525_n 0.00259183f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_137 N_D_N_M1013_g N_VPWR_c_521_n 0.00417489f $X=0.955 $Y=1.695 $X2=0 $Y2=0
cc_138 N_D_N_c_127_n N_VGND_c_599_n 0.00163f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_139 N_D_N_c_127_n N_VGND_c_600_n 0.00211678f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_140 N_D_N_c_127_n N_VGND_c_603_n 0.00510437f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_141 N_D_N_c_127_n N_VGND_c_607_n 0.00512902f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_205_93#_M1003_g N_A_27_410#_M1006_g 0.0226254f $X=1.89 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_205_93#_M1005_g N_A_27_410#_M1004_g 0.0243913f $X=1.89 $Y=2.275 $X2=0
+ $Y2=0
cc_144 N_A_205_93#_M1013_d N_A_27_410#_c_241_n 0.00247661f $X=1.03 $Y=1.485
+ $X2=0 $Y2=0
cc_145 N_A_205_93#_M1005_g N_A_27_410#_c_241_n 0.00812129f $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_146 N_A_205_93#_c_169_n N_A_27_410#_c_241_n 0.0398304f $X=1.405 $Y=1.61 $X2=0
+ $Y2=0
cc_147 N_A_205_93#_c_166_n N_A_27_410#_c_241_n 0.0045774f $X=1.645 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_A_205_93#_c_167_n N_A_27_410#_c_241_n 0.00315934f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_205_93#_M1005_g N_A_27_410#_c_242_n 0.010188f $X=1.89 $Y=2.275 $X2=0
+ $Y2=0
cc_150 N_A_205_93#_c_169_n N_A_27_410#_c_242_n 0.00913778f $X=1.405 $Y=1.61
+ $X2=0 $Y2=0
cc_151 N_A_205_93#_M1005_g N_A_27_410#_c_243_n 0.0065405f $X=1.89 $Y=2.275 $X2=0
+ $Y2=0
cc_152 N_A_205_93#_M1005_g N_A_27_410#_c_244_n 0.00882292f $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_153 N_A_205_93#_c_169_n N_A_27_410#_c_244_n 0.00554032f $X=1.405 $Y=1.61
+ $X2=0 $Y2=0
cc_154 N_A_205_93#_c_164_n N_A_27_410#_c_244_n 0.00921709f $X=1.49 $Y=1.525
+ $X2=0 $Y2=0
cc_155 N_A_205_93#_c_166_n N_A_27_410#_c_244_n 0.00673601f $X=1.645 $Y=1.16
+ $X2=0 $Y2=0
cc_156 N_A_205_93#_c_167_n N_A_27_410#_c_244_n 0.00178889f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_205_93#_M1005_g N_A_27_410#_c_235_n 8.16443e-19 $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_158 N_A_205_93#_c_163_n N_A_27_410#_c_235_n 0.00177015f $X=1.49 $Y=1.075
+ $X2=0 $Y2=0
cc_159 N_A_205_93#_c_164_n N_A_27_410#_c_235_n 0.00438503f $X=1.49 $Y=1.525
+ $X2=0 $Y2=0
cc_160 N_A_205_93#_c_166_n N_A_27_410#_c_235_n 0.006225f $X=1.645 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_205_93#_c_167_n N_A_27_410#_c_235_n 0.00131394f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_205_93#_c_166_n N_A_27_410#_c_236_n 4.75093e-19 $X=1.645 $Y=1.16
+ $X2=0 $Y2=0
cc_163 N_A_205_93#_c_167_n N_A_27_410#_c_236_n 0.0213915f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_205_93#_M1005_g N_B_M1001_g 0.00153736f $X=1.89 $Y=2.275 $X2=0 $Y2=0
cc_165 N_A_205_93#_M1005_g B 0.00223393f $X=1.89 $Y=2.275 $X2=0 $Y2=0
cc_166 N_A_205_93#_M1005_g N_B_c_327_n 0.00325164f $X=1.89 $Y=2.275 $X2=0 $Y2=0
cc_167 N_A_205_93#_M1005_g N_A_311_413#_c_416_n 0.00971256f $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_168 N_A_205_93#_M1005_g N_A_311_413#_c_417_n 0.00494253f $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_169 N_A_205_93#_M1003_g N_A_311_413#_c_408_n 0.00224864f $X=1.89 $Y=0.445
+ $X2=0 $Y2=0
cc_170 N_A_205_93#_c_165_n N_A_311_413#_c_408_n 0.00795991f $X=1.16 $Y=0.66
+ $X2=0 $Y2=0
cc_171 N_A_205_93#_M1005_g N_A_311_413#_c_426_n 0.00129708f $X=1.89 $Y=2.275
+ $X2=0 $Y2=0
cc_172 N_A_205_93#_M1005_g N_VPWR_c_525_n 0.00375986f $X=1.89 $Y=2.275 $X2=0
+ $Y2=0
cc_173 N_A_205_93#_M1005_g N_VPWR_c_521_n 0.00798404f $X=1.89 $Y=2.275 $X2=0
+ $Y2=0
cc_174 N_A_205_93#_c_165_n N_VGND_M1003_s 2.00035e-19 $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_175 N_A_205_93#_c_165_n N_VGND_c_599_n 8.07382e-19 $X=1.16 $Y=0.66 $X2=0
+ $Y2=0
cc_176 N_A_205_93#_M1003_g N_VGND_c_600_n 0.00915659f $X=1.89 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_205_93#_c_165_n N_VGND_c_600_n 0.0110792f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_178 N_A_205_93#_c_166_n N_VGND_c_600_n 0.0064624f $X=1.645 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_205_93#_c_167_n N_VGND_c_600_n 0.00452715f $X=1.89 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A_205_93#_M1003_g N_VGND_c_601_n 6.24108e-19 $X=1.89 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_205_93#_c_165_n N_VGND_c_603_n 0.0091771f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_182 N_A_205_93#_M1003_g N_VGND_c_604_n 0.0046653f $X=1.89 $Y=0.445 $X2=0
+ $Y2=0
cc_183 N_A_205_93#_M1003_g N_VGND_c_607_n 0.00803392f $X=1.89 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_A_205_93#_c_165_n N_VGND_c_607_n 0.0125849f $X=1.16 $Y=0.66 $X2=0 $Y2=0
cc_185 N_A_27_410#_c_243_n N_B_M1001_g 7.72856e-19 $X=2.225 $Y=1.5 $X2=0 $Y2=0
cc_186 N_A_27_410#_c_235_n N_B_M1001_g 8.95596e-19 $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_410#_c_236_n N_B_M1001_g 0.0641534f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_27_410#_M1006_g N_B_c_323_n 0.0136823f $X=2.325 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_27_410#_M1006_g N_B_c_324_n 0.0126742f $X=2.325 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_235_n N_A_c_367_n 0.0217601f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_27_410#_c_236_n N_A_c_367_n 0.00220685f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_410#_c_241_n N_A_311_413#_c_416_n 0.0272384f $X=1.745 $Y=1.95
+ $X2=0 $Y2=0
cc_193 N_A_27_410#_c_243_n N_A_311_413#_c_416_n 0.00376842f $X=2.225 $Y=1.5
+ $X2=0 $Y2=0
cc_194 N_A_27_410#_M1004_g N_A_311_413#_c_417_n 0.00197943f $X=2.37 $Y=1.695
+ $X2=0 $Y2=0
cc_195 N_A_27_410#_c_241_n N_A_311_413#_c_417_n 0.00625142f $X=1.745 $Y=1.95
+ $X2=0 $Y2=0
cc_196 N_A_27_410#_M1006_g N_A_311_413#_c_407_n 0.0112518f $X=2.325 $Y=0.445
+ $X2=0 $Y2=0
cc_197 N_A_27_410#_c_243_n N_A_311_413#_c_407_n 0.0012205f $X=2.225 $Y=1.5 $X2=0
+ $Y2=0
cc_198 N_A_27_410#_c_235_n N_A_311_413#_c_407_n 0.012736f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_27_410#_c_236_n N_A_311_413#_c_407_n 0.00313532f $X=2.31 $Y=1.16
+ $X2=0 $Y2=0
cc_200 N_A_27_410#_c_243_n N_A_311_413#_c_408_n 0.00589573f $X=2.225 $Y=1.5
+ $X2=0 $Y2=0
cc_201 N_A_27_410#_c_236_n N_A_311_413#_c_408_n 2.86694e-19 $X=2.31 $Y=1.16
+ $X2=0 $Y2=0
cc_202 N_A_27_410#_M1004_g N_A_311_413#_c_418_n 0.0121016f $X=2.37 $Y=1.695
+ $X2=0 $Y2=0
cc_203 N_A_27_410#_c_243_n N_A_311_413#_c_418_n 0.00656826f $X=2.225 $Y=1.5
+ $X2=0 $Y2=0
cc_204 N_A_27_410#_c_241_n N_A_311_413#_c_426_n 0.00786633f $X=1.745 $Y=1.95
+ $X2=0 $Y2=0
cc_205 N_A_27_410#_c_242_n N_A_311_413#_c_426_n 0.00628038f $X=1.83 $Y=1.865
+ $X2=0 $Y2=0
cc_206 N_A_27_410#_c_243_n N_A_311_413#_c_426_n 0.0109594f $X=2.225 $Y=1.5 $X2=0
+ $Y2=0
cc_207 N_A_27_410#_c_236_n N_A_311_413#_c_426_n 2.10144e-19 $X=2.31 $Y=1.16
+ $X2=0 $Y2=0
cc_208 N_A_27_410#_c_243_n N_A_311_413#_c_420_n 0.00276731f $X=2.225 $Y=1.5
+ $X2=0 $Y2=0
cc_209 N_A_27_410#_c_241_n N_VPWR_M1011_d 0.00538813f $X=1.745 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_210 N_A_27_410#_c_241_n N_VPWR_c_522_n 0.0229102f $X=1.745 $Y=1.95 $X2=0
+ $Y2=0
cc_211 N_A_27_410#_c_240_n N_VPWR_c_524_n 0.0168632f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_212 N_A_27_410#_c_241_n N_VPWR_c_524_n 0.00256078f $X=1.745 $Y=1.95 $X2=0
+ $Y2=0
cc_213 N_A_27_410#_M1004_g N_VPWR_c_525_n 0.00327927f $X=2.37 $Y=1.695 $X2=0
+ $Y2=0
cc_214 N_A_27_410#_c_241_n N_VPWR_c_525_n 0.0106725f $X=1.745 $Y=1.95 $X2=0
+ $Y2=0
cc_215 N_A_27_410#_M1004_g N_VPWR_c_521_n 0.00417489f $X=2.37 $Y=1.695 $X2=0
+ $Y2=0
cc_216 N_A_27_410#_c_240_n N_VPWR_c_521_n 0.00987599f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_217 N_A_27_410#_c_241_n N_VPWR_c_521_n 0.0238029f $X=1.745 $Y=1.95 $X2=0
+ $Y2=0
cc_218 N_A_27_410#_c_243_n A_393_413# 0.00263772f $X=2.225 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_27_410#_c_237_n N_VGND_c_599_n 0.0104991f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_220 N_A_27_410#_M1006_g N_VGND_c_600_n 6.22445e-19 $X=2.325 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_27_410#_M1006_g N_VGND_c_601_n 0.00728835f $X=2.325 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_27_410#_M1006_g N_VGND_c_604_n 0.00341689f $X=2.325 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_27_410#_M1006_g N_VGND_c_607_n 0.00409245f $X=2.325 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_27_410#_c_237_n N_VGND_c_607_n 0.0105585f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_225 N_A_27_410#_c_237_n N_VGND_c_608_n 0.00957361f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_226 N_B_M1001_g N_A_M1010_g 0.00392288f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_227 N_B_c_323_n N_A_M1010_g 0.0207641f $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_228 N_B_M1001_g N_A_M1012_g 0.0299871f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_229 B N_A_M1012_g 8.99686e-19 $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_230 N_B_M1001_g N_A_c_366_n 0.0213087f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_231 N_B_M1001_g N_A_c_367_n 0.0141584f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_232 N_B_c_324_n N_A_c_367_n 4.43208e-19 $X=2.737 $Y=0.91 $X2=0 $Y2=0
cc_233 B N_A_311_413#_c_416_n 0.0130053f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_234 N_B_c_327_n N_A_311_413#_c_416_n 6.32819e-19 $X=2.79 $Y=2.335 $X2=0 $Y2=0
cc_235 N_B_M1001_g N_A_311_413#_c_417_n 0.00201096f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_236 B N_A_311_413#_c_417_n 0.00542028f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_237 N_B_c_323_n N_A_311_413#_c_407_n 0.00699162f $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_238 N_B_c_324_n N_A_311_413#_c_407_n 0.00481812f $X=2.737 $Y=0.91 $X2=0 $Y2=0
cc_239 N_B_M1001_g N_A_311_413#_c_418_n 0.0107156f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_240 B N_A_311_413#_c_418_n 0.0349748f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_241 N_B_c_327_n N_A_311_413#_c_418_n 0.00101546f $X=2.79 $Y=2.335 $X2=0 $Y2=0
cc_242 N_B_M1001_g N_A_311_413#_c_420_n 0.00538706f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_243 B N_A_311_413#_c_420_n 0.0138251f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_244 N_B_M1001_g N_VPWR_c_523_n 0.00280623f $X=2.73 $Y=1.695 $X2=0 $Y2=0
cc_245 B N_VPWR_c_523_n 0.0285382f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_246 N_B_c_327_n N_VPWR_c_523_n 0.00108286f $X=2.79 $Y=2.335 $X2=0 $Y2=0
cc_247 B N_VPWR_c_525_n 0.0396304f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_248 N_B_c_327_n N_VPWR_c_525_n 0.00774997f $X=2.79 $Y=2.335 $X2=0 $Y2=0
cc_249 B N_VPWR_c_521_n 0.0238619f $X=2.905 $Y=2.125 $X2=0 $Y2=0
cc_250 N_B_c_327_n N_VPWR_c_521_n 0.0109691f $X=2.79 $Y=2.335 $X2=0 $Y2=0
cc_251 N_B_c_323_n N_VGND_c_601_n 0.00716819f $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_252 N_B_c_323_n N_VGND_c_602_n 6.24658e-19 $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_253 N_B_c_323_n N_VGND_c_605_n 0.00341689f $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_254 N_B_c_323_n N_VGND_c_607_n 0.00405445f $X=2.737 $Y=0.76 $X2=0 $Y2=0
cc_255 N_A_M1012_g N_A_311_413#_M1002_g 0.0189405f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_256 N_A_c_367_n N_A_311_413#_c_407_n 0.0189424f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_c_367_n N_A_311_413#_c_418_n 0.0101811f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_M1010_g N_A_311_413#_c_409_n 0.011795f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_c_366_n N_A_311_413#_c_409_n 0.00220162f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A_c_367_n N_A_311_413#_c_409_n 0.0166868f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_M1012_g N_A_311_413#_c_461_n 0.0112137f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_262 N_A_c_367_n N_A_311_413#_c_461_n 0.00969518f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_M1012_g N_A_311_413#_c_419_n 0.0034529f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_264 N_A_c_366_n N_A_311_413#_c_410_n 5.77159e-19 $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_c_367_n N_A_311_413#_c_410_n 0.0146254f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_M1012_g N_A_311_413#_c_420_n 0.00964298f $X=3.165 $Y=1.695 $X2=0
+ $Y2=0
cc_267 N_A_c_366_n N_A_311_413#_c_420_n 0.00156816f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_c_367_n N_A_311_413#_c_420_n 0.0112207f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_c_366_n N_A_311_413#_c_411_n 0.00186332f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_c_367_n N_A_311_413#_c_411_n 0.027072f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_c_366_n N_A_311_413#_c_412_n 0.0202671f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_c_367_n N_A_311_413#_c_412_n 3.56347e-19 $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_M1010_g N_A_311_413#_c_413_n 0.0034529f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_274 N_A_M1010_g N_A_311_413#_c_414_n 0.0177679f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_M1012_g N_VPWR_c_523_n 0.00293484f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_276 N_A_M1012_g N_VPWR_c_525_n 0.00264181f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_277 N_A_M1012_g N_VPWR_c_521_n 0.00333991f $X=3.165 $Y=1.695 $X2=0 $Y2=0
cc_278 N_A_M1010_g N_VGND_c_601_n 6.21849e-19 $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_279 N_A_M1010_g N_VGND_c_602_n 0.00746702f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_M1010_g N_VGND_c_605_n 0.00341689f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_281 N_A_M1010_g N_VGND_c_607_n 0.00405445f $X=3.165 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_311_413#_c_461_n N_VPWR_M1012_d 0.00526233f $X=3.44 $Y=1.58 $X2=0
+ $Y2=0
cc_283 N_A_311_413#_c_416_n N_VPWR_c_522_n 0.0057161f $X=2.085 $Y=2.29 $X2=0
+ $Y2=0
cc_284 N_A_311_413#_M1002_g N_VPWR_c_523_n 0.00485906f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_285 N_A_311_413#_c_461_n N_VPWR_c_523_n 0.0190361f $X=3.44 $Y=1.58 $X2=0
+ $Y2=0
cc_286 N_A_311_413#_c_420_n N_VPWR_c_523_n 0.00605542f $X=3.035 $Y=1.58 $X2=0
+ $Y2=0
cc_287 N_A_311_413#_c_412_n N_VPWR_c_523_n 2.11345e-19 $X=3.63 $Y=1.16 $X2=0
+ $Y2=0
cc_288 N_A_311_413#_c_416_n N_VPWR_c_525_n 0.0285048f $X=2.085 $Y=2.29 $X2=0
+ $Y2=0
cc_289 N_A_311_413#_M1002_g N_VPWR_c_526_n 0.00585385f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_311_413#_M1005_s N_VPWR_c_521_n 0.00217968f $X=1.555 $Y=2.065 $X2=0
+ $Y2=0
cc_291 N_A_311_413#_M1002_g N_VPWR_c_521_n 0.0128443f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_292 N_A_311_413#_c_416_n N_VPWR_c_521_n 0.0256417f $X=2.085 $Y=2.29 $X2=0
+ $Y2=0
cc_293 N_A_311_413#_c_418_n N_VPWR_c_521_n 0.00841166f $X=2.95 $Y=1.87 $X2=0
+ $Y2=0
cc_294 N_A_311_413#_c_416_n A_393_413# 0.0042428f $X=2.085 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_295 N_A_311_413#_c_417_n A_393_413# 0.00292122f $X=2.17 $Y=2.205 $X2=-0.19
+ $Y2=-0.24
cc_296 N_A_311_413#_c_426_n A_393_413# 0.00335245f $X=2.255 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_297 N_A_311_413#_c_418_n A_489_297# 0.00366293f $X=2.95 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_298 N_A_311_413#_c_418_n A_561_297# 0.00180544f $X=2.95 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_311_413#_c_420_n A_561_297# 0.00465932f $X=3.035 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_311_413#_M1002_g N_X_c_582_n 0.00349311f $X=3.655 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A_311_413#_c_409_n N_X_c_582_n 0.0035218f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_311_413#_c_419_n N_X_c_582_n 0.00841221f $X=3.525 $Y=1.495 $X2=0
+ $Y2=0
cc_303 N_A_311_413#_c_411_n N_X_c_582_n 0.024459f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_304 N_A_311_413#_c_412_n N_X_c_582_n 0.00753248f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_311_413#_c_413_n N_X_c_582_n 0.00836618f $X=3.577 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_311_413#_c_414_n N_X_c_582_n 0.00441003f $X=3.63 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_311_413#_c_409_n N_VGND_M1010_d 0.00464421f $X=3.44 $Y=0.74 $X2=0
+ $Y2=0
cc_308 N_A_311_413#_c_413_n N_VGND_M1010_d 6.98847e-19 $X=3.577 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_311_413#_c_502_p N_VGND_c_601_n 0.0124499f $X=2.1 $Y=0.47 $X2=0 $Y2=0
cc_310 N_A_311_413#_c_407_n N_VGND_c_601_n 0.020154f $X=2.87 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A_311_413#_c_409_n N_VGND_c_602_n 0.022675f $X=3.44 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_311_413#_c_412_n N_VGND_c_602_n 2.33671e-19 $X=3.63 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_311_413#_c_414_n N_VGND_c_602_n 0.0130203f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_311_413#_c_502_p N_VGND_c_604_n 0.00861358f $X=2.1 $Y=0.47 $X2=0
+ $Y2=0
cc_315 N_A_311_413#_c_407_n N_VGND_c_604_n 0.00299685f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_311_413#_c_407_n N_VGND_c_605_n 0.00273399f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_311_413#_c_510_p N_VGND_c_605_n 0.00846569f $X=2.955 $Y=0.47 $X2=0
+ $Y2=0
cc_318 N_A_311_413#_c_409_n N_VGND_c_605_n 0.00273399f $X=3.44 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_311_413#_c_409_n N_VGND_c_606_n 3.34073e-19 $X=3.44 $Y=0.74 $X2=0
+ $Y2=0
cc_320 N_A_311_413#_c_414_n N_VGND_c_606_n 0.00524631f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_321 N_A_311_413#_M1003_d N_VGND_c_607_n 0.0043277f $X=1.965 $Y=0.235 $X2=0
+ $Y2=0
cc_322 N_A_311_413#_M1007_d N_VGND_c_607_n 0.00256656f $X=2.82 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_311_413#_c_502_p N_VGND_c_607_n 0.00625722f $X=2.1 $Y=0.47 $X2=0
+ $Y2=0
cc_324 N_A_311_413#_c_407_n N_VGND_c_607_n 0.0101439f $X=2.87 $Y=0.74 $X2=0
+ $Y2=0
cc_325 N_A_311_413#_c_510_p N_VGND_c_607_n 0.00625722f $X=2.955 $Y=0.47 $X2=0
+ $Y2=0
cc_326 N_A_311_413#_c_409_n N_VGND_c_607_n 0.00638906f $X=3.44 $Y=0.74 $X2=0
+ $Y2=0
cc_327 N_A_311_413#_c_414_n N_VGND_c_607_n 0.00951738f $X=3.63 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_521_n A_393_413# 0.00214454f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_329 N_VPWR_c_521_n N_X_M1002_d 0.00399469f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_330 N_VPWR_c_526_n X 0.0190559f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_331 N_VPWR_c_521_n X 0.0105137f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_332 N_X_c_581_n N_VGND_c_606_n 0.00892672f $X=3.97 $Y=0.587 $X2=0 $Y2=0
cc_333 N_X_M1000_d N_VGND_c_607_n 0.00416042f $X=3.73 $Y=0.235 $X2=0 $Y2=0
cc_334 N_X_c_581_n N_VGND_c_607_n 0.00941771f $X=3.97 $Y=0.587 $X2=0 $Y2=0

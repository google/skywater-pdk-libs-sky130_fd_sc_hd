* NGSPICE file created from sky130_fd_sc_hd__a21bo_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_603_297# a_42_47# a_205_21# VPB phighvt w=1e+06u l=150000u
+  ad=1.06e+12p pd=1.012e+07u as=2.7e+11p ps=2.54e+06u
M1001 VPWR A1 a_603_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.38e+12p pd=1.276e+07u as=0p ps=0u
M1002 a_205_21# A1 a_861_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=1.495e+11p ps=1.76e+06u
M1003 a_205_21# a_42_47# a_603_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_861_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.261e+12p ps=1.038e+07u
M1005 VGND a_205_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.64e+11p ps=3.72e+06u
M1006 X a_205_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1007 X a_205_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_205_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_205_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_205_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_603_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1021_47# A1 a_205_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1013 VGND A2 a_1021_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_205_21# a_42_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_603_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_603_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR B1_N a_42_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1018 VPWR a_205_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_205_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_42_47# a_205_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND B1_N a_42_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.5025e+11p ps=2.07e+06u
.ends


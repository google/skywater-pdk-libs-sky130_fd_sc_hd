* File: sky130_fd_sc_hd__o21ba_4.spice.pex
* Created: Thu Aug 27 14:36:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BA_4%B1_N 1 3 6 8 9 13 15
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r42 9 15 10.0839 $w=2.78e-07 $l=2.45e-07 $layer=LI1_cond $X=0.745 $Y=1.53
+ $X2=0.745 $Y2=1.285
r43 8 15 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=0.69 $Y=1.18
+ $X2=0.745 $Y2=1.18
r44 8 14 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=1.18 $X2=0.59
+ $Y2=1.18
r45 4 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.325
+ $X2=0.59 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.59 $Y=1.325 $X2=0.59
+ $Y2=1.985
r47 1 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=0.995
+ $X2=0.59 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.59 $Y=0.995 $X2=0.59
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A_187_21# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 44 46 49 52 53 55 57 60 63 64 66 74
c162 74 0 1.22952e-19 $X=2.27 $Y=1.16
c163 64 0 7.57448e-20 $X=3.49 $Y=0.77
c164 46 0 1.12295e-19 $X=2.565 $Y=0.81
r165 71 72 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.85 $Y2=1.16
r166 69 71 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.01 $Y=1.16
+ $X2=1.43 $Y2=1.16
r167 62 64 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=3.42 $Y=0.77 $X2=3.49
+ $Y2=0.77
r168 62 63 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=3.42 $Y=0.77
+ $X2=3.235 $Y2=0.77
r169 55 68 3.19664 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=4.257 $Y=1.795
+ $X2=4.257 $Y2=1.96
r170 55 57 8.23174 $w=2.43e-07 $l=1.75e-07 $layer=LI1_cond $X=4.257 $Y=1.795
+ $X2=4.257 $Y2=1.62
r171 54 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.585 $Y=1.88
+ $X2=3.49 $Y2=1.88
r172 53 68 3.91346 $w=1.7e-07 $l=1.56984e-07 $layer=LI1_cond $X=4.135 $Y=1.88
+ $X2=4.257 $Y2=1.96
r173 53 54 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.135 $Y=1.88
+ $X2=3.585 $Y2=1.88
r174 52 66 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=1.795
+ $X2=3.49 $Y2=1.88
r175 51 64 2.34666 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.49 $Y=0.895
+ $X2=3.49 $Y2=0.77
r176 51 52 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=3.49 $Y=0.895
+ $X2=3.49 $Y2=1.795
r177 50 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=1.88
+ $X2=2.9 $Y2=1.88
r178 49 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.395 $Y=1.88
+ $X2=3.49 $Y2=1.88
r179 49 50 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.395 $Y=1.88
+ $X2=2.985 $Y2=1.88
r180 46 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.565 $Y=0.81
+ $X2=3.235 $Y2=0.81
r181 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.48 $Y=0.895
+ $X2=2.565 $Y2=0.81
r182 43 44 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.48 $Y=0.895
+ $X2=2.48 $Y2=1.075
r183 41 74 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.14 $Y=1.16
+ $X2=2.27 $Y2=1.16
r184 41 72 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.14 $Y=1.16
+ $X2=1.85 $Y2=1.16
r185 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.16 $X2=2.14 $Y2=1.16
r186 38 44 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.395 $Y=1.175
+ $X2=2.48 $Y2=1.075
r187 38 40 14.1409 $w=1.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.395 $Y=1.175
+ $X2=2.14 $Y2=1.175
r188 34 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.325
+ $X2=2.27 $Y2=1.16
r189 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.27 $Y=1.325
+ $X2=2.27 $Y2=1.985
r190 31 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=1.16
r191 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.27 $Y=0.995
+ $X2=2.27 $Y2=0.56
r192 27 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.325
+ $X2=1.85 $Y2=1.16
r193 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.85 $Y=1.325
+ $X2=1.85 $Y2=1.985
r194 24 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=0.995
+ $X2=1.85 $Y2=1.16
r195 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.85 $Y=0.995
+ $X2=1.85 $Y2=0.56
r196 20 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.16
r197 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.43 $Y=1.325
+ $X2=1.43 $Y2=1.985
r198 17 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.16
r199 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r200 13 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.325
+ $X2=1.01 $Y2=1.16
r201 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.01 $Y=1.325
+ $X2=1.01 $Y2=1.985
r202 10 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.16
r203 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r204 3 68 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=1.485 $X2=4.26 $Y2=1.96
r205 3 57 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.125
+ $Y=1.485 $X2=4.26 $Y2=1.62
r206 2 60 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=1.96
r207 1 62 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A_27_297# 1 2 9 13 15 17 18 20 24 27 29 32
+ 34 36 40 41 43 46 51 59
c110 51 0 1.22952e-19 $X=2.97 $Y=1.16
c111 18 0 1.80164e-19 $X=3.63 $Y=0.995
c112 9 0 1.55753e-19 $X=2.69 $Y=1.985
r113 58 59 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.21 $Y=1.16
+ $X2=3.63 $Y2=1.16
r114 57 58 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.11 $Y=1.16 $X2=3.21
+ $Y2=1.16
r115 52 57 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.97 $Y=1.16
+ $X2=3.11 $Y2=1.16
r116 52 54 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.97 $Y=1.16
+ $X2=2.69 $Y2=1.16
r117 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=1.16 $X2=2.97 $Y2=1.16
r118 48 51 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.82 $Y=1.16
+ $X2=2.97 $Y2=1.16
r119 44 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.48 $Y=1.53
+ $X2=2.82 $Y2=1.53
r120 40 41 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.62
+ $X2=0.26 $Y2=1.455
r121 38 41 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.17 $Y=0.855
+ $X2=0.17 $Y2=1.455
r122 36 38 17.0806 $w=4.58e-07 $l=4.65e-07 $layer=LI1_cond $X=0.315 $Y=0.39
+ $X2=0.315 $Y2=0.855
r123 34 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=1.445
+ $X2=2.82 $Y2=1.53
r124 33 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=1.245
+ $X2=2.82 $Y2=1.16
r125 33 34 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.82 $Y=1.245
+ $X2=2.82 $Y2=1.445
r126 31 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=1.615
+ $X2=2.48 $Y2=1.53
r127 31 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.48 $Y=1.615
+ $X2=2.48 $Y2=1.875
r128 30 43 4.03347 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=1.96
+ $X2=0.26 $Y2=1.96
r129 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=1.96
+ $X2=2.48 $Y2=1.875
r130 29 30 127.872 $w=1.68e-07 $l=1.96e-06 $layer=LI1_cond $X=2.395 $Y=1.96
+ $X2=0.435 $Y2=1.96
r131 25 43 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=1.96
r132 25 27 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=2.3
r133 24 43 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.875
+ $X2=0.26 $Y2=1.96
r134 23 40 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=1.62
r135 23 24 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=1.875
r136 18 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.63 $Y=0.995
+ $X2=3.63 $Y2=1.16
r137 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.63 $Y=0.995
+ $X2=3.63 $Y2=0.56
r138 15 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=1.16
r139 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.995
+ $X2=3.21 $Y2=0.56
r140 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r141 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r142 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r143 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.985
r144 2 43 600 $w=1.7e-07 $l=5.72495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=1.96
r145 2 40 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=1.62
r146 2 27 600 $w=1.7e-07 $l=9.16215e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=2.3
r147 1 36 91 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.38 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A2 1 3 6 8 10 13 15 22
c54 22 0 1.24925e-19 $X=4.47 $Y=1.16
c55 1 0 7.57448e-20 $X=4.05 $Y=0.995
r56 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.26 $Y=1.16
+ $X2=4.47 $Y2=1.16
r57 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.26
+ $Y=1.16 $X2=4.26 $Y2=1.16
r58 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.05 $Y=1.16
+ $X2=4.26 $Y2=1.16
r59 15 21 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=4.37 $Y=1.175 $X2=4.26
+ $Y2=1.175
r60 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=1.325
+ $X2=4.47 $Y2=1.16
r61 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.47 $Y=1.325
+ $X2=4.47 $Y2=1.985
r62 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=1.16
r63 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=0.56
r64 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=1.325
+ $X2=4.05 $Y2=1.16
r65 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.05 $Y=1.325 $X2=4.05
+ $Y2=1.985
r66 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.05 $Y=0.995
+ $X2=4.05 $Y2=1.16
r67 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.05 $Y=0.995 $X2=4.05
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A1 1 3 6 8 10 13 15 22
c38 15 0 1.24925e-19 $X=5.29 $Y=1.19
r39 20 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.155 $Y=1.16
+ $X2=5.31 $Y2=1.16
r40 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.16 $X2=5.155 $Y2=1.16
r41 17 20 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=5.155 $Y2=1.16
r42 15 21 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=5.29 $Y=1.175
+ $X2=5.155 $Y2=1.175
r43 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.325
+ $X2=5.31 $Y2=1.16
r44 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.31 $Y=1.325
+ $X2=5.31 $Y2=1.985
r45 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=0.995
+ $X2=5.31 $Y2=1.16
r46 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.31 $Y=0.995
+ $X2=5.31 $Y2=0.56
r47 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.325
+ $X2=4.89 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.89 $Y=1.325 $X2=4.89
+ $Y2=1.985
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=0.995
+ $X2=4.89 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.89 $Y=0.995 $X2=4.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%VPWR 1 2 3 4 5 20 24 28 32 36 39 40 42 43 44
+ 46 51 67 68 71 74 77
r105 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r107 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r108 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 62 65 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r112 61 64 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r113 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r114 59 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r115 59 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r116 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r117 56 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.48 $Y2=2.72
r118 56 58 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.99 $Y2=2.72
r119 55 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 55 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r121 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r122 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.64 $Y2=2.72
r123 52 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.48 $Y2=2.72
r125 51 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 50 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r127 50 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 47 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=0.8 $Y2=2.72
r130 47 49 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.965 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.64 $Y2=2.72
r132 46 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 44 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 42 64 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=4.83 $Y2=2.72
r135 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=5.1 $Y2=2.72
r136 41 67 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=2.72
+ $X2=5.1 $Y2=2.72
r138 40 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 39 58 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.2 $Y=2.72
+ $X2=2.99 $Y2=2.72
r140 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.2 $Y=2.72
+ $X2=3.325 $Y2=2.72
r141 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=2.635 $X2=5.1
+ $Y2=2.72
r142 34 36 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.1 $Y=2.635
+ $X2=5.1 $Y2=2
r143 30 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=2.72
r144 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=2.3
r145 26 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=2.635
+ $X2=2.48 $Y2=2.72
r146 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.48 $Y=2.635
+ $X2=2.48 $Y2=2.3
r147 22 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=2.635
+ $X2=1.64 $Y2=2.72
r148 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=2.635
+ $X2=1.64 $Y2=2.3
r149 18 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.635 $X2=0.8
+ $Y2=2.72
r150 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.8 $Y=2.635
+ $X2=0.8 $Y2=2.3
r151 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.965
+ $Y=1.485 $X2=5.1 $Y2=2
r152 4 32 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=2.3
r153 3 28 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.485 $X2=2.48 $Y2=2.3
r154 2 24 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.485 $X2=1.64 $Y2=2.3
r155 1 20 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.485 $X2=0.8 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%X 1 2 3 4 15 18 19 23 25 29 32
c57 23 0 1.55753e-19 $X=2.06 $Y=1.62
r58 29 32 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.06 $Y=0.51 $X2=2.06
+ $Y2=0.39
r59 28 29 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.06 $Y=0.725
+ $X2=2.06 $Y2=0.51
r60 21 27 4.37767 $w=2.6e-07 $l=2e-07 $layer=LI1_cond $X=1.455 $Y=1.575
+ $X2=1.255 $Y2=1.575
r61 21 23 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=1.455 $Y=1.575
+ $X2=2.06 $Y2=1.575
r62 20 25 3.9756 $w=1.8e-07 $l=2e-07 $layer=LI1_cond $X=1.455 $Y=0.815 $X2=1.255
+ $Y2=0.815
r63 19 28 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.895 $Y=0.815
+ $X2=2.06 $Y2=0.725
r64 19 20 27.1111 $w=1.78e-07 $l=4.4e-07 $layer=LI1_cond $X=1.895 $Y=0.815
+ $X2=1.455 $Y2=0.815
r65 18 27 2.84549 $w=4e-07 $l=1.3e-07 $layer=LI1_cond $X=1.255 $Y=1.445
+ $X2=1.255 $Y2=1.575
r66 17 25 2.77445 $w=3.65e-07 $l=9e-08 $layer=LI1_cond $X=1.255 $Y=0.905
+ $X2=1.255 $Y2=0.815
r67 17 18 15.558 $w=3.98e-07 $l=5.4e-07 $layer=LI1_cond $X=1.255 $Y=0.905
+ $X2=1.255 $Y2=1.445
r68 13 25 2.77445 $w=3.65e-07 $l=1.06066e-07 $layer=LI1_cond $X=1.22 $Y=0.725
+ $X2=1.255 $Y2=0.815
r69 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.22 $Y=0.725
+ $X2=1.22 $Y2=0.39
r70 4 23 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.925
+ $Y=1.485 $X2=2.06 $Y2=1.62
r71 3 27 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.22 $Y2=1.62
r72 2 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.925
+ $Y=0.235 $X2=2.06 $Y2=0.39
r73 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A_743_297# 1 2 3 10 12 13 14 16 18 21
r37 16 29 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=5.572 $Y=1.665
+ $X2=5.572 $Y2=1.56
r38 16 18 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=5.572 $Y=1.665
+ $X2=5.572 $Y2=2.3
r39 15 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.56
+ $X2=4.68 $Y2=1.56
r40 14 29 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=5.435 $Y=1.56
+ $X2=5.572 $Y2=1.56
r41 14 15 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=5.435 $Y=1.56
+ $X2=4.765 $Y2=1.56
r42 13 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.68 $Y=2.295
+ $X2=4.68 $Y2=2.38
r43 12 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.68 $Y=1.665
+ $X2=4.68 $Y2=1.56
r44 12 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.68 $Y=1.665
+ $X2=4.68 $Y2=2.295
r45 11 21 2.75731 $w=1.7e-07 $l=1.54919e-07 $layer=LI1_cond $X=3.925 $Y=2.38
+ $X2=3.805 $Y2=2.3
r46 10 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=2.38
+ $X2=4.68 $Y2=2.38
r47 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.595 $Y=2.38
+ $X2=3.925 $Y2=2.38
r48 3 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.485 $X2=5.52 $Y2=1.62
r49 3 18 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.485 $X2=5.52 $Y2=2.3
r50 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.485 $X2=4.68 $Y2=2.3
r51 2 25 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.485 $X2=4.68 $Y2=1.62
r52 1 21 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.485 $X2=3.84 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%VGND 1 2 3 4 5 18 20 24 28 32 36 38 39 41 42
+ 44 45 46 52 65 66 69 72
r98 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r99 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r100 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r101 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r102 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r103 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r104 60 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=2.53 $Y2=0
r105 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r106 57 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.48
+ $Y2=0
r107 57 59 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=3.91 $Y2=0
r108 56 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r109 56 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r110 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r111 53 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.64
+ $Y2=0
r112 53 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=2.07
+ $Y2=0
r113 52 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.48
+ $Y2=0
r114 52 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.07 $Y2=0
r115 50 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r116 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r117 46 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r118 44 62 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=4.83 $Y2=0
r119 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.015 $Y=0 $X2=5.1
+ $Y2=0
r120 43 65 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.75
+ $Y2=0
r121 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.1
+ $Y2=0
r122 41 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=3.91 $Y2=0
r123 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.26
+ $Y2=0
r124 40 62 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.345 $Y=0
+ $X2=4.83 $Y2=0
r125 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=0 $X2=4.26
+ $Y2=0
r126 38 49 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.69
+ $Y2=0
r127 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.8
+ $Y2=0
r128 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=0.085 $X2=5.1
+ $Y2=0
r129 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.1 $Y=0.085
+ $X2=5.1 $Y2=0.39
r130 30 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0
r131 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0.39
r132 26 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r133 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.39
r134 22 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0
r135 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.64 $Y=0.085
+ $X2=1.64 $Y2=0.39
r136 21 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.8
+ $Y2=0
r137 20 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.64
+ $Y2=0
r138 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=0.885 $Y2=0
r139 16 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r140 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.8 $Y=0.085
+ $X2=0.8 $Y2=0.39
r141 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.1 $Y2=0.39
r142 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.125
+ $Y=0.235 $X2=4.26 $Y2=0.39
r143 3 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.48 $Y2=0.39
r144 2 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.64 $Y2=0.39
r145 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.665
+ $Y=0.235 $X2=0.8 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_4%A_575_47# 1 2 3 4 13 17 18 19 23 25 29 35
c60 18 0 1.80164e-19 $X=3.88 $Y=0.725
r61 27 29 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=5.532 $Y=0.725
+ $X2=5.532 $Y2=0.39
r62 26 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.845 $Y=0.815
+ $X2=4.68 $Y2=0.815
r63 25 27 7.81092 $w=1.8e-07 $l=2.17391e-07 $layer=LI1_cond $X=5.355 $Y=0.815
+ $X2=5.532 $Y2=0.725
r64 25 26 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.355 $Y=0.815
+ $X2=4.845 $Y2=0.815
r65 21 35 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.68 $Y=0.725 $X2=4.68
+ $Y2=0.815
r66 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.68 $Y=0.725
+ $X2=4.68 $Y2=0.39
r67 20 34 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.005 $Y=0.815
+ $X2=3.88 $Y2=0.815
r68 19 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.515 $Y=0.815
+ $X2=4.68 $Y2=0.815
r69 19 20 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.515 $Y=0.815
+ $X2=4.005 $Y2=0.815
r70 18 34 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=3.88 $Y=0.725 $X2=3.88
+ $Y2=0.815
r71 17 32 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=3.88 $Y=0.475
+ $X2=3.88 $Y2=0.365
r72 17 18 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=3.88 $Y=0.475
+ $X2=3.88 $Y2=0.725
r73 13 32 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=3.755 $Y=0.365
+ $X2=3.88 $Y2=0.365
r74 13 15 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=3.755 $Y=0.365
+ $X2=3 $Y2=0.365
r75 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.385
+ $Y=0.235 $X2=5.52 $Y2=0.39
r76 3 23 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.545
+ $Y=0.235 $X2=4.68 $Y2=0.39
r77 2 34 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.84 $Y2=0.73
r78 2 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.84 $Y2=0.39
r79 1 15 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.235 $X2=3 $Y2=0.39
.ends


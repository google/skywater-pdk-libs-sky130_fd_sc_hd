* File: sky130_fd_sc_hd__clkdlybuf4s15_2.spice
* Created: Tue Sep  1 19:00:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s15_2.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s15_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.101055 AS=0.1134 PD=0.851776 PS=1.38 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_228_47#_M1003_d N_A_27_47#_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.65 AD=0.26325 AS=0.156395 PD=2.11 PS=1.31822 NRD=25.836 NRS=18.456 M=1
+ R=4.33333 SA=75000.6 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_228_47#_M1009_g N_A_362_333#_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.218175 AS=0.169 PD=1.65234 PS=1.82 NRD=64.608 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_362_333#_M1006_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.140975 PD=0.7 PS=1.06766 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_X_M1006_d N_A_362_333#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.2058 PD=0.7 PS=1.82 NRD=0 NRS=64.284 M=1 R=2.8 SA=75001.5
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_27_47#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.220714 AS=0.27 PD=1.57692 PS=2.54 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1001 N_A_228_47#_M1001_d N_A_27_47#_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.82 AD=0.3116 AS=0.180986 PD=2.4 PS=1.29308 NRD=27.6194 NRS=20.4092 M=1
+ R=5.46667 SA=75000.8 SB=75000.3 A=0.123 P=1.94 MULT=1
MM1004 N_VPWR_M1004_d N_A_228_47#_M1004_g N_A_362_333#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.82 AD=0.282585 AS=0.2173 PD=1.54088 PS=2.17 NRD=84.0796 NRS=0 M=1
+ R=5.46667 SA=75000.2 SB=75001.7 A=0.123 P=1.94 MULT=1
MM1002 N_VPWR_M1004_d N_A_362_333#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.344615 AS=0.14 PD=1.87912 PS=1.28 NRD=15.7403 NRS=0 M=1 R=6.66667
+ SA=75000.9 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_362_333#_M1007_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.49 AS=0.14 PD=2.98 PS=1.28 NRD=44.3053 NRS=0 M=1 R=6.66667 SA=75001.3
+ SB=75000.4 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__clkdlybuf4s15_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdlclkp_2.spice.pex
* Created: Thu Aug 27 14:47:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%SCE 3 7 9 10 17
r27 14 17 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r28 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.16
+ $X2=0.212 $Y2=1.53
r29 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r30 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r31 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.165
r32 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%GATE 3 7 9 10 15 16
c42 16 0 2.81318e-20 $X=0.94 $Y=1.16
c43 15 0 9.56754e-20 $X=0.94 $Y=1.16
r44 15 18 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=1.325
r45 15 17 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=0.915 $Y2=0.995
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r47 9 10 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.047 $Y=1.53
+ $X2=1.047 $Y2=1.87
r48 9 16 8.21746 $w=4.63e-07 $l=2.85e-07 $layer=LI1_cond $X=1.025 $Y=1.445
+ $X2=1.025 $Y2=1.16
r49 7 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.995
r50 3 18 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.83 $Y=2.165
+ $X2=0.83 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_147# 1 2 9 13 17 21 24 25 28 29 30
+ 33 35 37 41 44 53 54 57 60 68 74
c180 68 0 1.23968e-19 $X=1.78 $Y=1.74
c181 57 0 3.38573e-20 $X=1.615 $Y=1.53
c182 44 0 2.81939e-19 $X=4.08 $Y=1.19
c183 41 0 2.00517e-19 $X=1.615 $Y=1.325
c184 24 0 3.18278e-20 $X=1.45 $Y=0.87
c185 9 0 2.35132e-20 $X=1.375 $Y=0.415
r186 68 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.74
+ $X2=1.78 $Y2=1.905
r187 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=1.74 $X2=1.78 $Y2=1.74
r188 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.375 $Y=1.53
+ $X2=4.375 $Y2=1.53
r189 57 69 5.52036 $w=4.53e-07 $l=2.1e-07 $layer=LI1_cond $X=1.637 $Y=1.53
+ $X2=1.637 $Y2=1.74
r190 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.53
r191 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.76 $Y=1.53
+ $X2=1.615 $Y2=1.53
r192 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.23 $Y=1.53
+ $X2=4.375 $Y2=1.53
r193 53 54 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=4.23 $Y=1.53
+ $X2=1.76 $Y2=1.53
r194 44 74 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.08 $Y=1.19
+ $X2=4.08 $Y2=1.325
r195 44 73 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.08 $Y=1.19
+ $X2=4.08 $Y2=1.055
r196 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.08
+ $Y=1.19 $X2=4.08 $Y2=1.19
r197 41 57 5.38892 $w=4.53e-07 $l=2.05e-07 $layer=LI1_cond $X=1.637 $Y=1.325
+ $X2=1.637 $Y2=1.53
r198 40 41 3.94479 $w=4.53e-07 $l=1.2e-07 $layer=LI1_cond $X=1.615 $Y=1.205
+ $X2=1.615 $Y2=1.325
r199 35 37 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.71 $Y=0.615
+ $X2=4.71 $Y2=0.465
r200 31 61 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.46 $Y=1.62
+ $X2=4.335 $Y2=1.62
r201 31 33 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=4.46 $Y=1.62
+ $X2=4.845 $Y2=1.62
r202 30 61 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.335 $Y=1.495
+ $X2=4.335 $Y2=1.62
r203 29 30 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=4.335 $Y=1.275
+ $X2=4.335 $Y2=1.495
r204 28 29 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.315 $Y=1.19
+ $X2=4.335 $Y2=1.19
r205 28 43 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=1.19
+ $X2=4.08 $Y2=1.19
r206 27 35 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.315 $Y=0.7
+ $X2=4.71 $Y2=0.7
r207 27 28 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=4.315 $Y=0.785
+ $X2=4.315 $Y2=1.105
r208 25 63 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=0.87
+ $X2=1.375 $Y2=0.87
r209 24 40 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0.87
+ $X2=1.535 $Y2=1.205
r210 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=0.87 $X2=1.45 $Y2=0.87
r211 21 74 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.085 $Y=1.835
+ $X2=4.085 $Y2=1.325
r212 17 73 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.05 $Y=0.445
+ $X2=4.05 $Y2=1.055
r213 13 71 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.84 $Y=2.275
+ $X2=1.84 $Y2=1.905
r214 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=0.735
+ $X2=1.375 $Y2=0.87
r215 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.375 $Y=0.735
+ $X2=1.375 $Y2=0.415
r216 2 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.515 $X2=4.845 $Y2=1.66
r217 1 37 182 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.68 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_257_243# 1 2 9 11 12 15 17 20 23 24 26
+ 28 29 35 36 39 40 41
c120 40 0 1.47482e-19 $X=1.96 $Y=0.87
c121 36 0 1.27753e-19 $X=3.915 $Y=0.85
c122 35 0 5.81425e-21 $X=3.915 $Y=0.85
c123 26 0 1.45744e-19 $X=3.875 $Y=1.66
c124 17 0 2.81318e-20 $X=1.9 $Y=1.215
c125 12 0 2.67301e-20 $X=1.435 $Y=1.29
c126 9 0 3.17216e-20 $X=1.36 $Y=2.275
r127 39 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.87
+ $X2=1.96 $Y2=1.035
r128 39 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.87
+ $X2=1.96 $Y2=0.705
r129 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=0.87 $X2=1.96 $Y2=0.87
r130 36 48 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.787 $Y=0.85
+ $X2=3.787 $Y2=0.935
r131 36 47 2.69788 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.787 $Y=0.85
+ $X2=3.787 $Y2=0.765
r132 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.915 $Y=0.85
+ $X2=3.915 $Y2=0.85
r133 31 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.075 $Y=0.85
+ $X2=2.075 $Y2=0.85
r134 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.22 $Y=0.85
+ $X2=2.075 $Y2=0.85
r135 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.77 $Y=0.85
+ $X2=3.915 $Y2=0.85
r136 28 29 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=3.77 $Y=0.85
+ $X2=2.22 $Y2=0.85
r137 24 26 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.745 $Y=1.66
+ $X2=3.875 $Y2=1.66
r138 23 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.575
+ $X2=3.745 $Y2=1.66
r139 23 48 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.66 $Y=1.575
+ $X2=3.66 $Y2=0.935
r140 20 47 9.87808 $w=3.48e-07 $l=3e-07 $layer=LI1_cond $X=3.75 $Y=0.465
+ $X2=3.75 $Y2=0.765
r141 17 42 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.9 $Y=1.215
+ $X2=1.9 $Y2=1.035
r142 15 41 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.9 $Y=0.415
+ $X2=1.9 $Y2=0.705
r143 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.9 $Y2=1.215
r144 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.435 $Y2=1.29
r145 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.36 $Y=1.365
+ $X2=1.435 $Y2=1.29
r146 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.36 $Y=1.365
+ $X2=1.36 $Y2=2.275
r147 2 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.75
+ $Y=1.515 $X2=3.875 $Y2=1.66
r148 1 20 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=3.715
+ $Y=0.235 $X2=3.84 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_465_315# 1 2 9 13 17 21 23 27 31 33 36
+ 39 41 42 46 55
c128 46 0 1.8014e-19 $X=5.485 $Y=1.52
c129 39 0 1.77265e-19 $X=2.46 $Y=1.74
c130 36 0 4.48552e-20 $X=5.335 $Y=1.915
c131 33 0 9.5488e-20 $X=5.18 $Y=2
c132 13 0 1.38699e-19 $X=2.51 $Y=0.445
r133 47 55 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.485 $Y=1.52
+ $X2=5.575 $Y2=1.52
r134 47 52 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=5.485 $Y=1.52
+ $X2=5.435 $Y2=1.52
r135 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=1.52 $X2=5.485 $Y2=1.52
r136 39 51 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.74
+ $X2=2.46 $Y2=1.905
r137 39 50 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.46 $Y=1.74
+ $X2=2.46 $Y2=1.575
r138 38 41 3.38343 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=1.74
+ $X2=2.545 $Y2=1.74
r139 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.74 $X2=2.46 $Y2=1.74
r140 35 46 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.335 $Y=1.52
+ $X2=5.485 $Y2=1.52
r141 35 36 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=5.335 $Y=1.605
+ $X2=5.335 $Y2=1.915
r142 34 42 3.05 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.405 $Y=2
+ $X2=3.295 $Y2=1.86
r143 33 36 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=5.18 $Y=2
+ $X2=5.335 $Y2=1.915
r144 33 34 115.802 $w=1.68e-07 $l=1.775e-06 $layer=LI1_cond $X=5.18 $Y=2
+ $X2=3.405 $Y2=2
r145 29 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=1.86
r146 29 31 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.295 $Y=2.085
+ $X2=3.295 $Y2=2.205
r147 25 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.295 $Y=1.635
+ $X2=3.295 $Y2=1.86
r148 25 27 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=3.295 $Y=1.635
+ $X2=3.295 $Y2=0.42
r149 23 42 3.05 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.185 $Y=1.77
+ $X2=3.295 $Y2=1.86
r150 23 41 27.3172 $w=2.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.185 $Y=1.77
+ $X2=2.545 $Y2=1.77
r151 19 55 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.575 $Y=1.655
+ $X2=5.575 $Y2=1.52
r152 19 21 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.575 $Y=1.655
+ $X2=5.575 $Y2=2.165
r153 15 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.435 $Y=1.385
+ $X2=5.435 $Y2=1.52
r154 15 17 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.435 $Y=1.385
+ $X2=5.435 $Y2=0.445
r155 13 50 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.51 $Y=0.445
+ $X2=2.51 $Y2=1.575
r156 9 51 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.43 $Y=2.275
+ $X2=2.43 $Y2=1.905
r157 2 31 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=2.205
r158 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.235 $X2=3.32 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_287_413# 1 2 7 9 12 14 18 23 25 26 28 35
c99 28 0 1.77265e-19 $X=2.93 $Y=1.16
c100 26 0 3.17216e-20 $X=2.5 $Y=1.185
c101 25 0 3.18278e-20 $X=2.415 $Y=0.995
c102 14 0 2.67301e-20 $X=2.33 $Y=0.395
r103 31 32 14.6301 $w=2.46e-07 $l=2.95e-07 $layer=LI1_cond $X=2.12 $Y=1.205
+ $X2=2.415 $Y2=1.205
r104 29 35 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.93 $Y=1.16
+ $X2=3.11 $Y2=1.16
r105 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.16 $X2=2.93 $Y2=1.16
r106 26 32 4.2431 $w=3.8e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.5 $Y=1.185
+ $X2=2.415 $Y2=1.205
r107 26 28 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.5 $Y=1.185
+ $X2=2.93 $Y2=1.185
r108 25 32 2.90119 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.415 $Y=0.995
+ $X2=2.415 $Y2=1.205
r109 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.415 $Y=0.535
+ $X2=2.415 $Y2=0.995
r110 22 31 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.12 $Y=1.375
+ $X2=2.12 $Y2=1.205
r111 22 23 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.12 $Y=1.375
+ $X2=2.12 $Y2=2.125
r112 18 23 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.035 $Y=2.295
+ $X2=2.12 $Y2=2.125
r113 18 20 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.035 $Y=2.295
+ $X2=1.6 $Y2=2.295
r114 14 24 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.33 $Y=0.395
+ $X2=2.415 $Y2=0.535
r115 14 16 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=2.33 $Y=0.395
+ $X2=1.635 $Y2=0.395
r116 10 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r117 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r118 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r119 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=0.56
r120 2 20 600 $w=1.7e-07 $l=3.22102e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=2.065 $X2=1.6 $Y2=2.315
r121 1 16 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.635 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%CLK 3 5 8 11 15 17 18 21 24 27 29 33 38
c80 38 0 1.86451e-19 $X=4.925 $Y=1.14
c81 29 0 1.20889e-19 $X=4.715 $Y=1.325
c82 21 0 3.68683e-20 $X=5.885 $Y=1.05
c83 18 0 1.33567e-19 $X=4.66 $Y=0.88
c84 15 0 2.24995e-19 $X=5.995 $Y=2.165
r85 27 29 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.715 $Y=1.16
+ $X2=4.715 $Y2=1.325
r86 24 38 4.54172 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.79 $Y=1.14
+ $X2=4.925 $Y2=1.14
r87 24 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r88 22 33 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=5.885 $Y=1.05
+ $X2=5.995 $Y2=1.05
r89 22 30 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.885 $Y=1.05
+ $X2=5.795 $Y2=1.05
r90 21 38 35.6886 $w=3.08e-07 $l=9.6e-07 $layer=LI1_cond $X=5.885 $Y=1.11
+ $X2=4.925 $Y2=1.11
r91 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.885
+ $Y=1.05 $X2=5.885 $Y2=1.05
r92 17 18 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.66 $Y=0.73
+ $X2=4.66 $Y2=0.88
r93 13 33 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.995 $Y=1.185
+ $X2=5.995 $Y2=1.05
r94 13 15 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=5.995 $Y=1.185
+ $X2=5.995 $Y2=2.165
r95 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.795 $Y=0.915
+ $X2=5.795 $Y2=1.05
r96 9 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.795 $Y=0.915 $X2=5.795
+ $Y2=0.445
r97 8 29 163.88 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.635 $Y=1.835
+ $X2=4.635 $Y2=1.325
r98 5 27 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=4.715 $Y=1.115
+ $X2=4.715 $Y2=1.16
r99 5 18 31.1181 $w=4.2e-07 $l=2.35e-07 $layer=POLY_cond $X=4.715 $Y=1.115
+ $X2=4.715 $Y2=0.88
r100 3 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.47 $Y=0.445
+ $X2=4.47 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_1020_47# 1 2 7 9 12 14 16 19 23 25 26 27
+ 31 38
c82 7 0 3.68683e-20 $X=6.47 $Y=0.995
r83 37 38 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.47 $Y=1.16
+ $X2=6.89 $Y2=1.16
r84 34 37 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.415 $Y=1.16
+ $X2=6.47 $Y2=1.16
r85 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.16 $X2=6.415 $Y2=1.16
r86 31 33 9.57218 $w=4.78e-07 $l=2.09105e-07 $layer=LI1_cond $X=6.315 $Y=0.995
+ $X2=6.415 $Y2=1.16
r87 30 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.315 $Y=0.785
+ $X2=6.315 $Y2=0.995
r88 27 33 28.9697 $w=4.78e-07 $l=1.19932e-06 $layer=LI1_cond $X=5.785 $Y=2.085
+ $X2=6.415 $Y2=1.16
r89 27 29 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=5.785 $Y=2.085
+ $X2=5.785 $Y2=2.125
r90 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.23 $Y=0.7
+ $X2=6.315 $Y2=0.785
r91 25 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=6.23 $Y=0.7 $X2=5.31
+ $Y2=0.7
r92 21 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.205 $Y=0.615
+ $X2=5.31 $Y2=0.7
r93 21 23 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=5.205 $Y=0.615
+ $X2=5.205 $Y2=0.46
r94 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.16
r95 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.89 $Y=1.325
+ $X2=6.89 $Y2=1.985
r96 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=1.16
r97 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.89 $Y=0.995
+ $X2=6.89 $Y2=0.56
r98 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=1.325
+ $X2=6.47 $Y2=1.16
r99 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.47 $Y=1.325
+ $X2=6.47 $Y2=1.985
r100 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=0.995
+ $X2=6.47 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.47 $Y=0.995
+ $X2=6.47 $Y2=0.56
r102 2 29 600 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=1 $X=5.65
+ $Y=1.845 $X2=5.785 $Y2=2.125
r103 1 23 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.1
+ $Y=0.235 $X2=5.225 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%VPWR 1 2 3 4 5 6 19 21 25 27 29 33 35 36
+ 50 56 61 72 75 81 83 87
r98 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r99 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r100 80 81 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=2.53
+ $X2=5.53 $Y2=2.53
r101 77 80 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=5.29 $Y=2.53
+ $X2=5.365 $Y2=2.53
r102 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r103 74 75 11.8978 $w=7.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.795 $Y=2.44
+ $X2=3.015 $Y2=2.44
r104 70 74 4.34193 $w=7.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.795 $Y2=2.44
r105 70 72 10.8328 $w=7.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.375 $Y2=2.44
r106 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 65 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r108 65 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r109 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r110 62 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.4 $Y=2.72
+ $X2=6.235 $Y2=2.72
r111 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.4 $Y=2.72 $X2=6.67
+ $Y2=2.72
r112 61 86 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.185 $Y2=2.72
r113 61 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r114 60 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 60 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 59 81 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.53 $Y2=2.72
r117 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r118 56 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.07 $Y=2.72
+ $X2=6.235 $Y2=2.72
r119 56 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.07 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 53 78 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r121 52 55 9.7861 $w=5.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=4.36 $Y2=2.53
r122 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r123 50 77 0.761141 $w=5.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.255 $Y=2.53
+ $X2=5.29 $Y2=2.53
r124 50 55 19.4635 $w=5.48e-07 $l=8.95e-07 $layer=LI1_cond $X=5.255 $Y=2.53
+ $X2=4.36 $Y2=2.53
r125 49 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r126 49 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r127 48 75 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.015 $Y2=2.72
r128 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r129 45 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 44 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.375 $Y2=2.72
r131 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 42 45 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r133 41 44 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 39 67 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r136 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r137 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 36 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r139 35 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 33 52 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=3.85 $Y=2.53 $X2=3.91
+ $Y2=2.53
r141 33 35 12.2241 $w=5.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.85 $Y=2.53
+ $X2=3.575 $Y2=2.53
r142 29 32 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=7.142 $Y=1.66
+ $X2=7.142 $Y2=2.34
r143 27 86 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=7.142 $Y=2.635
+ $X2=7.185 $Y2=2.72
r144 27 32 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.142 $Y=2.635
+ $X2=7.142 $Y2=2.34
r145 23 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.235 $Y=2.635
+ $X2=6.235 $Y2=2.72
r146 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.235 $Y=2.635
+ $X2=6.235 $Y2=2.36
r147 19 67 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r148 19 21 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r149 6 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=2.34
r150 6 29 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.965
+ $Y=1.485 $X2=7.1 $Y2=1.66
r151 5 25 600 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.845 $X2=6.235 $Y2=2.36
r152 4 80 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=5.24
+ $Y=1.845 $X2=5.365 $Y2=2.34
r153 3 55 600 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=4.16
+ $Y=1.515 $X2=4.36 $Y2=2.34
r154 2 74 600 $w=1.7e-07 $l=4.15421e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=2.065 $X2=2.795 $Y2=2.36
r155 1 21 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%A_27_47# 1 2 3 12 15 16 17 18 20 24
r49 22 24 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.105 $Y=0.615
+ $X2=1.105 $Y2=0.42
r50 18 20 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=0.685 $Y=2.295
+ $X2=1.095 $Y2=2.295
r51 17 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.7 $X2=0.6
+ $Y2=0.7
r52 16 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=1.105 $Y2=0.615
r53 16 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.015 $Y=0.7
+ $X2=0.685 $Y2=0.7
r54 15 18 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.6 $Y=2.125
+ $X2=0.685 $Y2=2.295
r55 14 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=0.785 $X2=0.6
+ $Y2=0.7
r56 14 15 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=0.6 $Y=0.785
+ $X2=0.6 $Y2=2.125
r57 10 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.6 $Y2=0.7
r58 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r59 3 20 600 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.845 $X2=1.095 $Y2=2.29
r60 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%GCLK 1 2 8 12 13 14 16 17 18 19 20 26 37
r30 20 37 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=7.19 $Y=1.185 $X2=7.13
+ $Y2=1.185
r31 18 19 16.8598 $w=2.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.705 $Y=1.815
+ $X2=6.705 $Y2=2.21
r32 17 26 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=6.705 $Y=0.51
+ $X2=6.705 $Y2=0.42
r33 15 37 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=6.84 $Y=1.185
+ $X2=7.13 $Y2=1.185
r34 15 16 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=1.185
+ $X2=6.755 $Y2=1.185
r35 13 18 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.705 $Y=1.63
+ $X2=6.705 $Y2=1.815
r36 13 14 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=1.63
+ $X2=6.705 $Y2=1.495
r37 11 17 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.705 $Y=0.69
+ $X2=6.705 $Y2=0.51
r38 11 12 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=0.69
+ $X2=6.705 $Y2=0.825
r39 9 16 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.755 $Y=1.315
+ $X2=6.755 $Y2=1.185
r40 9 14 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.755 $Y=1.315
+ $X2=6.755 $Y2=1.495
r41 8 16 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.755 $Y=1.055
+ $X2=6.755 $Y2=1.185
r42 8 12 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.755 $Y=1.055
+ $X2=6.755 $Y2=0.825
r43 2 18 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=6.545
+ $Y=1.485 $X2=6.68 $Y2=1.815
r44 1 26 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.545
+ $Y=0.235 $X2=6.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__SDLCLKP_2%VGND 1 2 3 4 5 18 22 26 28 30 32 34 39 47
+ 57 63 66 69 73 77 80
r109 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r110 75 77 10.2686 $w=5.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.21 $Y=0.18
+ $X2=6.4 $Y2=0.18
r111 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r112 72 75 1.46689 $w=5.28e-07 $l=6.5e-08 $layer=LI1_cond $X=6.145 $Y=0.18
+ $X2=6.21 $Y2=0.18
r113 72 73 20.7625 $w=5.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6.145 $Y=0.18
+ $X2=5.49 $Y2=0.18
r114 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r115 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r116 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r117 61 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r118 61 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=6.21
+ $Y2=0
r119 60 77 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.4
+ $Y2=0
r120 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r121 57 79 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.01 $Y=0 $X2=7.185
+ $Y2=0
r122 57 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=0 $X2=6.67
+ $Y2=0
r123 56 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r124 56 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r125 55 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=5.49
+ $Y2=0
r126 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r127 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.26
+ $Y2=0
r128 53 55 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=4.425 $Y=0
+ $X2=5.29 $Y2=0
r129 51 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r130 51 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r131 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r132 48 66 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.015 $Y=0
+ $X2=2.842 $Y2=0
r133 48 50 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.015 $Y=0
+ $X2=3.91 $Y2=0
r134 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=4.26
+ $Y2=0
r135 47 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=3.91 $Y2=0
r136 46 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r137 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r138 43 46 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r139 43 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r140 42 45 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r141 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r142 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r143 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r144 39 66 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.842
+ $Y2=0
r145 39 45 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.67 $Y=0 $X2=2.53
+ $Y2=0
r146 34 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r147 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r148 32 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r149 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r150 28 79 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=7.142 $Y=0.085
+ $X2=7.185 $Y2=0
r151 28 30 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=7.142 $Y=0.085
+ $X2=7.142 $Y2=0.38
r152 24 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0
r153 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.26 $Y=0.085
+ $X2=4.26 $Y2=0.36
r154 20 66 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0
r155 20 22 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=2.842 $Y=0.085
+ $X2=2.842 $Y2=0.51
r156 16 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r157 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r158 5 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.965
+ $Y=0.235 $X2=7.1 $Y2=0.38
r159 4 72 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.145 $Y2=0.36
r160 3 26 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.125
+ $Y=0.235 $X2=4.26 $Y2=0.36
r161 2 22 182 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.815 $Y2=0.51
r162 1 18 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


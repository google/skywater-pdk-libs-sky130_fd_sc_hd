* File: sky130_fd_sc_hd__o311a_4.pxi.spice
* Created: Tue Sep  1 19:24:33 2020
* 
x_PM_SKY130_FD_SC_HD__O311A_4%A_79_21# N_A_79_21#_M1013_s N_A_79_21#_M1018_s
+ N_A_79_21#_M1008_s N_A_79_21#_M1004_s N_A_79_21#_c_128_n N_A_79_21#_M1012_g
+ N_A_79_21#_M1002_g N_A_79_21#_c_129_n N_A_79_21#_M1017_g N_A_79_21#_M1005_g
+ N_A_79_21#_c_130_n N_A_79_21#_M1019_g N_A_79_21#_M1020_g N_A_79_21#_c_131_n
+ N_A_79_21#_M1025_g N_A_79_21#_M1024_g N_A_79_21#_c_219_p N_A_79_21#_c_132_n
+ N_A_79_21#_c_142_n N_A_79_21#_c_235_p N_A_79_21#_c_149_p N_A_79_21#_c_180_p
+ N_A_79_21#_c_133_n N_A_79_21#_c_134_n N_A_79_21#_c_194_p N_A_79_21#_c_153_p
+ N_A_79_21#_c_196_p N_A_79_21#_c_143_n N_A_79_21#_c_234_p N_A_79_21#_c_135_n
+ N_A_79_21#_c_136_n N_A_79_21#_c_137_n N_A_79_21#_c_145_n N_A_79_21#_c_146_n
+ PM_SKY130_FD_SC_HD__O311A_4%A_79_21#
x_PM_SKY130_FD_SC_HD__O311A_4%C1 N_C1_M1018_g N_C1_c_266_n N_C1_M1013_g
+ N_C1_M1021_g N_C1_c_268_n N_C1_M1015_g C1 C1 N_C1_c_270_n
+ PM_SKY130_FD_SC_HD__O311A_4%C1
x_PM_SKY130_FD_SC_HD__O311A_4%B1 N_B1_c_322_n N_B1_M1008_g N_B1_c_318_n
+ N_B1_M1007_g N_B1_c_323_n N_B1_M1011_g N_B1_c_319_n N_B1_M1009_g B1 B1 B1
+ N_B1_c_321_n PM_SKY130_FD_SC_HD__O311A_4%B1
x_PM_SKY130_FD_SC_HD__O311A_4%A3 N_A3_M1004_g N_A3_M1000_g N_A3_M1016_g
+ N_A3_M1010_g N_A3_c_367_n A3 A3 A3 N_A3_c_369_n PM_SKY130_FD_SC_HD__O311A_4%A3
x_PM_SKY130_FD_SC_HD__O311A_4%A2 N_A2_M1022_g N_A2_M1006_g N_A2_M1023_g
+ N_A2_M1014_g A2 A2 N_A2_c_417_n PM_SKY130_FD_SC_HD__O311A_4%A2
x_PM_SKY130_FD_SC_HD__O311A_4%A1 N_A1_M1001_g N_A1_M1003_g N_A1_M1027_g
+ N_A1_M1026_g A1 A1 N_A1_c_463_n PM_SKY130_FD_SC_HD__O311A_4%A1
x_PM_SKY130_FD_SC_HD__O311A_4%VPWR N_VPWR_M1002_s N_VPWR_M1005_s N_VPWR_M1024_s
+ N_VPWR_M1021_d N_VPWR_M1011_d N_VPWR_M1003_d N_VPWR_c_499_n N_VPWR_c_500_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n N_VPWR_c_507_n VPWR N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_498_n N_VPWR_c_513_n N_VPWR_c_514_n
+ N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n PM_SKY130_FD_SC_HD__O311A_4%VPWR
x_PM_SKY130_FD_SC_HD__O311A_4%X N_X_M1012_s N_X_M1019_s N_X_M1002_d N_X_M1020_d
+ N_X_c_614_n N_X_c_617_n N_X_c_641_n N_X_c_626_n N_X_c_618_n N_X_c_645_n
+ N_X_c_654_p N_X_c_615_n N_X_c_635_n N_X_c_616_n X
+ PM_SKY130_FD_SC_HD__O311A_4%X
x_PM_SKY130_FD_SC_HD__O311A_4%A_875_297# N_A_875_297#_M1004_d
+ N_A_875_297#_M1016_d N_A_875_297#_M1006_s N_A_875_297#_c_660_n
+ N_A_875_297#_c_667_n N_A_875_297#_c_661_n N_A_875_297#_c_662_n
+ N_A_875_297#_c_663_n N_A_875_297#_c_680_n N_A_875_297#_c_664_n
+ PM_SKY130_FD_SC_HD__O311A_4%A_875_297#
x_PM_SKY130_FD_SC_HD__O311A_4%A_1147_297# N_A_1147_297#_M1006_d
+ N_A_1147_297#_M1014_d N_A_1147_297#_M1026_s N_A_1147_297#_c_706_n
+ N_A_1147_297#_c_713_n N_A_1147_297#_c_707_n N_A_1147_297#_c_725_n
+ N_A_1147_297#_c_708_n N_A_1147_297#_c_709_n N_A_1147_297#_c_710_n
+ PM_SKY130_FD_SC_HD__O311A_4%A_1147_297#
x_PM_SKY130_FD_SC_HD__O311A_4%VGND N_VGND_M1012_d N_VGND_M1017_d N_VGND_M1025_d
+ N_VGND_M1000_s N_VGND_M1022_s N_VGND_M1001_d N_VGND_c_742_n N_VGND_c_743_n
+ N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n
+ N_VGND_c_749_n VGND N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n
+ N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n N_VGND_c_757_n
+ N_VGND_c_758_n N_VGND_c_759_n PM_SKY130_FD_SC_HD__O311A_4%VGND
x_PM_SKY130_FD_SC_HD__O311A_4%A_467_47# N_A_467_47#_M1013_d N_A_467_47#_M1015_d
+ N_A_467_47#_M1009_d N_A_467_47#_c_868_n N_A_467_47#_c_869_n
+ N_A_467_47#_c_870_n N_A_467_47#_c_890_n PM_SKY130_FD_SC_HD__O311A_4%A_467_47#
x_PM_SKY130_FD_SC_HD__O311A_4%A_717_47# N_A_717_47#_M1007_s N_A_717_47#_M1000_d
+ N_A_717_47#_M1010_d N_A_717_47#_M1023_d N_A_717_47#_M1027_s
+ N_A_717_47#_c_896_n N_A_717_47#_c_908_n N_A_717_47#_c_915_n
+ N_A_717_47#_c_920_n N_A_717_47#_c_897_n N_A_717_47#_c_898_n
+ N_A_717_47#_c_899_n N_A_717_47#_c_900_n PM_SKY130_FD_SC_HD__O311A_4%A_717_47#
cc_1 VNB N_A_79_21#_c_128_n 0.0210045f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_129_n 0.0156962f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_130_n 0.0157154f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_131_n 0.0187698f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_132_n 0.00147908f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.055
cc_6 VNB N_A_79_21#_c_133_n 0.00305942f $X=-0.19 $Y=-0.24 $X2=2.3 $Y2=0.78
cc_7 VNB N_A_79_21#_c_134_n 7.99934e-19 $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.76
cc_8 VNB N_A_79_21#_c_135_n 0.00170727f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_9 VNB N_A_79_21#_c_136_n 0.0778587f $X=-0.19 $Y=-0.24 $X2=1.78 $Y2=1.16
cc_10 VNB N_A_79_21#_c_137_n 0.00389371f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=0.78
cc_11 VNB N_C1_M1018_g 3.83136e-19 $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=1.485
cc_12 VNB N_C1_c_266_n 0.017934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_C1_M1021_g 3.23752e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_C1_c_268_n 0.0144176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB C1 0.00485721f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_16 VNB N_C1_c_270_n 0.0587162f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_17 VNB N_B1_c_318_n 0.016229f $X=-0.19 $Y=-0.24 $X2=4.785 $Y2=1.485
cc_18 VNB N_B1_c_319_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB B1 0.0121465f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_20 VNB N_B1_c_321_n 0.0404816f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_21 VNB N_A3_M1004_g 5.14727e-19 $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=1.485
cc_22 VNB N_A3_M1000_g 0.0269785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A3_M1016_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A3_M1010_g 0.0204257f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_25 VNB N_A3_c_367_n 0.0398335f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_26 VNB A3 0.00266544f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_27 VNB N_A3_c_369_n 0.0355083f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_28 VNB N_A2_M1022_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=1.485
cc_29 VNB N_A2_M1006_g 4.5691e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A2_M1023_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A2_M1014_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_32 VNB A2 0.0036164f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_33 VNB N_A2_c_417_n 0.029894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A1_M1001_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=1.485
cc_35 VNB N_A1_M1003_g 4.25212e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A1_M1027_g 0.0232752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB A1 0.0112033f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_38 VNB N_A1_c_463_n 0.0478197f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_39 VNB N_VPWR_c_498_n 0.326667f $X=-0.19 $Y=-0.24 $X2=4.92 $Y2=1.815
cc_40 VNB N_X_c_614_n 0.00197742f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_41 VNB N_X_c_615_n 0.0141924f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_42 VNB N_X_c_616_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_43 VNB N_VGND_c_742_n 0.0102094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_743_n 0.0305153f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_45 VNB N_VGND_c_744_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_46 VNB N_VGND_c_745_n 0.00227952f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_47 VNB N_VGND_c_746_n 3.01556e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_747_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_49 VNB N_VGND_c_748_n 0.0118385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_749_n 0.0035381f $X=-0.19 $Y=-0.24 $X2=1.775 $Y2=1.185
cc_51 VNB N_VGND_c_750_n 0.0118385f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.16
cc_52 VNB N_VGND_c_751_n 0.0110732f $X=-0.19 $Y=-0.24 $X2=2.7 $Y2=1.815
cc_53 VNB N_VGND_c_752_n 0.0110791f $X=-0.19 $Y=-0.24 $X2=3.54 $Y2=1.815
cc_54 VNB N_VGND_c_753_n 0.0147997f $X=-0.19 $Y=-0.24 $X2=4.92 $Y2=1.815
cc_55 VNB N_VGND_c_754_n 0.376468f $X=-0.19 $Y=-0.24 $X2=1.86 $Y2=1.185
cc_56 VNB N_VGND_c_755_n 0.00436611f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_57 VNB N_VGND_c_756_n 0.0662108f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_58 VNB N_VGND_c_757_n 0.0124189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_758_n 0.0043639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_759_n 0.0043639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_467_47#_c_868_n 0.0052638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_467_47#_c_869_n 0.00135245f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_63 VNB N_A_467_47#_c_870_n 0.00287235f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_64 VNB N_A_717_47#_c_896_n 0.00653008f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_65 VNB N_A_717_47#_c_897_n 0.00905088f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_66 VNB N_A_717_47#_c_898_n 0.00207541f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_67 VNB N_A_717_47#_c_899_n 0.00151868f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_68 VNB N_A_717_47#_c_900_n 0.0279707f $X=-0.19 $Y=-0.24 $X2=1.775 $Y2=1.185
cc_69 VPB N_A_79_21#_M1002_g 0.0249926f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_70 VPB N_A_79_21#_M1005_g 0.0181826f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_71 VPB N_A_79_21#_M1020_g 0.0182107f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_72 VPB N_A_79_21#_M1024_g 0.02034f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_73 VPB N_A_79_21#_c_142_n 0.00198493f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.485
cc_74 VPB N_A_79_21#_c_143_n 0.0157355f $X=-0.19 $Y=1.305 $X2=4.835 $Y2=1.605
cc_75 VPB N_A_79_21#_c_136_n 0.0154697f $X=-0.19 $Y=1.305 $X2=1.78 $Y2=1.16
cc_76 VPB N_A_79_21#_c_145_n 0.00117749f $X=-0.19 $Y=1.305 $X2=2.7 $Y2=1.605
cc_77 VPB N_A_79_21#_c_146_n 0.00115444f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=1.605
cc_78 VPB N_C1_M1018_g 0.0224627f $X=-0.19 $Y=1.305 $X2=3.405 $Y2=1.485
cc_79 VPB N_C1_M1021_g 0.0195099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB C1 0.00626145f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_81 VPB N_B1_c_322_n 0.0141141f $X=-0.19 $Y=1.305 $X2=2.745 $Y2=0.235
cc_82 VPB N_B1_c_323_n 0.0190993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB B1 0.00460016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_84 VPB N_B1_c_321_n 0.0213427f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_85 VPB N_A3_M1004_g 0.0271907f $X=-0.19 $Y=1.305 $X2=3.405 $Y2=1.485
cc_86 VPB N_A3_M1016_g 0.0274617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB A3 0.0158394f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_88 VPB N_A2_M1006_g 0.0273218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A2_M1014_g 0.019782f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_90 VPB A2 0.00444715f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_91 VPB N_A1_M1003_g 0.0196045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A1_M1026_g 0.027097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_93 VPB A1 0.00591402f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_94 VPB N_A1_c_463_n 0.00614837f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_95 VPB N_VPWR_c_499_n 0.0101835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_500_n 0.0442414f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_97 VPB N_VPWR_c_501_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_98 VPB N_VPWR_c_502_n 0.0016795f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_99 VPB N_VPWR_c_503_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_504_n 3.12367e-19 $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.325
cc_101 VPB N_VPWR_c_505_n 0.0154476f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_102 VPB N_VPWR_c_506_n 0.00420258f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.16
cc_103 VPB N_VPWR_c_507_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.86 $Y2=1.055
cc_104 VPB N_VPWR_c_508_n 0.0124915f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=0.8
cc_105 VPB N_VPWR_c_509_n 0.0124915f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.76
cc_106 VPB N_VPWR_c_510_n 0.0702985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_511_n 0.0154931f $X=-0.19 $Y=1.305 $X2=4.92 $Y2=1.815
cc_108 VPB N_VPWR_c_498_n 0.0568917f $X=-0.19 $Y=1.305 $X2=4.92 $Y2=1.815
cc_109 VPB N_VPWR_c_513_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.54 $Y2=1.605
cc_110 VPB N_VPWR_c_514_n 0.0103759f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_111 VPB N_VPWR_c_515_n 0.00436868f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_112 VPB N_VPWR_c_516_n 0.00362871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_517_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_X_c_617_n 0.0028845f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_115 VPB N_X_c_618_n 0.00116994f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_116 VPB N_X_c_615_n 0.00326378f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_117 VPB N_A_875_297#_c_660_n 0.00443643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_875_297#_c_661_n 0.00204172f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_119 VPB N_A_875_297#_c_662_n 0.00962232f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_120 VPB N_A_875_297#_c_663_n 0.00898483f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_121 VPB N_A_875_297#_c_664_n 8.14146e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_1147_297#_c_706_n 0.00376319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_1147_297#_c_707_n 0.00489414f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_124 VPB N_A_1147_297#_c_708_n 0.0124504f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_125 VPB N_A_1147_297#_c_709_n 0.0293809f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_126 VPB N_A_1147_297#_c_710_n 0.0015191f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_127 N_A_79_21#_M1024_g N_C1_M1018_g 0.00946607f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_142_n N_C1_M1018_g 0.00267492f $X=1.86 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_149_p N_C1_M1018_g 0.0175453f $X=2.615 $Y=1.605 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_136_n N_C1_M1018_g 7.28283e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_132_n N_C1_c_266_n 0.00154333f $X=1.86 $Y=1.055 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_134_n N_C1_c_266_n 0.0119265f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_153_p N_C1_M1021_g 0.015604f $X=3.455 $Y=1.605 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_134_n N_C1_c_268_n 0.00297649f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_149_p C1 0.0341351f $X=2.615 $Y=1.605 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_153_p C1 0.018063f $X=3.455 $Y=1.605 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_135_n C1 0.0230019f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_136_n C1 0.00110264f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_137_n C1 0.0625269f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_145_n C1 0.013857f $X=2.7 $Y=1.605 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_131_n N_C1_c_270_n 6.75522e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_132_n N_C1_c_270_n 0.00111023f $X=1.86 $Y=1.055 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_149_p N_C1_c_270_n 5.19546e-19 $X=2.615 $Y=1.605 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_134_n N_C1_c_270_n 0.0102359f $X=2.88 $Y=0.76 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_153_p N_C1_c_270_n 0.00326608f $X=3.455 $Y=1.605 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_135_n N_C1_c_270_n 2.19242e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_136_n N_C1_c_270_n 0.009921f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_145_n N_C1_c_270_n 6.67081e-19 $X=2.7 $Y=1.605 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_153_p N_B1_c_322_n 0.015604f $X=3.455 $Y=1.605 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_79_21#_c_143_n N_B1_c_323_n 0.0195789f $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_153_p B1 0.0127963f $X=3.455 $Y=1.605 $X2=0 $Y2=0
cc_152 N_A_79_21#_c_143_n B1 0.0610748f $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_146_n B1 0.0131805f $X=3.54 $Y=1.605 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_143_n N_B1_c_321_n 0.00483899f $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_146_n N_B1_c_321_n 0.00274773f $X=3.54 $Y=1.605 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_143_n N_A3_M1004_g 0.016161f $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_143_n A3 0.0251507f $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_143_n N_A3_c_369_n 6.60094e-19 $X=4.835 $Y=1.605 $X2=0 $Y2=0
cc_159 N_A_79_21#_c_149_p N_VPWR_M1024_s 0.0132663f $X=2.615 $Y=1.605 $X2=0
+ $Y2=0
cc_160 N_A_79_21#_c_180_p N_VPWR_M1024_s 9.18498e-19 $X=1.945 $Y=1.605 $X2=0
+ $Y2=0
cc_161 N_A_79_21#_c_153_p N_VPWR_M1021_d 0.00452889f $X=3.455 $Y=1.605 $X2=0
+ $Y2=0
cc_162 N_A_79_21#_c_143_n N_VPWR_M1011_d 0.00626324f $X=4.835 $Y=1.605 $X2=0
+ $Y2=0
cc_163 N_A_79_21#_M1002_g N_VPWR_c_500_n 0.0157787f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_79_21#_M1005_g N_VPWR_c_500_n 8.36313e-19 $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_79_21#_M1002_g N_VPWR_c_501_n 6.54417e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_79_21#_M1005_g N_VPWR_c_501_n 0.0104025f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_79_21#_M1020_g N_VPWR_c_501_n 0.0104025f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_79_21#_M1024_g N_VPWR_c_501_n 6.54417e-19 $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_A_79_21#_M1020_g N_VPWR_c_502_n 6.67793e-19 $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_A_79_21#_M1024_g N_VPWR_c_502_n 0.0114196f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_149_p N_VPWR_c_502_n 0.0365821f $X=2.615 $Y=1.605 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_c_180_p N_VPWR_c_502_n 0.00989598f $X=1.945 $Y=1.605 $X2=0
+ $Y2=0
cc_173 N_A_79_21#_c_136_n N_VPWR_c_502_n 4.01766e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_194_p N_VPWR_c_503_n 0.0113958f $X=2.7 $Y=1.815 $X2=0 $Y2=0
cc_175 N_A_79_21#_c_153_p N_VPWR_c_504_n 0.017435f $X=3.455 $Y=1.605 $X2=0 $Y2=0
cc_176 N_A_79_21#_c_196_p N_VPWR_c_505_n 0.0113958f $X=3.54 $Y=1.815 $X2=0 $Y2=0
cc_177 N_A_79_21#_c_143_n N_VPWR_c_506_n 0.0134934f $X=4.835 $Y=1.605 $X2=0
+ $Y2=0
cc_178 N_A_79_21#_M1002_g N_VPWR_c_508_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_79_21#_M1005_g N_VPWR_c_508_n 0.0046653f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A_79_21#_M1020_g N_VPWR_c_509_n 0.0046653f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_79_21#_M1024_g N_VPWR_c_509_n 0.0046653f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A_79_21#_M1018_s N_VPWR_c_498_n 0.00570907f $X=2.565 $Y=1.485 $X2=0
+ $Y2=0
cc_183 N_A_79_21#_M1008_s N_VPWR_c_498_n 0.00570907f $X=3.405 $Y=1.485 $X2=0
+ $Y2=0
cc_184 N_A_79_21#_M1004_s N_VPWR_c_498_n 0.00216833f $X=4.785 $Y=1.485 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_M1002_g N_VPWR_c_498_n 0.00796766f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_79_21#_M1005_g N_VPWR_c_498_n 0.00796766f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_M1020_g N_VPWR_c_498_n 0.00796766f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_79_21#_M1024_g N_VPWR_c_498_n 0.00796766f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_79_21#_c_194_p N_VPWR_c_498_n 0.00646998f $X=2.7 $Y=1.815 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_196_p N_VPWR_c_498_n 0.00646998f $X=3.54 $Y=1.815 $X2=0
+ $Y2=0
cc_191 N_A_79_21#_c_128_n N_X_c_614_n 0.00260329f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_129_n N_X_c_614_n 0.00259917f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_136_n N_X_c_614_n 0.00805828f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_79_21#_M1002_g N_X_c_617_n 0.00379746f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_79_21#_M1005_g N_X_c_617_n 0.00379746f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_196 N_A_79_21#_c_136_n N_X_c_617_n 0.00310634f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_79_21#_c_129_n N_X_c_626_n 0.0112109f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_79_21#_c_130_n N_X_c_626_n 0.00967544f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_79_21#_c_219_p N_X_c_626_n 0.0298197f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_200 N_A_79_21#_c_136_n N_X_c_626_n 0.0021659f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_79_21#_M1005_g N_X_c_618_n 0.0167612f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_79_21#_M1020_g N_X_c_618_n 0.015224f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_79_21#_c_219_p N_X_c_618_n 0.0436667f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_204 N_A_79_21#_c_136_n N_X_c_618_n 0.00418025f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_79_21#_c_136_n N_X_c_615_n 0.0266688f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_79_21#_c_219_p N_X_c_635_n 0.0218399f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_207 N_A_79_21#_c_136_n N_X_c_635_n 0.0078907f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_219_p N_X_c_616_n 0.0131017f $X=1.775 $Y=1.185 $X2=0 $Y2=0
cc_209 N_A_79_21#_c_136_n N_X_c_616_n 0.00224547f $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_79_21#_c_143_n N_A_875_297#_M1004_d 0.00638585f $X=4.835 $Y=1.605
+ $X2=-0.19 $Y2=-0.24
cc_211 N_A_79_21#_c_143_n N_A_875_297#_c_660_n 0.0221881f $X=4.835 $Y=1.605
+ $X2=0 $Y2=0
cc_212 N_A_79_21#_M1004_s N_A_875_297#_c_667_n 0.00312348f $X=4.785 $Y=1.485
+ $X2=0 $Y2=0
cc_213 N_A_79_21#_c_143_n N_A_875_297#_c_667_n 0.0030597f $X=4.835 $Y=1.605
+ $X2=0 $Y2=0
cc_214 N_A_79_21#_c_234_p N_A_875_297#_c_667_n 0.011831f $X=4.92 $Y=1.725 $X2=0
+ $Y2=0
cc_215 N_A_79_21#_c_235_p N_VGND_M1025_d 8.94971e-19 $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_216 N_A_79_21#_c_137_n N_VGND_M1025_d 0.00423301f $X=2.195 $Y=0.78 $X2=0
+ $Y2=0
cc_217 N_A_79_21#_c_128_n N_VGND_c_743_n 0.0121301f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_129_n N_VGND_c_743_n 6.22847e-19 $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_79_21#_c_128_n N_VGND_c_744_n 5.71893e-19 $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_79_21#_c_129_n N_VGND_c_744_n 0.00748092f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_79_21#_c_130_n N_VGND_c_744_n 0.00748092f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_79_21#_c_131_n N_VGND_c_744_n 5.71893e-19 $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_79_21#_c_130_n N_VGND_c_745_n 5.66483e-19 $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_79_21#_c_131_n N_VGND_c_745_n 0.00840497f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_79_21#_c_235_p N_VGND_c_745_n 0.00946546f $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_226 N_A_79_21#_c_136_n N_VGND_c_745_n 4.90038e-19 $X=1.78 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_79_21#_c_137_n N_VGND_c_745_n 0.00613389f $X=2.195 $Y=0.78 $X2=0
+ $Y2=0
cc_228 N_A_79_21#_c_130_n N_VGND_c_748_n 0.00348405f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_229 N_A_79_21#_c_131_n N_VGND_c_748_n 0.0046653f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_79_21#_c_128_n N_VGND_c_750_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_79_21#_c_129_n N_VGND_c_750_n 0.00348405f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_79_21#_M1013_s N_VGND_c_754_n 0.00216833f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_A_79_21#_c_128_n N_VGND_c_754_n 0.00796766f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_79_21#_c_129_n N_VGND_c_754_n 0.00414556f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_79_21#_c_130_n N_VGND_c_754_n 0.00414556f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_79_21#_c_131_n N_VGND_c_754_n 0.00796766f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_79_21#_c_235_p N_VGND_c_754_n 7.30854e-19 $X=1.945 $Y=0.8 $X2=0 $Y2=0
cc_238 N_A_79_21#_c_137_n N_VGND_c_754_n 0.0048636f $X=2.195 $Y=0.78 $X2=0 $Y2=0
cc_239 N_A_79_21#_c_137_n N_VGND_c_756_n 0.00259545f $X=2.195 $Y=0.78 $X2=0
+ $Y2=0
cc_240 N_A_79_21#_c_134_n N_A_467_47#_M1013_d 0.00466238f $X=2.88 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_241 N_A_79_21#_M1013_s N_A_467_47#_c_868_n 0.00304422f $X=2.745 $Y=0.235
+ $X2=0 $Y2=0
cc_242 N_A_79_21#_c_133_n N_A_467_47#_c_868_n 0.0486965f $X=2.3 $Y=0.78 $X2=0
+ $Y2=0
cc_243 N_A_79_21#_c_143_n N_A_717_47#_c_896_n 2.9459e-19 $X=4.835 $Y=1.605 $X2=0
+ $Y2=0
cc_244 N_A_79_21#_c_143_n N_A_717_47#_c_897_n 0.00468137f $X=4.835 $Y=1.605
+ $X2=0 $Y2=0
cc_245 N_C1_c_268_n N_B1_c_318_n 0.00966181f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_246 C1 B1 0.0239247f $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_247 N_C1_c_270_n B1 0.00119363f $X=2.91 $Y=1.127 $X2=0 $Y2=0
cc_248 N_C1_M1021_g N_B1_c_321_n 0.0322492f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_249 C1 N_B1_c_321_n 6.79185e-19 $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_250 N_C1_c_270_n N_B1_c_321_n 0.0145602f $X=2.91 $Y=1.127 $X2=0 $Y2=0
cc_251 N_C1_M1018_g N_VPWR_c_502_n 0.0114208f $X=2.49 $Y=1.985 $X2=0 $Y2=0
cc_252 N_C1_M1021_g N_VPWR_c_502_n 6.67793e-19 $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_253 N_C1_M1018_g N_VPWR_c_503_n 0.0046653f $X=2.49 $Y=1.985 $X2=0 $Y2=0
cc_254 N_C1_M1021_g N_VPWR_c_503_n 0.0046653f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_255 N_C1_M1018_g N_VPWR_c_504_n 6.54417e-19 $X=2.49 $Y=1.985 $X2=0 $Y2=0
cc_256 N_C1_M1021_g N_VPWR_c_504_n 0.0103686f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_257 N_C1_M1018_g N_VPWR_c_498_n 0.00796766f $X=2.49 $Y=1.985 $X2=0 $Y2=0
cc_258 N_C1_M1021_g N_VPWR_c_498_n 0.00796766f $X=2.91 $Y=1.985 $X2=0 $Y2=0
cc_259 N_C1_c_266_n N_VGND_c_745_n 0.00201943f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_260 N_C1_c_266_n N_VGND_c_754_n 0.00655123f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_261 N_C1_c_268_n N_VGND_c_754_n 0.00525237f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_262 N_C1_c_266_n N_VGND_c_756_n 0.00357877f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_263 N_C1_c_268_n N_VGND_c_756_n 0.00357877f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_264 N_C1_c_266_n N_A_467_47#_c_868_n 0.00970685f $X=2.67 $Y=0.96 $X2=0 $Y2=0
cc_265 N_C1_c_268_n N_A_467_47#_c_868_n 0.0127039f $X=3.09 $Y=0.96 $X2=0 $Y2=0
cc_266 C1 N_A_467_47#_c_868_n 9.6287e-19 $X=2.91 $Y=1.105 $X2=0 $Y2=0
cc_267 B1 A3 0.0219825f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_268 B1 N_A3_c_369_n 0.00326544f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_269 N_B1_c_321_n N_A3_c_369_n 0.00445665f $X=3.75 $Y=1.202 $X2=0 $Y2=0
cc_270 N_B1_c_322_n N_VPWR_c_504_n 0.0105091f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B1_c_323_n N_VPWR_c_504_n 6.79288e-19 $X=3.75 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_322_n N_VPWR_c_505_n 0.0046653f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_323_n N_VPWR_c_505_n 0.00585385f $X=3.75 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_323_n N_VPWR_c_506_n 0.00770434f $X=3.75 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B1_c_322_n N_VPWR_c_498_n 0.00796766f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_323_n N_VPWR_c_498_n 0.0120155f $X=3.75 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_318_n N_VGND_c_754_n 0.00525237f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B1_c_319_n N_VGND_c_754_n 0.00655123f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B1_c_318_n N_VGND_c_756_n 0.00357877f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B1_c_319_n N_VGND_c_756_n 0.00357877f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_281 B1 N_A_467_47#_c_869_n 0.011084f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_282 N_B1_c_321_n N_A_467_47#_c_869_n 5.98235e-19 $X=3.75 $Y=1.202 $X2=0 $Y2=0
cc_283 N_B1_c_318_n N_A_467_47#_c_870_n 0.0112082f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B1_c_319_n N_A_467_47#_c_870_n 0.00970685f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_285 B1 N_A_467_47#_c_870_n 0.00417723f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_286 N_B1_c_318_n N_A_717_47#_c_896_n 0.00297649f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B1_c_319_n N_A_717_47#_c_896_n 0.0120278f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_288 B1 N_A_717_47#_c_896_n 0.0630075f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_289 N_B1_c_321_n N_A_717_47#_c_896_n 0.0025555f $X=3.75 $Y=1.202 $X2=0 $Y2=0
cc_290 N_B1_c_319_n N_A_717_47#_c_897_n 0.00358764f $X=3.93 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A3_M1010_g N_A2_M1022_g 0.0190692f $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A3_c_367_n A2 2.29814e-19 $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_293 A3 A2 0.0229587f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_294 N_A3_c_367_n N_A2_c_417_n 0.0190692f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_295 A3 N_A2_c_417_n 0.00223766f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_296 N_A3_M1004_g N_VPWR_c_506_n 0.00350651f $X=4.71 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A3_M1004_g N_VPWR_c_510_n 0.00357835f $X=4.71 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A3_M1016_g N_VPWR_c_510_n 0.00357877f $X=5.13 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A3_M1004_g N_VPWR_c_498_n 0.00664109f $X=4.71 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A3_M1016_g N_VPWR_c_498_n 0.00664112f $X=5.13 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A3_M1004_g N_A_875_297#_c_660_n 0.0067463f $X=4.71 $Y=1.985 $X2=0 $Y2=0
cc_302 N_A3_M1016_g N_A_875_297#_c_660_n 5.83107e-19 $X=5.13 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A3_M1004_g N_A_875_297#_c_667_n 0.00801314f $X=4.71 $Y=1.985 $X2=0
+ $Y2=0
cc_304 N_A3_M1016_g N_A_875_297#_c_667_n 0.0162905f $X=5.13 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A3_M1004_g N_A_875_297#_c_661_n 0.00415017f $X=4.71 $Y=1.985 $X2=0
+ $Y2=0
cc_306 N_A3_c_367_n N_A_875_297#_c_662_n 0.00199437f $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_307 A3 N_A_875_297#_c_662_n 0.0226698f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_308 N_A3_c_367_n N_A_1147_297#_c_707_n 2.20109e-19 $X=5.575 $Y=1.16 $X2=0
+ $Y2=0
cc_309 A3 N_A_1147_297#_c_707_n 0.0132149f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_310 N_A3_M1010_g N_VGND_c_746_n 5.59681e-19 $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A3_M1010_g N_VGND_c_751_n 0.00343969f $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_312 N_A3_M1000_g N_VGND_c_754_n 0.00542652f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A3_M1010_g N_VGND_c_754_n 0.0040777f $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_314 N_A3_M1000_g N_VGND_c_756_n 0.00343969f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A3_M1000_g N_VGND_c_757_n 0.00998459f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A3_M1010_g N_VGND_c_757_n 0.00820756f $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_317 N_A3_M1000_g N_A_717_47#_c_908_n 0.0124313f $X=4.88 $Y=0.56 $X2=0 $Y2=0
cc_318 N_A3_M1010_g N_A_717_47#_c_908_n 0.0124313f $X=5.65 $Y=0.56 $X2=0 $Y2=0
cc_319 A3 N_A_717_47#_c_908_n 0.0664264f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_320 N_A3_c_369_n N_A_717_47#_c_908_n 0.0106396f $X=5.205 $Y=1.16 $X2=0 $Y2=0
cc_321 A3 N_A_717_47#_c_897_n 0.00776161f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_322 N_A3_c_369_n N_A_717_47#_c_897_n 0.00347805f $X=5.205 $Y=1.16 $X2=0 $Y2=0
cc_323 A3 N_A_717_47#_c_898_n 0.0060421f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_324 N_A2_M1023_g N_A1_M1001_g 0.0268753f $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A2_M1014_g N_A1_M1003_g 0.0268753f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_326 A2 A1 0.0219796f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_327 A2 N_A1_c_463_n 0.00246182f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_328 N_A2_c_417_n N_A1_c_463_n 0.0268753f $X=6.49 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A2_M1014_g N_VPWR_c_507_n 0.00220481f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A2_M1006_g N_VPWR_c_510_n 0.00357835f $X=6.07 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A2_M1014_g N_VPWR_c_510_n 0.00539841f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A2_M1006_g N_VPWR_c_498_n 0.0066022f $X=6.07 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A2_M1014_g N_VPWR_c_498_n 0.00969144f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A2_M1006_g N_A_875_297#_c_662_n 0.00403388f $X=6.07 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A2_M1006_g N_A_875_297#_c_663_n 0.0108202f $X=6.07 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A2_M1014_g N_A_875_297#_c_663_n 0.00320695f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_337 N_A2_M1006_g N_A_875_297#_c_680_n 0.00649787f $X=6.07 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A2_M1014_g N_A_875_297#_c_680_n 0.00574261f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_339 N_A2_M1006_g N_A_1147_297#_c_713_n 0.0148475f $X=6.07 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A2_M1014_g N_A_1147_297#_c_713_n 0.0156313f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_341 A2 N_A_1147_297#_c_713_n 0.0385921f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_342 N_A2_c_417_n N_A_1147_297#_c_713_n 6.177e-19 $X=6.49 $Y=1.16 $X2=0 $Y2=0
cc_343 A2 N_A_1147_297#_c_710_n 0.0128337f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A2_M1022_g N_VGND_c_746_n 0.0070524f $X=6.07 $Y=0.56 $X2=0 $Y2=0
cc_345 N_A2_M1023_g N_VGND_c_746_n 0.00706261f $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A2_M1023_g N_VGND_c_747_n 5.60103e-19 $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A2_M1022_g N_VGND_c_751_n 0.00343969f $X=6.07 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A2_M1023_g N_VGND_c_752_n 0.00343969f $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_349 N_A2_M1022_g N_VGND_c_754_n 0.00409398f $X=6.07 $Y=0.56 $X2=0 $Y2=0
cc_350 N_A2_M1023_g N_VGND_c_754_n 0.00409398f $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_351 N_A2_M1022_g N_VGND_c_757_n 5.75836e-19 $X=6.07 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A2_M1022_g N_A_717_47#_c_915_n 0.0109681f $X=6.07 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A2_M1023_g N_A_717_47#_c_915_n 0.0106382f $X=6.49 $Y=0.56 $X2=0 $Y2=0
cc_354 A2 N_A_717_47#_c_915_n 0.0371643f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_355 N_A2_c_417_n N_A_717_47#_c_915_n 0.00201657f $X=6.49 $Y=1.16 $X2=0 $Y2=0
cc_356 A2 N_A_717_47#_c_899_n 0.0128184f $X=6.59 $Y=1.105 $X2=0 $Y2=0
cc_357 N_A1_M1003_g N_VPWR_c_507_n 0.0139764f $X=6.91 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A1_M1026_g N_VPWR_c_507_n 0.0123094f $X=7.33 $Y=1.985 $X2=0 $Y2=0
cc_359 N_A1_M1003_g N_VPWR_c_510_n 0.0046653f $X=6.91 $Y=1.985 $X2=0 $Y2=0
cc_360 N_A1_M1026_g N_VPWR_c_511_n 0.0046653f $X=7.33 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A1_M1003_g N_VPWR_c_498_n 0.00799591f $X=6.91 $Y=1.985 $X2=0 $Y2=0
cc_362 N_A1_M1026_g N_VPWR_c_498_n 0.00897796f $X=7.33 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A1_M1003_g N_A_875_297#_c_663_n 4.97148e-19 $X=6.91 $Y=1.985 $X2=0
+ $Y2=0
cc_364 N_A1_M1003_g N_A_875_297#_c_680_n 5.65979e-19 $X=6.91 $Y=1.985 $X2=0
+ $Y2=0
cc_365 N_A1_M1003_g N_A_1147_297#_c_708_n 0.0172227f $X=6.91 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_A1_M1026_g N_A_1147_297#_c_708_n 0.0168728f $X=7.33 $Y=1.985 $X2=0
+ $Y2=0
cc_367 A1 N_A_1147_297#_c_708_n 0.0557881f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_368 N_A1_c_463_n N_A_1147_297#_c_708_n 0.00187137f $X=7.33 $Y=1.16 $X2=0
+ $Y2=0
cc_369 N_A1_M1001_g N_VGND_c_746_n 5.60103e-19 $X=6.91 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A1_M1001_g N_VGND_c_747_n 0.00706261f $X=6.91 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A1_M1027_g N_VGND_c_747_n 0.00878851f $X=7.33 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A1_M1001_g N_VGND_c_752_n 0.00343969f $X=6.91 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A1_M1027_g N_VGND_c_753_n 0.00343969f $X=7.33 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A1_M1001_g N_VGND_c_754_n 0.00409398f $X=6.91 $Y=0.56 $X2=0 $Y2=0
cc_375 N_A1_M1027_g N_VGND_c_754_n 0.00507603f $X=7.33 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A1_M1001_g N_A_717_47#_c_920_n 0.0122054f $X=6.91 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A1_M1027_g N_A_717_47#_c_920_n 0.0106382f $X=7.33 $Y=0.56 $X2=0 $Y2=0
cc_378 A1 N_A_717_47#_c_920_n 0.0305584f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_379 N_A1_c_463_n N_A_717_47#_c_920_n 0.00201657f $X=7.33 $Y=1.16 $X2=0 $Y2=0
cc_380 A1 N_A_717_47#_c_900_n 0.022872f $X=7.51 $Y=1.105 $X2=0 $Y2=0
cc_381 N_A1_c_463_n N_A_717_47#_c_900_n 0.00389396f $X=7.33 $Y=1.16 $X2=0 $Y2=0
cc_382 N_VPWR_c_498_n N_X_M1002_d 0.00570907f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_498_n N_X_M1020_d 0.00570907f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_508_n N_X_c_641_n 0.0113958f $X=0.935 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_498_n N_X_c_641_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_M1005_s N_X_c_618_n 0.00314561f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_387 N_VPWR_c_501_n N_X_c_618_n 0.017435f $X=1.1 $Y=2.02 $X2=0 $Y2=0
cc_388 N_VPWR_c_509_n N_X_c_645_n 0.0113958f $X=1.775 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_498_n N_X_c_645_n 0.00646998f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_500_n N_X_c_615_n 0.0260916f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_391 N_VPWR_c_498_n N_A_875_297#_M1004_d 0.00210122f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_392 N_VPWR_c_498_n N_A_875_297#_M1016_d 0.00210127f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_498_n N_A_875_297#_M1006_s 0.00215201f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_506_n N_A_875_297#_c_660_n 0.02144f $X=3.96 $Y=2.06 $X2=0 $Y2=0
cc_395 N_VPWR_c_510_n N_A_875_297#_c_667_n 0.0322563f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_498_n N_A_875_297#_c_667_n 0.0207396f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_506_n N_A_875_297#_c_661_n 0.0097139f $X=3.96 $Y=2.06 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_510_n N_A_875_297#_c_661_n 0.0209659f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_498_n N_A_875_297#_c_661_n 0.0125139f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_507_n N_A_875_297#_c_663_n 0.00551528f $X=7.12 $Y=2.02 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_510_n N_A_875_297#_c_663_n 0.0545209f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_498_n N_A_875_297#_c_663_n 0.033645f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_507_n N_A_875_297#_c_680_n 0.00518536f $X=7.12 $Y=2.02 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_510_n N_A_875_297#_c_664_n 0.0188252f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_498_n N_A_875_297#_c_664_n 0.0103982f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_498_n N_A_1147_297#_M1006_d 0.00210147f $X=7.59 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_407 N_VPWR_c_498_n N_A_1147_297#_M1014_d 0.00622412f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_498_n N_A_1147_297#_M1026_s 0.00387172f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_510_n N_A_1147_297#_c_725_n 0.0034111f $X=6.955 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_498_n N_A_1147_297#_c_725_n 0.00519041f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_M1003_d N_A_1147_297#_c_708_n 0.00315342f $X=6.985 $Y=1.485 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_507_n N_A_1147_297#_c_708_n 0.017435f $X=7.12 $Y=2.02 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_511_n N_A_1147_297#_c_709_n 0.0194349f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_498_n N_A_1147_297#_c_709_n 0.0107063f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_X_c_626_n N_VGND_M1017_d 0.00305927f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_416 N_X_c_615_n N_VGND_c_743_n 0.0260916f $X=0.595 $Y=1.185 $X2=0 $Y2=0
cc_417 N_X_c_626_n N_VGND_c_744_n 0.0163351f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_418 N_X_c_626_n N_VGND_c_748_n 0.0020257f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_419 N_X_c_616_n N_VGND_c_748_n 0.0113346f $X=1.52 $Y=0.72 $X2=0 $Y2=0
cc_420 N_X_c_626_n N_VGND_c_750_n 0.0020257f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_421 N_X_c_654_p N_VGND_c_750_n 0.0113958f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_422 N_X_M1012_s N_VGND_c_754_n 0.00417167f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_423 N_X_M1019_s N_VGND_c_754_n 0.00417167f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_424 N_X_c_626_n N_VGND_c_754_n 0.00913773f $X=1.435 $Y=0.8 $X2=0 $Y2=0
cc_425 N_X_c_654_p N_VGND_c_754_n 0.00646998f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_426 N_X_c_616_n N_VGND_c_754_n 0.00645703f $X=1.52 $Y=0.72 $X2=0 $Y2=0
cc_427 N_A_875_297#_c_663_n N_A_1147_297#_M1006_d 0.00480843f $X=6.115 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_428 N_A_875_297#_c_662_n N_A_1147_297#_c_706_n 0.0320836f $X=5.34 $Y=1.805
+ $X2=0 $Y2=0
cc_429 N_A_875_297#_c_663_n N_A_1147_297#_c_706_n 0.0184655f $X=6.115 $Y=2.38
+ $X2=0 $Y2=0
cc_430 N_A_875_297#_M1006_s N_A_1147_297#_c_713_n 0.00315342f $X=6.145 $Y=1.485
+ $X2=0 $Y2=0
cc_431 N_A_875_297#_c_663_n N_A_1147_297#_c_713_n 0.0030597f $X=6.115 $Y=2.38
+ $X2=0 $Y2=0
cc_432 N_A_875_297#_c_680_n N_A_1147_297#_c_713_n 0.0171917f $X=6.28 $Y=2.02
+ $X2=0 $Y2=0
cc_433 N_A_875_297#_c_662_n N_A_1147_297#_c_707_n 0.0209301f $X=5.34 $Y=1.805
+ $X2=0 $Y2=0
cc_434 N_A_1147_297#_c_713_n N_A_717_47#_c_915_n 6.10904e-19 $X=6.615 $Y=1.605
+ $X2=0 $Y2=0
cc_435 N_A_1147_297#_c_708_n N_A_717_47#_c_920_n 0.00285457f $X=7.455 $Y=1.605
+ $X2=0 $Y2=0
cc_436 N_A_1147_297#_c_707_n N_A_717_47#_c_898_n 0.00304105f $X=5.945 $Y=1.605
+ $X2=0 $Y2=0
cc_437 N_A_1147_297#_c_710_n N_A_717_47#_c_899_n 2.76459e-19 $X=6.7 $Y=1.605
+ $X2=0 $Y2=0
cc_438 N_VGND_c_754_n N_A_467_47#_M1013_d 0.00209344f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_439 N_VGND_c_754_n N_A_467_47#_M1015_d 0.0021521f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_754_n N_A_467_47#_M1009_d 0.00209344f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_745_n N_A_467_47#_c_868_n 0.0211533f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_442 N_VGND_c_754_n N_A_467_47#_c_868_n 0.0367981f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_756_n N_A_467_47#_c_868_n 0.0592983f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_444 N_VGND_c_754_n N_A_467_47#_c_870_n 0.0330421f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_756_n N_A_467_47#_c_870_n 0.0526799f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_446 N_VGND_c_754_n N_A_467_47#_c_890_n 0.00653405f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_756_n N_A_467_47#_c_890_n 0.0114055f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_448 N_VGND_c_754_n N_A_717_47#_M1007_s 0.00216833f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_449 N_VGND_c_754_n N_A_717_47#_M1000_d 0.00230473f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_754_n N_A_717_47#_M1010_d 0.00257509f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_754_n N_A_717_47#_M1023_d 0.00257509f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_754_n N_A_717_47#_M1027_s 0.00230473f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_754_n N_A_717_47#_c_896_n 0.00633184f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_756_n N_A_717_47#_c_896_n 0.00306647f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_455 N_VGND_M1000_s N_A_717_47#_c_908_n 0.0125147f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_VGND_c_751_n N_A_717_47#_c_908_n 0.00224243f $X=6.115 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_c_754_n N_A_717_47#_c_908_n 0.011033f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_458 N_VGND_c_756_n N_A_717_47#_c_908_n 0.00224243f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_459 N_VGND_c_757_n N_A_717_47#_c_908_n 0.0436983f $X=5.605 $Y=0.21 $X2=0
+ $Y2=0
cc_460 N_VGND_M1022_s N_A_717_47#_c_915_n 0.00307587f $X=6.145 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_VGND_c_746_n N_A_717_47#_c_915_n 0.0163829f $X=6.28 $Y=0.36 $X2=0 $Y2=0
cc_462 N_VGND_c_751_n N_A_717_47#_c_915_n 0.00224243f $X=6.115 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_c_752_n N_A_717_47#_c_915_n 0.00224243f $X=6.955 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_754_n N_A_717_47#_c_915_n 0.00960972f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_M1001_d N_A_717_47#_c_920_n 0.00307587f $X=6.985 $Y=0.235 $X2=0
+ $Y2=0
cc_466 N_VGND_c_747_n N_A_717_47#_c_920_n 0.0163829f $X=7.12 $Y=0.36 $X2=0 $Y2=0
cc_467 N_VGND_c_752_n N_A_717_47#_c_920_n 0.00224243f $X=6.955 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_753_n N_A_717_47#_c_920_n 0.00224243f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_754_n N_A_717_47#_c_920_n 0.00960972f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_754_n N_A_717_47#_c_897_n 0.0103005f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_756_n N_A_717_47#_c_897_n 0.0186139f $X=4.925 $Y=0.21 $X2=0
+ $Y2=0
cc_472 N_VGND_c_751_n N_A_717_47#_c_898_n 0.0113346f $X=6.115 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_754_n N_A_717_47#_c_898_n 0.00645703f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_752_n N_A_717_47#_c_899_n 0.0113346f $X=6.955 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_754_n N_A_717_47#_c_899_n 0.00645703f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_753_n N_A_717_47#_c_900_n 0.0193268f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_c_754_n N_A_717_47#_c_900_n 0.0106848f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_478 N_A_467_47#_c_870_n N_A_717_47#_M1007_s 0.00305418f $X=4.14 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_479 N_A_467_47#_M1009_d N_A_717_47#_c_896_n 0.00520747f $X=4.005 $Y=0.235
+ $X2=0 $Y2=0
cc_480 N_A_467_47#_c_870_n N_A_717_47#_c_896_n 0.0411983f $X=4.14 $Y=0.38 $X2=0
+ $Y2=0
cc_481 N_A_467_47#_c_870_n N_A_717_47#_c_897_n 0.0207686f $X=4.14 $Y=0.38 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__dlrbp_2.pxi.spice
* Created: Thu Aug 27 14:17:00 2020
* 
x_PM_SKY130_FD_SC_HD__DLRBP_2%GATE N_GATE_c_176_n N_GATE_c_171_n N_GATE_M1024_g
+ N_GATE_c_177_n N_GATE_M1012_g N_GATE_c_172_n N_GATE_c_178_n GATE GATE
+ N_GATE_c_174_n N_GATE_c_175_n PM_SKY130_FD_SC_HD__DLRBP_2%GATE
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1012_s
+ N_A_27_47#_M1014_g N_A_27_47#_M1000_g N_A_27_47#_M1001_g N_A_27_47#_c_215_n
+ N_A_27_47#_c_216_n N_A_27_47#_M1006_g N_A_27_47#_c_228_n N_A_27_47#_c_218_n
+ N_A_27_47#_c_219_n N_A_27_47#_c_220_n N_A_27_47#_c_229_n N_A_27_47#_c_230_n
+ N_A_27_47#_c_221_n N_A_27_47#_c_222_n N_A_27_47#_c_232_n N_A_27_47#_c_233_n
+ N_A_27_47#_c_234_n N_A_27_47#_c_235_n N_A_27_47#_c_236_n N_A_27_47#_c_237_n
+ N_A_27_47#_c_223_n PM_SKY130_FD_SC_HD__DLRBP_2%A_27_47#
x_PM_SKY130_FD_SC_HD__DLRBP_2%D N_D_M1005_g N_D_M1020_g D N_D_c_363_n
+ N_D_c_364_n PM_SKY130_FD_SC_HD__DLRBP_2%D
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_299_47# N_A_299_47#_M1005_s N_A_299_47#_M1020_s
+ N_A_299_47#_M1010_g N_A_299_47#_M1015_g N_A_299_47#_c_409_n
+ N_A_299_47#_c_402_n N_A_299_47#_c_410_n N_A_299_47#_c_411_n
+ N_A_299_47#_c_403_n N_A_299_47#_c_404_n N_A_299_47#_c_405_n
+ N_A_299_47#_c_406_n N_A_299_47#_c_407_n PM_SKY130_FD_SC_HD__DLRBP_2%A_299_47#
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_193_47# N_A_193_47#_M1014_d N_A_193_47#_M1000_d
+ N_A_193_47#_M1018_g N_A_193_47#_M1026_g N_A_193_47#_c_487_n
+ N_A_193_47#_c_488_n N_A_193_47#_c_495_n N_A_193_47#_c_489_n
+ N_A_193_47#_c_490_n N_A_193_47#_c_496_n N_A_193_47#_c_497_n
+ N_A_193_47#_c_498_n N_A_193_47#_c_499_n N_A_193_47#_c_491_n
+ N_A_193_47#_c_500_n N_A_193_47#_c_501_n PM_SKY130_FD_SC_HD__DLRBP_2%A_193_47#
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_711_307# N_A_711_307#_M1007_s
+ N_A_711_307#_M1002_d N_A_711_307#_M1013_g N_A_711_307#_M1019_g
+ N_A_711_307#_c_613_n N_A_711_307#_M1003_g N_A_711_307#_M1011_g
+ N_A_711_307#_c_614_n N_A_711_307#_M1023_g N_A_711_307#_M1027_g
+ N_A_711_307#_c_615_n N_A_711_307#_c_616_n N_A_711_307#_M1021_g
+ N_A_711_307#_M1025_g N_A_711_307#_c_618_n N_A_711_307#_c_630_n
+ N_A_711_307#_c_631_n N_A_711_307#_c_638_p N_A_711_307#_c_642_p
+ N_A_711_307#_c_657_p N_A_711_307#_c_632_n N_A_711_307#_c_619_n
+ N_A_711_307#_c_661_p N_A_711_307#_c_620_n N_A_711_307#_c_621_n
+ PM_SKY130_FD_SC_HD__DLRBP_2%A_711_307#
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_561_413# N_A_561_413#_M1018_d
+ N_A_561_413#_M1001_d N_A_561_413#_c_758_n N_A_561_413#_M1007_g
+ N_A_561_413#_M1002_g N_A_561_413#_c_759_n N_A_561_413#_c_760_n
+ N_A_561_413#_c_769_n N_A_561_413#_c_770_n N_A_561_413#_c_761_n
+ N_A_561_413#_c_767_n N_A_561_413#_c_762_n N_A_561_413#_c_763_n
+ PM_SKY130_FD_SC_HD__DLRBP_2%A_561_413#
x_PM_SKY130_FD_SC_HD__DLRBP_2%RESET_B N_RESET_B_M1016_g N_RESET_B_M1008_g
+ RESET_B N_RESET_B_c_840_n N_RESET_B_c_841_n N_RESET_B_c_842_n
+ PM_SKY130_FD_SC_HD__DLRBP_2%RESET_B
x_PM_SKY130_FD_SC_HD__DLRBP_2%A_1316_47# N_A_1316_47#_M1021_s
+ N_A_1316_47#_M1025_s N_A_1316_47#_c_877_n N_A_1316_47#_M1004_g
+ N_A_1316_47#_M1017_g N_A_1316_47#_c_878_n N_A_1316_47#_M1009_g
+ N_A_1316_47#_M1022_g N_A_1316_47#_c_881_n N_A_1316_47#_c_886_n
+ N_A_1316_47#_c_882_n N_A_1316_47#_c_896_n
+ PM_SKY130_FD_SC_HD__DLRBP_2%A_1316_47#
x_PM_SKY130_FD_SC_HD__DLRBP_2%VPWR N_VPWR_M1012_d N_VPWR_M1020_d N_VPWR_M1013_d
+ N_VPWR_M1002_s N_VPWR_M1008_d N_VPWR_M1027_d N_VPWR_M1025_d N_VPWR_M1022_d
+ N_VPWR_c_947_n N_VPWR_c_948_n N_VPWR_c_949_n N_VPWR_c_950_n N_VPWR_c_951_n
+ N_VPWR_c_952_n N_VPWR_c_953_n VPWR N_VPWR_c_954_n N_VPWR_c_955_n
+ N_VPWR_c_956_n N_VPWR_c_957_n N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n
+ N_VPWR_c_961_n N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n
+ N_VPWR_c_966_n N_VPWR_c_946_n PM_SKY130_FD_SC_HD__DLRBP_2%VPWR
x_PM_SKY130_FD_SC_HD__DLRBP_2%Q N_Q_M1003_d N_Q_M1011_s N_Q_c_1079_n
+ N_Q_c_1081_n N_Q_c_1093_n Q Q Q N_Q_c_1100_n PM_SKY130_FD_SC_HD__DLRBP_2%Q
x_PM_SKY130_FD_SC_HD__DLRBP_2%Q_N N_Q_N_M1004_d N_Q_N_M1017_s N_Q_N_c_1118_n
+ N_Q_N_c_1126_n N_Q_N_c_1128_n N_Q_N_c_1120_n N_Q_N_c_1132_n Q_N Q_N Q_N Q_N
+ Q_N PM_SKY130_FD_SC_HD__DLRBP_2%Q_N
x_PM_SKY130_FD_SC_HD__DLRBP_2%VGND N_VGND_M1024_d N_VGND_M1005_d N_VGND_M1019_d
+ N_VGND_M1016_d N_VGND_M1023_s N_VGND_M1021_d N_VGND_M1009_s N_VGND_c_1147_n
+ N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ N_VGND_c_1152_n N_VGND_c_1153_n N_VGND_c_1154_n VGND N_VGND_c_1155_n
+ N_VGND_c_1156_n N_VGND_c_1157_n N_VGND_c_1158_n N_VGND_c_1159_n
+ N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n
+ N_VGND_c_1168_n PM_SKY130_FD_SC_HD__DLRBP_2%VGND
cc_1 VNB N_GATE_c_171_n 0.0172359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_GATE_c_172_n 0.0231104f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB GATE 0.0128731f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_GATE_c_174_n 0.0212744f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_GATE_c_175_n 0.0148062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_27_47#_M1014_g 0.0397896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.135
cc_7 VNB N_A_27_47#_c_215_n 0.0133352f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_c_216_n 0.00520223f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_9 VNB N_A_27_47#_M1006_g 0.0463995f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_10 VNB N_A_27_47#_c_218_n 0.0112465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_219_n 0.00225297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_220_n 0.00793517f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_221_n 7.86136e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_222_n 0.00419087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_223_n 0.0230671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1005_g 0.025905f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_17 VNB N_D_M1020_g 0.00623929f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_18 VNB N_D_c_363_n 0.00407935f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_19 VNB N_D_c_364_n 0.0421785f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_20 VNB N_A_299_47#_M1015_g 0.0129409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_299_47#_c_402_n 0.00285527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_299_47#_c_403_n 0.00496114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_299_47#_c_404_n 0.0033094f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.235
cc_24 VNB N_A_299_47#_c_405_n 0.00265154f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_25 VNB N_A_299_47#_c_406_n 0.0274388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_299_47#_c_407_n 0.01709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_193_47#_c_487_n 0.0140955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_193_47#_c_488_n 0.00466868f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_29 VNB N_A_193_47#_c_489_n 0.0271289f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_30 VNB N_A_193_47#_c_490_n 0.00380485f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_31 VNB N_A_193_47#_c_491_n 0.0176114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_711_307#_M1019_g 0.050573f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_33 VNB N_A_711_307#_c_613_n 0.0159621f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_34 VNB N_A_711_307#_c_614_n 0.0187611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_711_307#_c_615_n 0.0472642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_711_307#_c_616_n 0.0289705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_711_307#_M1021_g 0.035711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_711_307#_c_618_n 0.00814735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_711_307#_c_619_n 0.00595002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_711_307#_c_620_n 0.00184091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_711_307#_c_621_n 0.00106791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_561_413#_c_758_n 0.0223177f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_43 VNB N_A_561_413#_c_759_n 0.042106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_561_413#_c_760_n 0.00807173f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.665
cc_45 VNB N_A_561_413#_c_761_n 0.0073863f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_46 VNB N_A_561_413#_c_762_n 0.00349711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_561_413#_c_763_n 0.0110602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_RESET_B_c_840_n 0.020032f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_49 VNB N_RESET_B_c_841_n 0.0019514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_842_n 0.0167388f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_51 VNB N_A_1316_47#_c_877_n 0.0164712f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_52 VNB N_A_1316_47#_c_878_n 0.0410818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1316_47#_M1009_g 0.0237845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1316_47#_M1022_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_55 VNB N_A_1316_47#_c_881_n 0.00889151f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_56 VNB N_A_1316_47#_c_882_n 0.0040705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_946_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_Q_c_1079_n 0.00226542f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_59 VNB N_Q_N_c_1118_n 0.00121055f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.74
cc_60 VNB Q_N 0.015424f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_61 VNB N_VGND_c_1147_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_62 VNB N_VGND_c_1148_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_63 VNB N_VGND_c_1149_n 0.00700347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1150_n 3.99405e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1151_n 0.00491053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1152_n 0.00204791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1153_n 0.00991007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1154_n 0.0315363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1155_n 0.0146858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1156_n 0.0271747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1157_n 0.0409479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1158_n 0.0276212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1159_n 0.0125407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1160_n 0.018206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1161_n 0.0153644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1162_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1163_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1164_n 0.00507544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1165_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1166_n 0.00526381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1167_n 0.00462184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1168_n 0.416824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VPB N_GATE_c_176_n 0.0128877f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.59
cc_84 VPB N_GATE_c_177_n 0.0186098f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.74
cc_85 VPB N_GATE_c_178_n 0.0238684f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_86 VPB GATE 0.0128465f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_87 VPB N_GATE_c_174_n 0.0108705f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_88 VPB N_A_27_47#_M1000_g 0.0394963f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_89 VPB N_A_27_47#_M1001_g 0.0300673f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.665
cc_90 VPB N_A_27_47#_c_215_n 0.0174193f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_91 VPB N_A_27_47#_c_216_n 0.00955572f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_92 VPB N_A_27_47#_c_228_n 0.0121288f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_93 VPB N_A_27_47#_c_229_n 0.00126297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_c_230_n 0.0300266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_221_n 6.01599e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_c_232_n 0.0224566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_27_47#_c_233_n 0.00376537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_27_47#_c_234_n 0.00546179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_47#_c_235_n 0.00344459f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_27_47#_c_236_n 0.00529835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_27_47#_c_237_n 0.00947367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_47#_c_223_n 0.0115914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_D_M1020_g 0.0462501f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_104 VPB N_D_c_363_n 0.00235013f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_105 VPB N_A_299_47#_M1015_g 0.0366983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_299_47#_c_409_n 0.00712099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_299_47#_c_410_n 0.00409088f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_108 VPB N_A_299_47#_c_411_n 0.00290124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_299_47#_c_404_n 0.00355393f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_110 VPB N_A_193_47#_M1026_g 0.0205785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_193_47#_c_487_n 0.00804665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_193_47#_c_488_n 0.00254424f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_113 VPB N_A_193_47#_c_495_n 0.00293933f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_114 VPB N_A_193_47#_c_496_n 0.00872299f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_115 VPB N_A_193_47#_c_497_n 0.00238602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_193_47#_c_498_n 0.00711634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_193_47#_c_499_n 0.00237469f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_193_47#_c_500_n 0.0267112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_193_47#_c_501_n 0.00795904f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_711_307#_M1013_g 0.0291104f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_121 VPB N_A_711_307#_M1019_g 0.0183333f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_122 VPB N_A_711_307#_M1011_g 0.0183857f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_123 VPB N_A_711_307#_M1027_g 0.0225684f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_124 VPB N_A_711_307#_c_615_n 0.0230116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_711_307#_c_616_n 0.00603343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_711_307#_M1025_g 0.0474712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_711_307#_c_618_n 5.1591e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_711_307#_c_630_n 0.00523696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_711_307#_c_631_n 0.04731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_711_307#_c_632_n 0.00155778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_561_413#_M1002_g 0.0255039f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_561_413#_c_759_n 0.0151075f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_561_413#_c_760_n 5.1126e-19 $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.665
cc_134 VPB N_A_561_413#_c_767_n 0.00880061f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_135 VPB N_A_561_413#_c_762_n 0.00182699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_M1008_g 0.0195094f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_137 VPB N_RESET_B_c_840_n 0.00406721f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_138 VPB N_RESET_B_c_841_n 0.00209991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_1316_47#_M1017_g 0.0191443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_1316_47#_c_878_n 0.00447364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_1316_47#_M1022_g 0.0264718f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_142 VPB N_A_1316_47#_c_886_n 0.0129935f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_143 VPB N_A_1316_47#_c_882_n 0.0044458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_947_n 0.00126149f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_145 VPB N_VPWR_c_948_n 0.00343394f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_146 VPB N_VPWR_c_949_n 3.18587e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_950_n 0.0111729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_951_n 0.00288228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_952_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_953_n 0.0425526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_954_n 0.0146514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_955_n 0.0295132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_956_n 0.0125756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_957_n 0.0158421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_958_n 0.0184742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_959_n 0.0153644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_960_n 0.00473435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_961_n 0.00440565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_962_n 0.0387638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_963_n 0.0281605f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_964_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_965_n 0.00497181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_966_n 0.00443372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_946_n 0.0598897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_Q_c_1079_n 0.00325141f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_166 VPB N_Q_c_1081_n 0.00338591f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.135
cc_167 VPB N_Q_N_c_1120_n 0.00148895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB Q_N 0.00509247f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_169 N_GATE_c_171_n N_A_27_47#_M1014_g 0.0187834f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_170 N_GATE_c_175_n N_A_27_47#_M1014_g 0.0041981f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_171 N_GATE_c_178_n N_A_27_47#_M1000_g 0.0260359f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_172 N_GATE_c_174_n N_A_27_47#_M1000_g 0.00527228f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_173 N_GATE_c_171_n N_A_27_47#_c_219_n 0.00674622f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_174 N_GATE_c_172_n N_A_27_47#_c_219_n 0.0105293f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_175 N_GATE_c_172_n N_A_27_47#_c_220_n 0.00672951f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_176 GATE N_A_27_47#_c_220_n 0.0202563f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_177 N_GATE_c_174_n N_A_27_47#_c_220_n 7.62625e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_178 N_GATE_c_177_n N_A_27_47#_c_229_n 0.0135762f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_179 N_GATE_c_178_n N_A_27_47#_c_229_n 0.00220936f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_180 N_GATE_c_177_n N_A_27_47#_c_230_n 2.2048e-19 $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_181 N_GATE_c_178_n N_A_27_47#_c_230_n 0.00396f $X=0.47 $Y=1.665 $X2=0 $Y2=0
cc_182 GATE N_A_27_47#_c_230_n 0.0221922f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_183 N_GATE_c_174_n N_A_27_47#_c_230_n 5.90345e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_184 N_GATE_c_174_n N_A_27_47#_c_221_n 0.00319708f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_185 N_GATE_c_172_n N_A_27_47#_c_222_n 0.00179331f $X=0.47 $Y=0.805 $X2=0
+ $Y2=0
cc_186 GATE N_A_27_47#_c_222_n 0.0288709f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_187 N_GATE_c_175_n N_A_27_47#_c_222_n 0.0015185f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_188 N_GATE_c_176_n N_A_27_47#_c_233_n 0.0033897f $X=0.305 $Y=1.59 $X2=0 $Y2=0
cc_189 N_GATE_c_178_n N_A_27_47#_c_233_n 0.00102562f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_190 GATE N_A_27_47#_c_233_n 0.00653918f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_191 N_GATE_c_176_n N_A_27_47#_c_234_n 7.60515e-19 $X=0.305 $Y=1.59 $X2=0
+ $Y2=0
cc_192 N_GATE_c_178_n N_A_27_47#_c_234_n 0.00427582f $X=0.47 $Y=1.665 $X2=0
+ $Y2=0
cc_193 GATE N_A_27_47#_c_223_n 9.06759e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_194 N_GATE_c_174_n N_A_27_47#_c_223_n 0.0165992f $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_195 N_GATE_c_177_n N_VPWR_c_947_n 0.00946555f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_196 N_GATE_c_177_n N_VPWR_c_954_n 0.00332278f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_197 N_GATE_c_177_n N_VPWR_c_946_n 0.00484884f $X=0.47 $Y=1.74 $X2=0 $Y2=0
cc_198 N_GATE_c_171_n N_VGND_c_1147_n 0.0112612f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_199 N_GATE_c_171_n N_VGND_c_1155_n 0.00339367f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_200 N_GATE_c_172_n N_VGND_c_1155_n 4.74473e-19 $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_201 N_GATE_c_171_n N_VGND_c_1168_n 0.00497794f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_232_n N_D_M1020_g 0.00583826f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_232_n N_D_c_363_n 0.0087134f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_204 N_A_27_47#_M1014_g N_D_c_364_n 0.00520956f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A_27_47#_M1001_g N_A_299_47#_M1015_g 0.0353942f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_216_n N_A_299_47#_M1015_g 0.0248435f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_232_n N_A_299_47#_M1015_g 0.00493352f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_235_n N_A_299_47#_M1015_g 0.00140912f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_236_n N_A_299_47#_M1015_g 0.00239179f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_232_n N_A_299_47#_c_410_n 0.0116439f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_211 N_A_27_47#_c_235_n N_A_299_47#_c_410_n 0.00130924f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_236_n N_A_299_47#_c_410_n 0.00675603f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_232_n N_A_299_47#_c_411_n 0.0115067f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_232_n N_A_299_47#_c_403_n 0.00675641f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_232_n N_A_299_47#_c_404_n 0.0108494f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_c_235_n N_A_299_47#_c_404_n 0.00124596f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_236_n N_A_299_47#_c_404_n 0.00570493f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_232_n N_A_299_47#_c_406_n 0.00107604f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_M1001_g N_A_193_47#_M1026_g 0.019647f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1014_g N_A_193_47#_c_487_n 0.00779983f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_219_n N_A_193_47#_c_487_n 0.0100297f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_c_221_n N_A_193_47#_c_487_n 0.023541f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_222_n N_A_193_47#_c_487_n 0.0158341f $X=0.725 $Y=1.07 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_232_n N_A_193_47#_c_487_n 0.0184539f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_233_n N_A_193_47#_c_487_n 0.00230203f $X=0.84 $Y=1.53 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_234_n N_A_193_47#_c_487_n 0.0208179f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_215_n N_A_193_47#_c_488_n 0.0127601f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_228 N_A_27_47#_M1006_g N_A_193_47#_c_488_n 0.00492704f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_235_n N_A_193_47#_c_488_n 0.00101104f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_236_n N_A_193_47#_c_488_n 0.0151027f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_237_n N_A_193_47#_c_488_n 0.00406305f $X=2.67 $Y=1.52 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_229_n N_A_193_47#_c_495_n 0.00294892f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_232_n N_A_193_47#_c_495_n 0.00195186f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_223_n N_A_193_47#_c_495_n 0.00779983f $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_216_n N_A_193_47#_c_489_n 0.0188813f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1006_g N_A_193_47#_c_489_n 0.0192792f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_236_n N_A_193_47#_c_489_n 4.13927e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_215_n N_A_193_47#_c_490_n 7.03475e-19 $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_216_n N_A_193_47#_c_490_n 0.00136198f $X=2.805 $Y=1.32 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1006_g N_A_193_47#_c_490_n 0.00256371f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_c_236_n N_A_193_47#_c_490_n 0.00180905f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_M1001_g N_A_193_47#_c_496_n 0.00736818f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_215_n N_A_193_47#_c_496_n 0.00118095f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_228_n N_A_193_47#_c_496_n 0.00185018f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_232_n N_A_193_47#_c_496_n 0.0871075f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_235_n N_A_193_47#_c_496_n 0.0266068f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_236_n N_A_193_47#_c_496_n 0.00864674f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1000_g N_A_193_47#_c_497_n 0.00458322f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_229_n N_A_193_47#_c_497_n 0.00551586f $X=0.61 $Y=1.88 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_232_n N_A_193_47#_c_497_n 0.0259095f $X=2.41 $Y=1.53 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_234_n N_A_193_47#_c_497_n 0.00110517f $X=0.695 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1000_g N_A_193_47#_c_498_n 0.00779983f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_M1001_g N_A_193_47#_c_499_n 0.00145116f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_215_n N_A_193_47#_c_499_n 0.00113693f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1006_g N_A_193_47#_c_491_n 0.0126141f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_215_n N_A_193_47#_c_500_n 0.0184363f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_228_n N_A_193_47#_c_500_n 0.0166555f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_215_n N_A_193_47#_c_501_n 0.00399682f $X=3.145 $Y=1.32 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_228_n N_A_193_47#_c_501_n 0.00596961f $X=2.67 $Y=1.685 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_235_n N_A_193_47#_c_501_n 4.76211e-19 $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_236_n N_A_193_47#_c_501_n 0.00815409f $X=2.555 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1006_g N_A_711_307#_M1019_g 0.0425869f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1001_g N_A_561_413#_c_769_n 0.0049672f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1006_g N_A_561_413#_c_770_n 0.0125275f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1006_g N_A_561_413#_c_761_n 0.00562201f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_c_215_n N_A_561_413#_c_767_n 6.99098e-19 $X=3.145 $Y=1.32
+ $X2=0 $Y2=0
cc_267 N_A_27_47#_M1006_g N_A_561_413#_c_763_n 0.00352817f $X=3.22 $Y=0.415
+ $X2=0 $Y2=0
cc_268 N_A_27_47#_c_229_n N_VPWR_M1012_d 0.00193227f $X=0.61 $Y=1.88 $X2=-0.19
+ $Y2=-0.24
cc_269 N_A_27_47#_M1000_g N_VPWR_c_947_n 0.00964955f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_229_n N_VPWR_c_947_n 0.015089f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_230_n N_VPWR_c_947_n 0.0127436f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_233_n N_VPWR_c_947_n 0.0031008f $X=0.84 $Y=1.53 $X2=0 $Y2=0
cc_273 N_A_27_47#_M1001_g N_VPWR_c_948_n 0.00401328f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_232_n N_VPWR_c_948_n 0.0019389f $X=2.41 $Y=1.53 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_229_n N_VPWR_c_954_n 0.0018545f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_230_n N_VPWR_c_954_n 0.0184766f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_277 N_A_27_47#_M1000_g N_VPWR_c_955_n 0.00442511f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1001_g N_VPWR_c_962_n 0.00497675f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1000_g N_VPWR_c_946_n 0.00889084f $X=0.89 $Y=2.135 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_M1001_g N_VPWR_c_946_n 0.00611433f $X=2.73 $Y=2.275 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_229_n N_VPWR_c_946_n 0.00483676f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_230_n N_VPWR_c_946_n 0.00993215f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_219_n N_VGND_M1024_d 0.00166538f $X=0.61 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_284 N_A_27_47#_M1014_g N_VGND_c_1147_n 0.011777f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_219_n N_VGND_c_1147_n 0.0150802f $X=0.61 $Y=0.72 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_221_n N_VGND_c_1147_n 0.00124842f $X=0.755 $Y=1.235 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_223_n N_VGND_c_1147_n 5.79361e-19 $X=0.89 $Y=1.235 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1006_g N_VGND_c_1149_n 0.0017297f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_218_n N_VGND_c_1155_n 0.0110793f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_219_n N_VGND_c_1155_n 0.00243651f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1014_g N_VGND_c_1156_n 0.0046653f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_M1006_g N_VGND_c_1157_n 0.0037981f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1024_s N_VGND_c_1168_n 0.00234409f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1014_g N_VGND_c_1168_n 0.00934473f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1006_g N_VGND_c_1168_n 0.00555936f $X=3.22 $Y=0.415 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_218_n N_VGND_c_1168_n 0.00934849f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_219_n N_VGND_c_1168_n 0.00549708f $X=0.61 $Y=0.72 $X2=0
+ $Y2=0
cc_298 N_D_c_364_n N_A_299_47#_M1015_g 0.03863f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_299 N_D_M1020_g N_A_299_47#_c_409_n 0.012851f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_300 N_D_M1005_g N_A_299_47#_c_402_n 0.0144498f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_301 N_D_c_363_n N_A_299_47#_c_402_n 0.00627239f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_302 N_D_c_364_n N_A_299_47#_c_402_n 0.00123166f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_303 N_D_M1020_g N_A_299_47#_c_410_n 0.00794545f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_304 N_D_M1020_g N_A_299_47#_c_411_n 0.00412429f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_305 N_D_c_363_n N_A_299_47#_c_411_n 0.0229667f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_306 N_D_c_364_n N_A_299_47#_c_411_n 0.00131849f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_307 N_D_M1005_g N_A_299_47#_c_403_n 0.00563568f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_308 N_D_c_363_n N_A_299_47#_c_403_n 0.0107593f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_309 N_D_c_363_n N_A_299_47#_c_404_n 0.0164827f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_310 N_D_c_364_n N_A_299_47#_c_404_n 0.00552652f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_311 N_D_M1005_g N_A_299_47#_c_405_n 0.00120855f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_312 N_D_c_363_n N_A_299_47#_c_405_n 0.0138491f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_313 N_D_c_364_n N_A_299_47#_c_405_n 0.0042466f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_314 N_D_M1005_g N_A_299_47#_c_406_n 0.0197208f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_315 N_D_M1005_g N_A_299_47#_c_407_n 0.015283f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_316 N_D_M1005_g N_A_193_47#_c_487_n 0.00203374f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_317 N_D_M1020_g N_A_193_47#_c_487_n 0.00459933f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_318 N_D_c_363_n N_A_193_47#_c_487_n 0.0209974f $X=1.625 $Y=1.04 $X2=0 $Y2=0
cc_319 N_D_c_364_n N_A_193_47#_c_487_n 0.00256393f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_320 N_D_M1020_g N_A_193_47#_c_495_n 0.00134564f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_321 N_D_M1020_g N_A_193_47#_c_496_n 0.00294239f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_322 N_D_M1020_g N_VPWR_c_948_n 0.00304701f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_323 N_D_M1020_g N_VPWR_c_955_n 0.00543342f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_324 N_D_M1020_g N_VPWR_c_946_n 0.00734866f $X=1.83 $Y=2.165 $X2=0 $Y2=0
cc_325 N_D_M1005_g N_VGND_c_1148_n 0.0110406f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_326 N_D_M1005_g N_VGND_c_1156_n 0.00337001f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_327 N_D_M1005_g N_VGND_c_1168_n 0.0053254f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_328 N_D_c_364_n N_VGND_c_1168_n 0.00103829f $X=1.83 $Y=1.04 $X2=0 $Y2=0
cc_329 N_A_299_47#_c_409_n N_A_193_47#_c_487_n 0.0010921f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_330 N_A_299_47#_c_411_n N_A_193_47#_c_487_n 0.00859001f $X=1.785 $Y=1.58
+ $X2=0 $Y2=0
cc_331 N_A_299_47#_c_405_n N_A_193_47#_c_487_n 0.0191833f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_332 N_A_299_47#_M1015_g N_A_193_47#_c_488_n 0.00370009f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_333 N_A_299_47#_c_403_n N_A_193_47#_c_488_n 0.00178567f $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_334 N_A_299_47#_c_406_n N_A_193_47#_c_488_n 9.9633e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_335 N_A_299_47#_c_409_n N_A_193_47#_c_495_n 0.0471072f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_336 N_A_299_47#_c_403_n N_A_193_47#_c_489_n 9.56555e-19 $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_337 N_A_299_47#_c_406_n N_A_193_47#_c_489_n 0.0117556f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_338 N_A_299_47#_c_407_n N_A_193_47#_c_489_n 0.00200147f $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_339 N_A_299_47#_c_403_n N_A_193_47#_c_490_n 0.0129081f $X=2.055 $Y=1.095
+ $X2=0 $Y2=0
cc_340 N_A_299_47#_c_406_n N_A_193_47#_c_490_n 9.50608e-19 $X=2.255 $Y=0.93
+ $X2=0 $Y2=0
cc_341 N_A_299_47#_c_407_n N_A_193_47#_c_490_n 2.04855e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_342 N_A_299_47#_M1015_g N_A_193_47#_c_496_n 0.00365242f $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_343 N_A_299_47#_c_409_n N_A_193_47#_c_496_n 0.022748f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_344 N_A_299_47#_c_410_n N_A_193_47#_c_496_n 0.00551435f $X=1.97 $Y=1.58 $X2=0
+ $Y2=0
cc_345 N_A_299_47#_c_409_n N_A_193_47#_c_497_n 0.00273055f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_346 N_A_299_47#_c_407_n N_A_193_47#_c_491_n 0.0197019f $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_347 N_A_299_47#_M1015_g N_A_561_413#_c_769_n 5.24267e-19 $X=2.25 $Y=2.165
+ $X2=0 $Y2=0
cc_348 N_A_299_47#_c_407_n N_A_561_413#_c_770_n 7.34833e-19 $X=2.255 $Y=0.765
+ $X2=0 $Y2=0
cc_349 N_A_299_47#_M1015_g N_VPWR_c_948_n 0.0234057f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_350 N_A_299_47#_c_409_n N_VPWR_c_948_n 0.0232987f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_351 N_A_299_47#_c_410_n N_VPWR_c_948_n 0.013562f $X=1.97 $Y=1.58 $X2=0 $Y2=0
cc_352 N_A_299_47#_c_409_n N_VPWR_c_955_n 0.0159418f $X=1.62 $Y=1.99 $X2=0 $Y2=0
cc_353 N_A_299_47#_M1015_g N_VPWR_c_962_n 0.00212864f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_354 N_A_299_47#_M1020_s N_VPWR_c_946_n 0.00174533f $X=1.495 $Y=1.845 $X2=0
+ $Y2=0
cc_355 N_A_299_47#_M1015_g N_VPWR_c_946_n 0.00262666f $X=2.25 $Y=2.165 $X2=0
+ $Y2=0
cc_356 N_A_299_47#_c_409_n N_VPWR_c_946_n 0.00576627f $X=1.62 $Y=1.99 $X2=0
+ $Y2=0
cc_357 N_A_299_47#_c_403_n N_VGND_M1005_d 0.00156939f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_358 N_A_299_47#_c_402_n N_VGND_c_1148_n 0.00259081f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_359 N_A_299_47#_c_403_n N_VGND_c_1148_n 0.0141976f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_A_299_47#_c_407_n N_VGND_c_1148_n 0.00955875f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_361 N_A_299_47#_c_402_n N_VGND_c_1156_n 0.00255672f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_362 N_A_299_47#_c_405_n N_VGND_c_1156_n 0.00711582f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_363 N_A_299_47#_c_406_n N_VGND_c_1157_n 9.84895e-19 $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_364 N_A_299_47#_c_407_n N_VGND_c_1157_n 0.0046653f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_365 N_A_299_47#_M1005_s N_VGND_c_1168_n 0.00283248f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_A_299_47#_c_402_n N_VGND_c_1168_n 0.00473142f $X=1.97 $Y=0.7 $X2=0
+ $Y2=0
cc_367 N_A_299_47#_c_403_n N_VGND_c_1168_n 0.00552372f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_368 N_A_299_47#_c_405_n N_VGND_c_1168_n 0.00607883f $X=1.62 $Y=0.51 $X2=0
+ $Y2=0
cc_369 N_A_299_47#_c_406_n N_VGND_c_1168_n 0.00117722f $X=2.255 $Y=0.93 $X2=0
+ $Y2=0
cc_370 N_A_299_47#_c_407_n N_VGND_c_1168_n 0.00454932f $X=2.255 $Y=0.765 $X2=0
+ $Y2=0
cc_371 N_A_193_47#_M1026_g N_A_711_307#_M1013_g 0.0263455f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_372 N_A_193_47#_c_501_n N_A_711_307#_M1013_g 2.14526e-19 $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_373 N_A_193_47#_c_500_n N_A_711_307#_c_631_n 0.0167148f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_374 N_A_193_47#_c_501_n N_A_711_307#_c_631_n 3.98623e-19 $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_375 N_A_193_47#_M1026_g N_A_561_413#_c_769_n 0.00895296f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_376 N_A_193_47#_c_496_n N_A_561_413#_c_769_n 0.00281719f $X=2.87 $Y=1.87
+ $X2=0 $Y2=0
cc_377 N_A_193_47#_c_499_n N_A_561_413#_c_769_n 0.00272719f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_378 N_A_193_47#_c_501_n N_A_561_413#_c_769_n 0.0119883f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_379 N_A_193_47#_c_489_n N_A_561_413#_c_770_n 0.00144439f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_380 N_A_193_47#_c_490_n N_A_561_413#_c_770_n 0.021036f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_381 N_A_193_47#_c_491_n N_A_561_413#_c_770_n 0.00674639f $X=2.8 $Y=0.705
+ $X2=0 $Y2=0
cc_382 N_A_193_47#_c_490_n N_A_561_413#_c_761_n 0.0184898f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_383 N_A_193_47#_M1026_g N_A_561_413#_c_767_n 0.00377053f $X=3.15 $Y=2.275
+ $X2=0 $Y2=0
cc_384 N_A_193_47#_c_488_n N_A_561_413#_c_767_n 0.0113318f $X=3.01 $Y=1.575
+ $X2=0 $Y2=0
cc_385 N_A_193_47#_c_499_n N_A_561_413#_c_767_n 0.00286078f $X=3.015 $Y=1.87
+ $X2=0 $Y2=0
cc_386 N_A_193_47#_c_500_n N_A_561_413#_c_767_n 0.00425391f $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_387 N_A_193_47#_c_501_n N_A_561_413#_c_767_n 0.02751f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_388 N_A_193_47#_c_488_n N_A_561_413#_c_763_n 0.0167533f $X=3.01 $Y=1.575
+ $X2=0 $Y2=0
cc_389 N_A_193_47#_c_490_n N_A_561_413#_c_763_n 0.0027819f $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_390 N_A_193_47#_c_500_n N_A_561_413#_c_763_n 4.91178e-19 $X=3.18 $Y=1.74
+ $X2=0 $Y2=0
cc_391 N_A_193_47#_c_496_n N_VPWR_M1020_d 6.81311e-19 $X=2.87 $Y=1.87 $X2=0
+ $Y2=0
cc_392 N_A_193_47#_c_498_n N_VPWR_c_947_n 0.0127357f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_393 N_A_193_47#_c_496_n N_VPWR_c_948_n 0.0184713f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_394 N_A_193_47#_c_499_n N_VPWR_c_948_n 9.60597e-19 $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_395 N_A_193_47#_c_501_n N_VPWR_c_948_n 0.00216895f $X=3.18 $Y=1.74 $X2=0
+ $Y2=0
cc_396 N_A_193_47#_c_498_n N_VPWR_c_955_n 0.015988f $X=1.155 $Y=1.87 $X2=0 $Y2=0
cc_397 N_A_193_47#_M1026_g N_VPWR_c_962_n 0.00366111f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_398 N_A_193_47#_M1026_g N_VPWR_c_946_n 0.00538229f $X=3.15 $Y=2.275 $X2=0
+ $Y2=0
cc_399 N_A_193_47#_c_496_n N_VPWR_c_946_n 0.0750488f $X=2.87 $Y=1.87 $X2=0 $Y2=0
cc_400 N_A_193_47#_c_497_n N_VPWR_c_946_n 0.0151526f $X=1.3 $Y=1.87 $X2=0 $Y2=0
cc_401 N_A_193_47#_c_498_n N_VPWR_c_946_n 0.00389918f $X=1.155 $Y=1.87 $X2=0
+ $Y2=0
cc_402 N_A_193_47#_c_499_n N_VPWR_c_946_n 0.0148792f $X=3.015 $Y=1.87 $X2=0
+ $Y2=0
cc_403 N_A_193_47#_c_496_n A_465_369# 0.00388705f $X=2.87 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_404 N_A_193_47#_c_491_n N_VGND_c_1148_n 0.0017371f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_405 N_A_193_47#_c_487_n N_VGND_c_1156_n 0.00732874f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_406 N_A_193_47#_c_489_n N_VGND_c_1157_n 9.43262e-19 $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_407 N_A_193_47#_c_490_n N_VGND_c_1157_n 8.03214e-19 $X=3.01 $Y=0.87 $X2=0
+ $Y2=0
cc_408 N_A_193_47#_c_491_n N_VGND_c_1157_n 0.00400086f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_409 N_A_193_47#_M1014_d N_VGND_c_1168_n 0.00535012f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_410 N_A_193_47#_c_487_n N_VGND_c_1168_n 0.00616598f $X=1.1 $Y=0.51 $X2=0
+ $Y2=0
cc_411 N_A_193_47#_c_489_n N_VGND_c_1168_n 0.00121904f $X=2.8 $Y=0.87 $X2=0
+ $Y2=0
cc_412 N_A_193_47#_c_490_n N_VGND_c_1168_n 0.00182f $X=3.01 $Y=0.87 $X2=0 $Y2=0
cc_413 N_A_193_47#_c_491_n N_VGND_c_1168_n 0.0059606f $X=2.8 $Y=0.705 $X2=0
+ $Y2=0
cc_414 N_A_711_307#_c_638_p N_A_561_413#_c_758_n 0.00990518f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_415 N_A_711_307#_c_619_n N_A_561_413#_c_758_n 0.00595161f $X=4.425 $Y=0.58
+ $X2=0 $Y2=0
cc_416 N_A_711_307#_c_630_n N_A_561_413#_M1002_g 0.0166068f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_417 N_A_711_307#_c_631_n N_A_561_413#_M1002_g 0.0064088f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_418 N_A_711_307#_c_642_p N_A_561_413#_M1002_g 0.00661649f $X=4.855 $Y=2.27
+ $X2=0 $Y2=0
cc_419 N_A_711_307#_M1019_g N_A_561_413#_c_759_n 0.0214321f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_420 N_A_711_307#_c_630_n N_A_561_413#_c_759_n 0.0145126f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_421 N_A_711_307#_c_631_n N_A_561_413#_c_759_n 0.00487525f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_422 N_A_711_307#_c_619_n N_A_561_413#_c_759_n 0.00885226f $X=4.425 $Y=0.58
+ $X2=0 $Y2=0
cc_423 N_A_711_307#_M1019_g N_A_561_413#_c_770_n 0.00160594f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_424 N_A_711_307#_M1019_g N_A_561_413#_c_761_n 0.010318f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_425 N_A_711_307#_M1013_g N_A_561_413#_c_767_n 0.0213969f $X=3.63 $Y=2.275
+ $X2=0 $Y2=0
cc_426 N_A_711_307#_M1019_g N_A_561_413#_c_767_n 0.00744096f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_427 N_A_711_307#_c_630_n N_A_561_413#_c_767_n 0.0192637f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_428 N_A_711_307#_c_631_n N_A_561_413#_c_767_n 0.0103945f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_429 N_A_711_307#_M1019_g N_A_561_413#_c_762_n 0.0244229f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_430 N_A_711_307#_c_630_n N_A_561_413#_c_762_n 0.02399f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_431 N_A_711_307#_c_631_n N_A_561_413#_c_762_n 0.00672107f $X=3.925 $Y=1.7
+ $X2=0 $Y2=0
cc_432 N_A_711_307#_M1011_g N_RESET_B_M1008_g 0.0227734f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_A_711_307#_c_657_p N_RESET_B_M1008_g 0.0128217f $X=5.32 $Y=1.62 $X2=0
+ $Y2=0
cc_434 N_A_711_307#_c_632_n N_RESET_B_M1008_g 0.00443134f $X=5.415 $Y=1.535
+ $X2=0 $Y2=0
cc_435 N_A_711_307#_c_616_n N_RESET_B_c_840_n 0.0203089f $X=6.05 $Y=1.16 $X2=0
+ $Y2=0
cc_436 N_A_711_307#_c_638_p N_RESET_B_c_840_n 0.00144439f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_437 N_A_711_307#_c_661_p N_RESET_B_c_840_n 4.32398e-19 $X=4.855 $Y=1.755
+ $X2=0 $Y2=0
cc_438 N_A_711_307#_c_620_n N_RESET_B_c_840_n 0.00197689f $X=5.535 $Y=1.16 $X2=0
+ $Y2=0
cc_439 N_A_711_307#_c_616_n N_RESET_B_c_841_n 3.21195e-19 $X=6.05 $Y=1.16 $X2=0
+ $Y2=0
cc_440 N_A_711_307#_c_630_n N_RESET_B_c_841_n 0.0202313f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_441 N_A_711_307#_c_638_p N_RESET_B_c_841_n 0.0384833f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_711_307#_c_657_p N_RESET_B_c_841_n 0.0109472f $X=5.32 $Y=1.62 $X2=0
+ $Y2=0
cc_443 N_A_711_307#_c_619_n N_RESET_B_c_841_n 0.0109732f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_444 N_A_711_307#_c_661_p N_RESET_B_c_841_n 0.012291f $X=4.855 $Y=1.755 $X2=0
+ $Y2=0
cc_445 N_A_711_307#_c_620_n N_RESET_B_c_841_n 0.0273265f $X=5.535 $Y=1.16 $X2=0
+ $Y2=0
cc_446 N_A_711_307#_c_613_n N_RESET_B_c_842_n 0.0211574f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A_711_307#_c_638_p N_RESET_B_c_842_n 0.0117784f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_711_307#_c_619_n N_RESET_B_c_842_n 0.00108664f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_449 N_A_711_307#_c_621_n N_RESET_B_c_842_n 0.00357987f $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_450 N_A_711_307#_M1021_g N_A_1316_47#_c_877_n 0.0197646f $X=6.915 $Y=0.445
+ $X2=0 $Y2=0
cc_451 N_A_711_307#_M1025_g N_A_1316_47#_M1017_g 0.0225541f $X=6.915 $Y=2.165
+ $X2=0 $Y2=0
cc_452 N_A_711_307#_c_618_n N_A_1316_47#_c_878_n 0.0209606f $X=6.915 $Y=1.16
+ $X2=0 $Y2=0
cc_453 N_A_711_307#_c_614_n N_A_1316_47#_c_881_n 0.00559975f $X=5.975 $Y=0.995
+ $X2=0 $Y2=0
cc_454 N_A_711_307#_M1021_g N_A_1316_47#_c_881_n 0.019901f $X=6.915 $Y=0.445
+ $X2=0 $Y2=0
cc_455 N_A_711_307#_M1027_g N_A_1316_47#_c_886_n 0.0054592f $X=5.975 $Y=1.985
+ $X2=0 $Y2=0
cc_456 N_A_711_307#_M1025_g N_A_1316_47#_c_886_n 0.0273964f $X=6.915 $Y=2.165
+ $X2=0 $Y2=0
cc_457 N_A_711_307#_c_618_n N_A_1316_47#_c_882_n 0.0181222f $X=6.915 $Y=1.16
+ $X2=0 $Y2=0
cc_458 N_A_711_307#_c_615_n N_A_1316_47#_c_896_n 0.0248708f $X=6.84 $Y=1.16
+ $X2=0 $Y2=0
cc_459 N_A_711_307#_c_618_n N_A_1316_47#_c_896_n 0.0011918f $X=6.915 $Y=1.16
+ $X2=0 $Y2=0
cc_460 N_A_711_307#_c_630_n N_VPWR_M1002_s 0.00639144f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_461 N_A_711_307#_c_657_p N_VPWR_M1008_d 0.00685929f $X=5.32 $Y=1.62 $X2=0
+ $Y2=0
cc_462 N_A_711_307#_c_632_n N_VPWR_M1008_d 5.79934e-19 $X=5.415 $Y=1.535 $X2=0
+ $Y2=0
cc_463 N_A_711_307#_M1011_g N_VPWR_c_949_n 0.0113184f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_464 N_A_711_307#_M1027_g N_VPWR_c_949_n 4.79945e-19 $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_465 N_A_711_307#_c_657_p N_VPWR_c_949_n 0.0219885f $X=5.32 $Y=1.62 $X2=0
+ $Y2=0
cc_466 N_A_711_307#_M1027_g N_VPWR_c_950_n 0.00314703f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_467 N_A_711_307#_c_615_n N_VPWR_c_950_n 0.00146061f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_468 N_A_711_307#_M1025_g N_VPWR_c_950_n 0.00326926f $X=6.915 $Y=2.165 $X2=0
+ $Y2=0
cc_469 N_A_711_307#_M1025_g N_VPWR_c_951_n 0.00297479f $X=6.915 $Y=2.165 $X2=0
+ $Y2=0
cc_470 N_A_711_307#_c_642_p N_VPWR_c_956_n 0.00972841f $X=4.855 $Y=2.27 $X2=0
+ $Y2=0
cc_471 N_A_711_307#_M1011_g N_VPWR_c_957_n 0.0046653f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_472 N_A_711_307#_M1027_g N_VPWR_c_957_n 0.00541359f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_A_711_307#_M1025_g N_VPWR_c_958_n 0.00541359f $X=6.915 $Y=2.165 $X2=0
+ $Y2=0
cc_474 N_A_711_307#_M1013_g N_VPWR_c_962_n 0.00520872f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_475 N_A_711_307#_M1013_g N_VPWR_c_963_n 0.00483063f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_476 N_A_711_307#_c_630_n N_VPWR_c_963_n 0.039758f $X=4.77 $Y=1.7 $X2=0 $Y2=0
cc_477 N_A_711_307#_c_631_n N_VPWR_c_963_n 0.00809172f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_478 N_A_711_307#_c_642_p N_VPWR_c_963_n 0.0235008f $X=4.855 $Y=2.27 $X2=0
+ $Y2=0
cc_479 N_A_711_307#_M1002_d N_VPWR_c_946_n 0.00443507f $X=4.71 $Y=1.485 $X2=0
+ $Y2=0
cc_480 N_A_711_307#_M1013_g N_VPWR_c_946_n 0.0103589f $X=3.63 $Y=2.275 $X2=0
+ $Y2=0
cc_481 N_A_711_307#_M1011_g N_VPWR_c_946_n 0.00794405f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_482 N_A_711_307#_M1027_g N_VPWR_c_946_n 0.0108799f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_483 N_A_711_307#_M1025_g N_VPWR_c_946_n 0.0109968f $X=6.915 $Y=2.165 $X2=0
+ $Y2=0
cc_484 N_A_711_307#_c_630_n N_VPWR_c_946_n 0.00825301f $X=4.77 $Y=1.7 $X2=0
+ $Y2=0
cc_485 N_A_711_307#_c_631_n N_VPWR_c_946_n 0.00123717f $X=3.925 $Y=1.7 $X2=0
+ $Y2=0
cc_486 N_A_711_307#_c_642_p N_VPWR_c_946_n 0.00637538f $X=4.855 $Y=2.27 $X2=0
+ $Y2=0
cc_487 N_A_711_307#_c_613_n N_Q_c_1079_n 0.00205731f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_A_711_307#_c_614_n N_Q_c_1079_n 0.0152777f $X=5.975 $Y=0.995 $X2=0
+ $Y2=0
cc_489 N_A_711_307#_c_615_n N_Q_c_1079_n 0.0223633f $X=6.84 $Y=1.16 $X2=0 $Y2=0
cc_490 N_A_711_307#_c_616_n N_Q_c_1079_n 0.0162799f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_491 N_A_711_307#_M1021_g N_Q_c_1079_n 0.00133246f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_492 N_A_711_307#_c_638_p N_Q_c_1079_n 0.0136f $X=5.32 $Y=0.74 $X2=0 $Y2=0
cc_493 N_A_711_307#_c_620_n N_Q_c_1079_n 0.0257936f $X=5.535 $Y=1.16 $X2=0 $Y2=0
cc_494 N_A_711_307#_c_621_n N_Q_c_1079_n 0.0093605f $X=5.47 $Y=0.995 $X2=0 $Y2=0
cc_495 N_A_711_307#_M1011_g N_Q_c_1081_n 0.00120596f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_496 N_A_711_307#_M1027_g N_Q_c_1081_n 0.00584713f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_497 N_A_711_307#_c_632_n N_Q_c_1081_n 0.00870075f $X=5.415 $Y=1.535 $X2=0
+ $Y2=0
cc_498 N_A_711_307#_M1011_g N_Q_c_1093_n 0.00731262f $X=5.535 $Y=1.985 $X2=0
+ $Y2=0
cc_499 N_A_711_307#_M1027_g N_Q_c_1093_n 0.0124021f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_500 N_A_711_307#_c_616_n N_Q_c_1093_n 0.0027047f $X=6.05 $Y=1.16 $X2=0 $Y2=0
cc_501 N_A_711_307#_c_657_p N_Q_c_1093_n 0.0140134f $X=5.32 $Y=1.62 $X2=0 $Y2=0
cc_502 N_A_711_307#_c_632_n N_Q_c_1093_n 0.00298593f $X=5.415 $Y=1.535 $X2=0
+ $Y2=0
cc_503 N_A_711_307#_c_613_n Q 0.0040044f $X=5.535 $Y=0.995 $X2=0 $Y2=0
cc_504 N_A_711_307#_c_638_p Q 7.49507e-19 $X=5.32 $Y=0.74 $X2=0 $Y2=0
cc_505 N_A_711_307#_M1027_g N_Q_c_1100_n 0.0118052f $X=5.975 $Y=1.985 $X2=0
+ $Y2=0
cc_506 N_A_711_307#_c_638_p N_VGND_M1016_d 0.00679393f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_711_307#_c_621_n N_VGND_M1016_d 6.98288e-19 $X=5.47 $Y=0.995 $X2=0
+ $Y2=0
cc_508 N_A_711_307#_M1019_g N_VGND_c_1149_n 0.0115145f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_711_307#_c_619_n N_VGND_c_1149_n 0.0084822f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_510 N_A_711_307#_c_613_n N_VGND_c_1150_n 0.00771894f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_511 N_A_711_307#_c_614_n N_VGND_c_1150_n 7.60567e-19 $X=5.975 $Y=0.995 $X2=0
+ $Y2=0
cc_512 N_A_711_307#_c_638_p N_VGND_c_1150_n 0.0207574f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_711_307#_c_619_n N_VGND_c_1150_n 0.00204313f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_514 N_A_711_307#_c_613_n N_VGND_c_1151_n 7.4812e-19 $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_515 N_A_711_307#_c_614_n N_VGND_c_1151_n 0.00840969f $X=5.975 $Y=0.995 $X2=0
+ $Y2=0
cc_516 N_A_711_307#_c_615_n N_VGND_c_1151_n 0.00119981f $X=6.84 $Y=1.16 $X2=0
+ $Y2=0
cc_517 N_A_711_307#_M1021_g N_VGND_c_1151_n 0.00215585f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_518 N_A_711_307#_M1021_g N_VGND_c_1152_n 0.00164839f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_519 N_A_711_307#_M1019_g N_VGND_c_1157_n 0.0046653f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_520 N_A_711_307#_c_638_p N_VGND_c_1158_n 0.0078938f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_711_307#_c_619_n N_VGND_c_1158_n 0.00903426f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_522 N_A_711_307#_c_613_n N_VGND_c_1159_n 0.00446579f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_523 N_A_711_307#_c_614_n N_VGND_c_1159_n 0.0034272f $X=5.975 $Y=0.995 $X2=0
+ $Y2=0
cc_524 N_A_711_307#_c_638_p N_VGND_c_1159_n 3.34073e-19 $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_711_307#_M1021_g N_VGND_c_1160_n 0.0054895f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_526 N_A_711_307#_M1007_s N_VGND_c_1168_n 0.00233038f $X=4.3 $Y=0.235 $X2=0
+ $Y2=0
cc_527 N_A_711_307#_M1019_g N_VGND_c_1168_n 0.00813035f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_528 N_A_711_307#_c_613_n N_VGND_c_1168_n 0.00733753f $X=5.535 $Y=0.995 $X2=0
+ $Y2=0
cc_529 N_A_711_307#_c_614_n N_VGND_c_1168_n 0.00409821f $X=5.975 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_711_307#_M1021_g N_VGND_c_1168_n 0.0112465f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_531 N_A_711_307#_c_638_p N_VGND_c_1168_n 0.0160201f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_532 N_A_711_307#_c_619_n N_VGND_c_1168_n 0.0102202f $X=4.425 $Y=0.58 $X2=0
+ $Y2=0
cc_533 N_A_711_307#_c_638_p A_942_47# 0.00470094f $X=5.32 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_534 N_A_561_413#_M1002_g N_RESET_B_M1008_g 0.0228015f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_535 N_A_561_413#_c_760_n N_RESET_B_c_840_n 0.0214965f $X=4.635 $Y=1.16 $X2=0
+ $Y2=0
cc_536 N_A_561_413#_c_759_n N_RESET_B_c_841_n 0.0115911f $X=4.56 $Y=1.16 $X2=0
+ $Y2=0
cc_537 N_A_561_413#_c_760_n N_RESET_B_c_841_n 0.012104f $X=4.635 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_A_561_413#_c_762_n N_RESET_B_c_841_n 0.0243426f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_539 N_A_561_413#_c_758_n N_RESET_B_c_842_n 0.0410517f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_561_413#_c_769_n N_VPWR_c_948_n 0.00578043f $X=3.27 $Y=2.34 $X2=0
+ $Y2=0
cc_541 N_A_561_413#_M1002_g N_VPWR_c_949_n 6.67854e-19 $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_542 N_A_561_413#_M1002_g N_VPWR_c_956_n 0.00427505f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_543 N_A_561_413#_c_769_n N_VPWR_c_962_n 0.0226583f $X=3.27 $Y=2.34 $X2=0
+ $Y2=0
cc_544 N_A_561_413#_c_767_n N_VPWR_c_962_n 0.0156263f $X=3.52 $Y=1.96 $X2=0
+ $Y2=0
cc_545 N_A_561_413#_M1002_g N_VPWR_c_963_n 0.0108273f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_546 N_A_561_413#_M1001_d N_VPWR_c_946_n 0.00173835f $X=2.805 $Y=2.065 $X2=0
+ $Y2=0
cc_547 N_A_561_413#_M1002_g N_VPWR_c_946_n 0.00413985f $X=4.635 $Y=1.985 $X2=0
+ $Y2=0
cc_548 N_A_561_413#_c_769_n N_VPWR_c_946_n 0.00997071f $X=3.27 $Y=2.34 $X2=0
+ $Y2=0
cc_549 N_A_561_413#_c_767_n N_VPWR_c_946_n 0.0121128f $X=3.52 $Y=1.96 $X2=0
+ $Y2=0
cc_550 N_A_561_413#_c_767_n A_645_413# 0.0058803f $X=3.52 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_551 N_A_561_413#_c_770_n N_VGND_c_1148_n 0.00233934f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_552 N_A_561_413#_c_758_n N_VGND_c_1149_n 0.00644915f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_553 N_A_561_413#_c_759_n N_VGND_c_1149_n 0.00169847f $X=4.56 $Y=1.16 $X2=0
+ $Y2=0
cc_554 N_A_561_413#_c_770_n N_VGND_c_1149_n 0.0104492f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_555 N_A_561_413#_c_762_n N_VGND_c_1149_n 0.0119873f $X=4.115 $Y=1.16 $X2=0
+ $Y2=0
cc_556 N_A_561_413#_c_758_n N_VGND_c_1150_n 0.00213078f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_557 N_A_561_413#_c_770_n N_VGND_c_1157_n 0.0246608f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_558 N_A_561_413#_c_758_n N_VGND_c_1158_n 0.00426723f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_559 N_A_561_413#_M1018_d N_VGND_c_1168_n 0.00237979f $X=2.865 $Y=0.235 $X2=0
+ $Y2=0
cc_560 N_A_561_413#_c_758_n N_VGND_c_1168_n 0.00731201f $X=4.635 $Y=0.995 $X2=0
+ $Y2=0
cc_561 N_A_561_413#_c_770_n N_VGND_c_1168_n 0.0243863f $X=3.33 $Y=0.45 $X2=0
+ $Y2=0
cc_562 N_A_561_413#_c_770_n A_659_47# 0.00373396f $X=3.33 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_563 N_A_561_413#_c_761_n A_659_47# 0.00149829f $X=3.415 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_564 N_RESET_B_M1008_g N_VPWR_c_949_n 0.0110144f $X=5.065 $Y=1.985 $X2=0 $Y2=0
cc_565 N_RESET_B_M1008_g N_VPWR_c_956_n 0.0046653f $X=5.065 $Y=1.985 $X2=0 $Y2=0
cc_566 N_RESET_B_M1008_g N_VPWR_c_963_n 6.22549e-19 $X=5.065 $Y=1.985 $X2=0
+ $Y2=0
cc_567 N_RESET_B_M1008_g N_VPWR_c_946_n 0.00802136f $X=5.065 $Y=1.985 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_842_n N_VGND_c_1150_n 0.0101341f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_842_n N_VGND_c_1158_n 0.00341689f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_570 N_RESET_B_c_842_n N_VGND_c_1168_n 0.0040799f $X=5.055 $Y=0.995 $X2=0
+ $Y2=0
cc_571 N_A_1316_47#_c_886_n N_VPWR_c_950_n 0.0509455f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_572 N_A_1316_47#_M1017_g N_VPWR_c_951_n 0.0110571f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_573 N_A_1316_47#_c_878_n N_VPWR_c_951_n 0.00179383f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_574 N_A_1316_47#_M1022_g N_VPWR_c_951_n 7.50638e-19 $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_575 N_A_1316_47#_c_886_n N_VPWR_c_951_n 0.0235095f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_576 N_A_1316_47#_c_882_n N_VPWR_c_951_n 0.00978589f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_577 N_A_1316_47#_M1022_g N_VPWR_c_953_n 0.00312874f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_578 N_A_1316_47#_c_886_n N_VPWR_c_958_n 0.0213966f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_579 N_A_1316_47#_M1017_g N_VPWR_c_959_n 0.00486043f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_580 N_A_1316_47#_M1022_g N_VPWR_c_959_n 0.00541359f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_581 N_A_1316_47#_M1025_s N_VPWR_c_946_n 0.00209319f $X=6.58 $Y=1.845 $X2=0
+ $Y2=0
cc_582 N_A_1316_47#_M1017_g N_VPWR_c_946_n 0.0082748f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_583 N_A_1316_47#_M1022_g N_VPWR_c_946_n 0.0104946f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_584 N_A_1316_47#_c_886_n N_VPWR_c_946_n 0.0126193f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_585 N_A_1316_47#_c_881_n N_Q_c_1079_n 0.01964f $X=6.705 $Y=0.51 $X2=0 $Y2=0
cc_586 N_A_1316_47#_c_896_n N_Q_c_1079_n 0.0269233f $X=6.702 $Y=1.16 $X2=0 $Y2=0
cc_587 N_A_1316_47#_c_886_n N_Q_c_1081_n 0.0100636f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_588 N_A_1316_47#_c_886_n N_Q_c_1100_n 0.005053f $X=6.705 $Y=2 $X2=0 $Y2=0
cc_589 N_A_1316_47#_c_877_n N_Q_N_c_1118_n 0.00385723f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_590 N_A_1316_47#_c_878_n N_Q_N_c_1118_n 0.00314449f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_591 N_A_1316_47#_M1009_g N_Q_N_c_1118_n 0.00768995f $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_592 N_A_1316_47#_c_882_n N_Q_N_c_1118_n 0.00456865f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_593 N_A_1316_47#_c_878_n N_Q_N_c_1126_n 0.00163737f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_594 N_A_1316_47#_M1009_g N_Q_N_c_1126_n 0.00199113f $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_595 N_A_1316_47#_c_878_n N_Q_N_c_1128_n 0.00149964f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_596 N_A_1316_47#_M1022_g N_Q_N_c_1128_n 0.00155059f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_597 N_A_1316_47#_M1017_g N_Q_N_c_1120_n 0.00601018f $X=7.39 $Y=1.985 $X2=0
+ $Y2=0
cc_598 N_A_1316_47#_M1022_g N_Q_N_c_1120_n 0.0100205f $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_599 N_A_1316_47#_c_878_n N_Q_N_c_1132_n 0.00862745f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_600 N_A_1316_47#_M1022_g N_Q_N_c_1132_n 2.76149e-19 $X=7.81 $Y=1.985 $X2=0
+ $Y2=0
cc_601 N_A_1316_47#_c_882_n N_Q_N_c_1132_n 0.0226854f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_602 N_A_1316_47#_M1009_g Q_N 0.00609939f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_603 N_A_1316_47#_M1022_g Q_N 0.00928793f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_604 N_A_1316_47#_c_878_n Q_N 0.0130776f $X=7.81 $Y=1.025 $X2=0 $Y2=0
cc_605 N_A_1316_47#_M1022_g Q_N 0.00643425f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_606 N_A_1316_47#_c_881_n N_VGND_c_1151_n 0.0171711f $X=6.705 $Y=0.51 $X2=0
+ $Y2=0
cc_607 N_A_1316_47#_c_877_n N_VGND_c_1152_n 0.00756765f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_608 N_A_1316_47#_c_878_n N_VGND_c_1152_n 0.00188342f $X=7.81 $Y=1.025 $X2=0
+ $Y2=0
cc_609 N_A_1316_47#_M1009_g N_VGND_c_1152_n 6.49537e-19 $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_610 N_A_1316_47#_c_882_n N_VGND_c_1152_n 0.0108724f $X=7.34 $Y=1.16 $X2=0
+ $Y2=0
cc_611 N_A_1316_47#_M1009_g N_VGND_c_1154_n 0.00312874f $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_612 N_A_1316_47#_c_881_n N_VGND_c_1160_n 0.0210884f $X=6.705 $Y=0.51 $X2=0
+ $Y2=0
cc_613 N_A_1316_47#_c_877_n N_VGND_c_1161_n 0.00486043f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_614 N_A_1316_47#_M1009_g N_VGND_c_1161_n 0.00541359f $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_615 N_A_1316_47#_M1021_s N_VGND_c_1168_n 0.00210122f $X=6.58 $Y=0.235 $X2=0
+ $Y2=0
cc_616 N_A_1316_47#_c_877_n N_VGND_c_1168_n 0.0082748f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_617 N_A_1316_47#_M1009_g N_VGND_c_1168_n 0.0104946f $X=7.81 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_1316_47#_c_881_n N_VGND_c_1168_n 0.0125221f $X=6.705 $Y=0.51 $X2=0
+ $Y2=0
cc_619 N_VPWR_c_946_n A_465_369# 0.00476473f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_620 N_VPWR_c_946_n A_645_413# 0.00267862f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_621 N_VPWR_c_946_n N_Q_M1011_s 0.00474271f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_622 N_VPWR_c_950_n N_Q_c_1079_n 0.00936314f $X=6.185 $Y=2 $X2=0 $Y2=0
cc_623 N_VPWR_c_949_n N_Q_c_1100_n 0.0415928f $X=5.275 $Y=2.02 $X2=0 $Y2=0
cc_624 N_VPWR_c_957_n N_Q_c_1100_n 0.0153589f $X=6.1 $Y=2.72 $X2=0 $Y2=0
cc_625 N_VPWR_c_946_n N_Q_c_1100_n 0.00934584f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_626 N_VPWR_c_946_n N_Q_N_M1017_s 0.00393857f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_627 N_VPWR_c_959_n Q_N 0.0151826f $X=7.935 $Y=2.72 $X2=0 $Y2=0
cc_628 N_VPWR_c_946_n Q_N 0.00941829f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_629 N_VPWR_c_953_n Q_N 0.021861f $X=8.02 $Y=1.66 $X2=0 $Y2=0
cc_630 N_Q_c_1079_n N_VGND_M1023_s 0.00645199f $X=5.927 $Y=1.325 $X2=0 $Y2=0
cc_631 Q N_VGND_c_1150_n 0.0106188f $X=5.68 $Y=0.425 $X2=0 $Y2=0
cc_632 N_Q_c_1079_n N_VGND_c_1151_n 0.0144491f $X=5.927 $Y=1.325 $X2=0 $Y2=0
cc_633 N_Q_c_1079_n N_VGND_c_1159_n 0.00245167f $X=5.927 $Y=1.325 $X2=0 $Y2=0
cc_634 Q N_VGND_c_1159_n 0.00770732f $X=5.68 $Y=0.425 $X2=0 $Y2=0
cc_635 N_Q_M1003_d N_VGND_c_1168_n 0.00502936f $X=5.61 $Y=0.235 $X2=0 $Y2=0
cc_636 N_Q_c_1079_n N_VGND_c_1168_n 0.00506428f $X=5.927 $Y=1.325 $X2=0 $Y2=0
cc_637 Q N_VGND_c_1168_n 0.00618204f $X=5.68 $Y=0.425 $X2=0 $Y2=0
cc_638 Q_N N_VGND_c_1154_n 0.021861f $X=7.995 $Y=1.105 $X2=0 $Y2=0
cc_639 Q_N N_VGND_c_1161_n 0.0151169f $X=7.535 $Y=0.425 $X2=0 $Y2=0
cc_640 N_Q_N_M1004_d N_VGND_c_1168_n 0.00393857f $X=7.465 $Y=0.235 $X2=0 $Y2=0
cc_641 Q_N N_VGND_c_1168_n 0.00940437f $X=7.535 $Y=0.425 $X2=0 $Y2=0
cc_642 N_VGND_c_1168_n A_465_47# 0.0139156f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_643 N_VGND_c_1168_n A_659_47# 0.00687059f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24
cc_644 N_VGND_c_1168_n A_942_47# 0.00335103f $X=8.05 $Y=0 $X2=-0.19 $Y2=-0.24

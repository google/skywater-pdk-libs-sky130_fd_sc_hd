* File: sky130_fd_sc_hd__o21ba_4.spice
* Created: Thu Aug 27 14:36:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ba_4.pex.spice"
.subckt sky130_fd_sc_hd__o21ba_4  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_B1_N_M1020_g N_A_27_297#_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.19825 PD=0.92 PS=1.91 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1020_d N_A_187_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_187_21#_M1011_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1011_d N_A_187_21#_M1015_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_187_21#_M1021_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_575_47#_M1012_d N_A_27_297#_M1012_g N_A_187_21#_M1012_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1016 N_A_575_47#_M1016_d N_A_27_297#_M1016_g N_A_187_21#_M1012_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_575_47#_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1010_d N_A2_M1017_g N_A_575_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A1_M1013_g N_A_575_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1013_d N_A1_M1014_g N_A_575_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_27_297#_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.38 PD=1.27 PS=2.76 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75000.3
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1005_d N_A_187_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A_187_21#_M1007_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.1
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1007_d N_A_187_21#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1018_d N_A_187_21#_M1018_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1018_d N_A_27_297#_M1000_g N_A_187_21#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A_27_297#_M1002_g N_A_187_21#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_743_297#_M1001_d N_A2_M1001_g N_A_187_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_A_743_297#_M1004_d N_A2_M1004_g N_A_187_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1009 N_A_743_297#_M1004_d N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1019 N_A_743_297#_M1019_d N_A1_M1019_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_53 VNB 0 1.12295e-19 $X=0.145 $Y=-0.085
*
.include "sky130_fd_sc_hd__o21ba_4.pxi.spice"
*
.ends
*
*

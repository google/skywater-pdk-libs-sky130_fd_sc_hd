* File: sky130_fd_sc_hd__einvn_2.spice.SKY130_FD_SC_HD__EINVN_2.pxi
* Created: Thu Aug 27 14:20:15 2020
* 
x_PM_SKY130_FD_SC_HD__EINVN_2%TE_B N_TE_B_M1008_g N_TE_B_c_61_n N_TE_B_M1006_g
+ N_TE_B_c_65_n N_TE_B_c_66_n N_TE_B_M1002_g N_TE_B_c_67_n N_TE_B_c_68_n
+ N_TE_B_M1004_g N_TE_B_c_69_n TE_B PM_SKY130_FD_SC_HD__EINVN_2%TE_B
x_PM_SKY130_FD_SC_HD__EINVN_2%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_102_n N_A_27_47#_M1003_g N_A_27_47#_c_103_n N_A_27_47#_c_104_n
+ N_A_27_47#_c_105_n N_A_27_47#_M1005_g N_A_27_47#_c_106_n N_A_27_47#_c_111_n
+ N_A_27_47#_c_107_n N_A_27_47#_c_108_n N_A_27_47#_c_109_n N_A_27_47#_c_110_n
+ PM_SKY130_FD_SC_HD__EINVN_2%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVN_2%A N_A_M1007_g N_A_M1000_g N_A_M1009_g N_A_M1001_g
+ N_A_c_169_n A N_A_c_171_n PM_SKY130_FD_SC_HD__EINVN_2%A
x_PM_SKY130_FD_SC_HD__EINVN_2%VPWR N_VPWR_M1006_d N_VPWR_M1004_d N_VPWR_c_214_n
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n VPWR N_VPWR_c_218_n
+ N_VPWR_c_219_n N_VPWR_c_213_n N_VPWR_c_221_n N_VPWR_c_222_n
+ PM_SKY130_FD_SC_HD__EINVN_2%VPWR
x_PM_SKY130_FD_SC_HD__EINVN_2%A_204_309# N_A_204_309#_M1002_s
+ N_A_204_309#_M1000_s N_A_204_309#_c_277_n N_A_204_309#_c_262_n
+ N_A_204_309#_c_282_n N_A_204_309#_c_263_n
+ PM_SKY130_FD_SC_HD__EINVN_2%A_204_309#
x_PM_SKY130_FD_SC_HD__EINVN_2%Z N_Z_M1007_s N_Z_M1000_d N_Z_M1001_d Z Z Z Z Z Z
+ Z N_Z_c_296_n Z PM_SKY130_FD_SC_HD__EINVN_2%Z
x_PM_SKY130_FD_SC_HD__EINVN_2%VGND N_VGND_M1008_d N_VGND_M1003_s N_VGND_c_332_n
+ N_VGND_c_333_n VGND N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n
+ N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n PM_SKY130_FD_SC_HD__EINVN_2%VGND
x_PM_SKY130_FD_SC_HD__EINVN_2%A_214_120# N_A_214_120#_M1003_d
+ N_A_214_120#_M1005_d N_A_214_120#_M1009_d N_A_214_120#_c_382_n
+ N_A_214_120#_c_378_n N_A_214_120#_c_408_n N_A_214_120#_c_379_n
+ N_A_214_120#_c_380_n PM_SKY130_FD_SC_HD__EINVN_2%A_214_120#
cc_1 VNB N_TE_B_M1008_g 0.0429947f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_B_c_61_n 0.0401369f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.47
cc_3 VNB TE_B 0.0133203f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_c_102_n 0.017541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_5 VNB N_A_27_47#_c_103_n 0.0118932f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.395
cc_6 VNB N_A_27_47#_c_104_n 0.00902397f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.47
cc_7 VNB N_A_27_47#_c_105_n 0.0147779f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_8 VNB N_A_27_47#_c_106_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_9 VNB N_A_27_47#_c_107_n 0.00110654f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_10 VNB N_A_27_47#_c_108_n 0.0183891f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.395
cc_11 VNB N_A_27_47#_c_109_n 0.0186942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_110_n 0.034244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_M1007_g 0.0179476f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_14 VNB N_A_M1000_g 6.82813e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_15 VNB N_A_M1009_g 0.0235444f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.47
cc_16 VNB N_A_c_169_n 0.0267194f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_17 VNB A 0.0078301f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_A_c_171_n 0.0276634f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_19 VNB N_VPWR_c_213_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB Z 0.00141716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_332_n 0.00475141f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.395
cc_22 VNB N_VGND_c_333_n 4.11703e-19 $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=2.015
cc_23 VNB N_VGND_c_334_n 0.0143218f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_24 VNB N_VGND_c_335_n 0.0149333f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_25 VNB N_VGND_c_336_n 0.0347876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_337_n 0.188074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_338_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_339_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_214_120#_c_378_n 0.00772857f $X=-0.19 $Y=-0.24 $X2=1.365 $Y2=2.015
cc_30 VNB N_A_214_120#_c_379_n 0.0139808f $X=-0.19 $Y=-0.24 $X2=0.325 $Y2=1.16
cc_31 VNB N_A_214_120#_c_380_n 0.00702719f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.395
cc_32 VPB N_TE_B_c_61_n 0.0184868f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.47
cc_33 VPB N_TE_B_M1006_g 0.0367521f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_34 VPB N_TE_B_c_65_n 0.0185273f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.395
cc_35 VPB N_TE_B_c_66_n 0.0141524f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.47
cc_36 VPB N_TE_B_c_67_n 0.0260828f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_37 VPB N_TE_B_c_68_n 0.016581f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.47
cc_38 VPB N_TE_B_c_69_n 0.00618823f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.395
cc_39 VPB TE_B 0.0054315f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_40 VPB N_A_27_47#_c_111_n 0.03055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_107_n 0.0140666f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_42 VPB N_A_M1000_g 0.0252558f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_43 VPB N_A_M1001_g 0.026587f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.395
cc_44 VPB N_A_c_171_n 0.00701784f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_45 VPB N_VPWR_c_214_n 3.9647e-19 $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.395
cc_46 VPB N_VPWR_c_215_n 0.0130026f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.47
cc_47 VPB N_VPWR_c_216_n 0.00455076f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=2.015
cc_48 VPB N_VPWR_c_217_n 0.0118766f $X=-0.19 $Y=1.305 $X2=1.365 $Y2=1.47
cc_49 VPB N_VPWR_c_218_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.395
cc_50 VPB N_VPWR_c_219_n 0.0254149f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_213_n 0.0436139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_221_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_222_n 0.0046501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_204_309#_c_262_n 0.00597804f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=1.47
cc_55 VPB N_A_204_309#_c_263_n 0.00976501f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_56 VPB Z 0.0141095f $X=-0.19 $Y=1.305 $X2=1.29 $Y2=1.395
cc_57 VPB Z 0.0311552f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.395
cc_58 VPB N_Z_c_296_n 0.00723959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB Z 0.00195684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_TE_B_c_67_n N_A_27_47#_c_104_n 0.00721886f $X=1.29 $Y=1.395 $X2=0 $Y2=0
cc_61 N_TE_B_M1006_g N_A_27_47#_c_111_n 0.00933515f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_62 N_TE_B_c_61_n N_A_27_47#_c_107_n 0.0103412f $X=0.47 $Y=1.47 $X2=0 $Y2=0
cc_63 N_TE_B_M1006_g N_A_27_47#_c_107_n 0.023602f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_64 N_TE_B_c_65_n N_A_27_47#_c_107_n 0.015458f $X=0.87 $Y=1.395 $X2=0 $Y2=0
cc_65 N_TE_B_c_66_n N_A_27_47#_c_107_n 0.00647698f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_66 N_TE_B_c_69_n N_A_27_47#_c_107_n 0.00701012f $X=0.945 $Y=1.395 $X2=0 $Y2=0
cc_67 TE_B N_A_27_47#_c_107_n 0.0275866f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_68 N_TE_B_M1008_g N_A_27_47#_c_108_n 0.0280377f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_69 N_TE_B_c_61_n N_A_27_47#_c_108_n 0.016812f $X=0.47 $Y=1.47 $X2=0 $Y2=0
cc_70 TE_B N_A_27_47#_c_108_n 0.042038f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_TE_B_c_69_n N_A_27_47#_c_109_n 0.0168237f $X=0.945 $Y=1.395 $X2=0 $Y2=0
cc_72 N_TE_B_M1006_g N_VPWR_c_214_n 0.0125686f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_73 N_TE_B_c_66_n N_VPWR_c_214_n 0.010303f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_74 N_TE_B_c_68_n N_VPWR_c_214_n 6.0115e-19 $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_75 N_TE_B_c_66_n N_VPWR_c_216_n 5.67858e-19 $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_76 N_TE_B_c_68_n N_VPWR_c_216_n 0.00831127f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_77 N_TE_B_c_66_n N_VPWR_c_217_n 0.00486043f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_78 N_TE_B_c_68_n N_VPWR_c_217_n 0.00339367f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_79 N_TE_B_M1006_g N_VPWR_c_218_n 0.0046653f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_80 N_TE_B_M1006_g N_VPWR_c_213_n 0.00895857f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_81 N_TE_B_c_66_n N_VPWR_c_213_n 0.0082748f $X=0.945 $Y=1.47 $X2=0 $Y2=0
cc_82 N_TE_B_c_68_n N_VPWR_c_213_n 0.00397141f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_83 N_TE_B_c_66_n N_A_204_309#_c_263_n 0.00136389f $X=0.945 $Y=1.47 $X2=0
+ $Y2=0
cc_84 N_TE_B_c_67_n N_A_204_309#_c_263_n 0.00684228f $X=1.29 $Y=1.395 $X2=0
+ $Y2=0
cc_85 N_TE_B_c_68_n N_A_204_309#_c_263_n 0.0274422f $X=1.365 $Y=1.47 $X2=0 $Y2=0
cc_86 N_TE_B_c_67_n N_Z_c_296_n 9.7292e-19 $X=1.29 $Y=1.395 $X2=0 $Y2=0
cc_87 N_TE_B_M1008_g N_VGND_c_332_n 0.00966829f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_88 N_TE_B_M1008_g N_VGND_c_334_n 0.00341574f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_89 N_TE_B_M1008_g N_VGND_c_337_n 0.00501514f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_90 N_TE_B_M1008_g N_A_214_120#_c_380_n 0.00250093f $X=0.47 $Y=0.445 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_c_105_n N_A_M1007_g 0.0186064f $X=1.825 $Y=0.96 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_109_n N_A_M1007_g 2.53393e-19 $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_109_n N_A_c_169_n 0.00108159f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_110_n N_A_c_169_n 0.0181805f $X=1.87 $Y=1.035 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_107_n N_VPWR_M1006_d 0.00310745f $X=0.695 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_27_47#_c_107_n N_VPWR_c_214_n 0.0232987f $X=0.695 $Y=1.555 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_111_n N_VPWR_c_218_n 0.018001f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1006_s N_VPWR_c_213_n 0.00387172f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_111_n N_VPWR_c_213_n 0.00993603f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_109_n N_A_204_309#_c_262_n 0.00501044f $X=1.87 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_110_n N_A_204_309#_c_262_n 0.00324962f $X=1.87 $Y=1.035
+ $X2=0 $Y2=0
cc_102 N_A_27_47#_c_104_n N_A_204_309#_c_263_n 0.00147672f $X=1.48 $Y=1.035
+ $X2=0 $Y2=0
cc_103 N_A_27_47#_c_107_n N_A_204_309#_c_263_n 0.00848719f $X=0.695 $Y=1.555
+ $X2=0 $Y2=0
cc_104 N_A_27_47#_c_109_n N_A_204_309#_c_263_n 0.0590727f $X=1.87 $Y=1.16 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_110_n N_A_204_309#_c_263_n 0.0019454f $X=1.87 $Y=1.035 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_105_n Z 4.96653e-19 $X=1.825 $Y=0.96 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_109_n N_Z_c_296_n 0.00688424f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_110_n N_Z_c_296_n 0.00200161f $X=1.87 $Y=1.035 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_109_n Z 0.0128722f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_110_n Z 8.2894e-19 $X=1.87 $Y=1.035 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_108_n N_VGND_M1008_d 0.002671f $X=0.895 $Y=1.135 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_27_47#_c_102_n N_VGND_c_332_n 0.00197049f $X=1.405 $Y=0.96 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_108_n N_VGND_c_332_n 0.0249115f $X=0.895 $Y=1.135 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_102_n N_VGND_c_333_n 0.00723954f $X=1.405 $Y=0.96 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_105_n N_VGND_c_333_n 0.00808417f $X=1.825 $Y=0.96 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_106_n N_VGND_c_334_n 0.0177719f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_108_n N_VGND_c_334_n 0.00273425f $X=0.895 $Y=1.135 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_102_n N_VGND_c_335_n 0.00341689f $X=1.405 $Y=0.96 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_105_n N_VGND_c_336_n 0.00341689f $X=1.825 $Y=0.96 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_M1008_s N_VGND_c_337_n 0.00228937f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_102_n N_VGND_c_337_n 0.00540327f $X=1.405 $Y=0.96 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_105_n N_VGND_c_337_n 0.00423453f $X=1.825 $Y=0.96 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_106_n N_VGND_c_337_n 0.00989054f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_108_n N_VGND_c_337_n 0.00577733f $X=0.895 $Y=1.135 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_102_n N_A_214_120#_c_382_n 0.00940897f $X=1.405 $Y=0.96
+ $X2=0 $Y2=0
cc_126 N_A_27_47#_c_103_n N_A_214_120#_c_382_n 0.00179137f $X=1.705 $Y=1.035
+ $X2=0 $Y2=0
cc_127 N_A_27_47#_c_105_n N_A_214_120#_c_382_n 0.0103011f $X=1.825 $Y=0.96 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_c_109_n N_A_214_120#_c_382_n 0.0475193f $X=1.87 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_110_n N_A_214_120#_c_382_n 5.90934e-19 $X=1.87 $Y=1.035
+ $X2=0 $Y2=0
cc_130 N_A_27_47#_c_108_n N_A_214_120#_c_380_n 0.0156017f $X=0.895 $Y=1.135
+ $X2=0 $Y2=0
cc_131 N_A_27_47#_c_109_n N_A_214_120#_c_380_n 0.0221828f $X=1.87 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_M1000_g N_VPWR_c_219_n 0.00339367f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1001_g N_VPWR_c_219_n 0.00541359f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1000_g N_VPWR_c_213_n 0.00397141f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1001_g N_VPWR_c_213_n 0.0107398f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1000_g N_VPWR_c_222_n 0.0151087f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1001_g N_VPWR_c_222_n 0.0012662f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1000_g N_A_204_309#_c_262_n 0.0153218f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_A_204_309#_c_263_n 0.00426715f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1007_g Z 0.00319905f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_M1009_g Z 0.00617133f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A_M1000_g Z 0.00406561f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1001_g Z 0.0210047f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_c_169_n Z 4.74471e-19 $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_145 A Z 0.0260514f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A_c_171_n Z 0.00683006f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_M1000_g Z 9.99223e-19 $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1001_g Z 0.0120957f $X=2.74 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1000_g N_Z_c_296_n 0.0106702f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1007_g Z 0.00447149f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_M1000_g Z 0.00772664f $X=2.32 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1009_g Z 0.00358678f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_c_169_n Z 0.0226659f $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_154 A Z 0.0146926f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_M1007_g N_VGND_c_333_n 0.00112941f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_VGND_c_336_n 0.00357877f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_M1009_g N_VGND_c_336_n 0.00357877f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A_M1007_g N_VGND_c_337_n 0.00547239f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A_M1009_g N_VGND_c_337_n 0.0062648f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_M1007_g N_A_214_120#_c_378_n 0.0125883f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_161 N_A_M1009_g N_A_214_120#_c_378_n 0.0130314f $X=2.74 $Y=0.56 $X2=0 $Y2=0
cc_162 N_A_c_169_n N_A_214_120#_c_378_n 2.64617e-19 $X=2.815 $Y=1.16 $X2=0 $Y2=0
cc_163 A N_A_214_120#_c_378_n 0.00121919f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_164 A N_A_214_120#_c_379_n 0.0135366f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A_c_171_n N_A_214_120#_c_379_n 0.00554784f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_166 N_VPWR_c_213_n N_A_204_309#_M1002_s 0.00408188f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_167 N_VPWR_c_213_n N_A_204_309#_M1000_s 0.00411295f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_217_n N_A_204_309#_c_277_n 0.0109464f $X=1.41 $Y=2.53 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_213_n N_A_204_309#_c_277_n 0.00637602f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_215_n N_A_204_309#_c_262_n 0.0300999f $X=2 $Y=2.53 $X2=0 $Y2=0
cc_171 N_VPWR_c_219_n N_A_204_309#_c_262_n 0.00246817f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_213_n N_A_204_309#_c_262_n 0.00424653f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_219_n N_A_204_309#_c_282_n 0.0112958f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_213_n N_A_204_309#_c_282_n 0.00644886f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_175 N_VPWR_M1004_d N_A_204_309#_c_263_n 0.00435154f $X=1.44 $Y=1.545 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_216_n N_A_204_309#_c_263_n 0.0300999f $X=1.685 $Y=2.53 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_217_n N_A_204_309#_c_263_n 0.00263233f $X=1.41 $Y=2.53 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_213_n N_A_204_309#_c_263_n 0.008611f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_179 N_VPWR_c_222_n N_Z_M1000_d 0.00290085f $X=2.275 $Y=2.53 $X2=0 $Y2=0
cc_180 N_VPWR_c_213_n N_Z_M1001_d 0.00210122f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_181 N_VPWR_c_219_n Z 0.0225048f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_182 N_VPWR_c_213_n Z 0.0132695f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_183 N_A_204_309#_c_262_n N_Z_M1000_d 0.004872f $X=2.445 $Y=1.975 $X2=0 $Y2=0
cc_184 N_A_204_309#_M1000_s Z 0.00167813f $X=2.395 $Y=1.485 $X2=0 $Y2=0
cc_185 N_A_204_309#_c_262_n Z 0.0129015f $X=2.445 $Y=1.975 $X2=0 $Y2=0
cc_186 N_A_204_309#_c_262_n N_Z_c_296_n 0.0291967f $X=2.445 $Y=1.975 $X2=0 $Y2=0
cc_187 N_A_204_309#_c_263_n N_Z_c_296_n 0.0232998f $X=1.775 $Y=1.765 $X2=0 $Y2=0
cc_188 N_Z_M1007_s N_VGND_c_337_n 0.00216833f $X=2.395 $Y=0.235 $X2=0 $Y2=0
cc_189 N_Z_c_296_n N_A_214_120#_c_382_n 0.00512817f $X=2.365 $Y=1.57 $X2=0 $Y2=0
cc_190 N_Z_M1007_s N_A_214_120#_c_378_n 0.00304167f $X=2.395 $Y=0.235 $X2=0
+ $Y2=0
cc_191 Z N_A_214_120#_c_378_n 0.0158016f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_192 N_VGND_c_337_n N_A_214_120#_M1003_d 0.00220811f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_193 N_VGND_c_337_n N_A_214_120#_M1005_d 0.00296726f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_337_n N_A_214_120#_M1009_d 0.00210127f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_M1003_s N_A_214_120#_c_382_n 0.00304947f $X=1.48 $Y=0.235 $X2=0
+ $Y2=0
cc_196 N_VGND_c_333_n N_A_214_120#_c_382_n 0.0160613f $X=1.615 $Y=0.36 $X2=0
+ $Y2=0
cc_197 N_VGND_c_335_n N_A_214_120#_c_382_n 0.00232396f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_336_n N_A_214_120#_c_382_n 0.00232396f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_337_n N_A_214_120#_c_382_n 0.00970544f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_336_n N_A_214_120#_c_378_n 0.0543564f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_201 N_VGND_c_337_n N_A_214_120#_c_378_n 0.0339092f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_336_n N_A_214_120#_c_408_n 0.0165329f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_337_n N_A_214_120#_c_408_n 0.00939218f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_332_n N_A_214_120#_c_380_n 0.0188389f $X=0.68 $Y=0.38 $X2=0
+ $Y2=0
cc_205 N_VGND_c_335_n N_A_214_120#_c_380_n 0.0181389f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_337_n N_A_214_120#_c_380_n 0.0100822f $X=2.99 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__lpflow_inputisolatch_1.spice
* Created: Thu Aug 27 14:25:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__lpflow_inputisolatch_1.pex.spice"
.subckt sky130_fd_sc_hd__lpflow_inputisolatch_1  VNB VPB SLEEP_B D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* SLEEP_B	SLEEP_B
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_SLEEP_B_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_193_47#_M1010_d N_A_27_47#_M1010_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_381_47# N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.1092 PD=0.802308 PS=1.36 NRD=32.628 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_A_476_47#_M1014_d N_A_193_47#_M1014_g A_381_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0621 AS=0.0609231 PD=0.705 PS=0.687692 NRD=21.66 NRS=38.076 M=1
+ R=2.4 SA=75000.7 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1001 A_575_47# N_A_27_47#_M1001_g N_A_476_47#_M1014_d VNB NSHORT L=0.15 W=0.36
+ AD=0.0486 AS=0.0621 PD=0.63 PS=0.705 NRD=26.664 NRS=0 M=1 R=2.4 SA=75001.2
+ SB=75000.6 A=0.054 P=1.02 MULT=1
MM1005 N_VGND_M1005_d N_A_629_21#_M1005_g A_575_47# VNB NSHORT L=0.15 W=0.36
+ AD=0.0936 AS=0.0486 PD=1.24 PS=0.63 NRD=0 NRS=26.664 M=1 R=2.4 SA=75001.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1008 N_VGND_M1008_d N_A_476_47#_M1008_g N_A_629_21#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_Q_M1006_d N_A_476_47#_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_VPWR_M1012_d N_SLEEP_B_M1012_g N_A_27_47#_M1012_s VPB PHIGHVT L=0.15
+ W=0.55 AD=0.07425 AS=0.143 PD=0.82 PS=1.62 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_A_193_47#_M1002_d N_A_27_47#_M1002_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.55 AD=0.143 AS=0.07425 PD=1.62 PS=0.82 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1013 A_381_369# N_D_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.115623 AS=0.1664 PD=1.16528 PS=1.8 NRD=38.6711 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_A_476_47#_M1009_d N_A_27_47#_M1009_g A_381_369# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.0758774 PD=0.69 PS=0.764717 NRD=0 NRS=58.9227 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_560_413# N_A_193_47#_M1003_g N_A_476_47#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07245 AS=0.0567 PD=0.765 PS=0.69 NRD=55.1009 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_629_21#_M1011_g A_560_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1134 AS=0.07245 PD=1.38 PS=0.765 NRD=2.3443 NRS=55.1009 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_476_47#_M1007_g N_A_629_21#_M1007_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1000 N_Q_M1000_d N_A_476_47#_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
c_110 VPB 0 1.54137e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__lpflow_inputisolatch_1.pxi.spice"
*
.ends
*
*

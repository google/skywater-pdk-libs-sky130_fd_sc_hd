* File: sky130_fd_sc_hd__a21boi_4.spice.pex
* Created: Thu Aug 27 14:00:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BOI_4%B1_N 3 7 8 11 13
c34 3 0 1.29412e-19 $X=0.505 $Y=1.985
r35 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=1.325
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.16
+ $X2=0.565 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.16 $X2=0.565 $Y2=1.16
r38 8 12 9.79176 $w=4.61e-07 $l=3.7e-07 $layer=LI1_cond $X=0.397 $Y=1.53
+ $X2=0.397 $Y2=1.16
r39 7 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.625 $Y=0.56
+ $X2=0.625 $Y2=0.995
r40 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=1.985
+ $X2=0.505 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 35 37 41 43 46 48 54 60 61 72
c117 61 0 1.29412e-19 $X=0.962 $Y=1.19
c118 12 0 2.99299e-20 $X=1.455 $Y=1.985
r119 71 72 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.445 $Y=1.16
+ $X2=2.745 $Y2=1.16
r120 70 71 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.315 $Y=1.16
+ $X2=2.445 $Y2=1.16
r121 67 68 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.885 $Y=1.16
+ $X2=2.015 $Y2=1.16
r122 66 67 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=1.585 $Y=1.16
+ $X2=1.885 $Y2=1.16
r123 65 66 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.455 $Y=1.16
+ $X2=1.585 $Y2=1.16
r124 55 70 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.235 $Y=1.16
+ $X2=2.315 $Y2=1.16
r125 55 68 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.235 $Y=1.16
+ $X2=2.015 $Y2=1.16
r126 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.235
+ $Y=1.16 $X2=2.235 $Y2=1.16
r127 52 65 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.215 $Y=1.16
+ $X2=1.455 $Y2=1.16
r128 52 62 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.215 $Y=1.16
+ $X2=1.155 $Y2=1.16
r129 51 54 37.9191 $w=3.08e-07 $l=1.02e-06 $layer=LI1_cond $X=1.215 $Y=1.19
+ $X2=2.235 $Y2=1.19
r130 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r131 49 61 0.255944 $w=3.1e-07 $l=1.43e-07 $layer=LI1_cond $X=1.105 $Y=1.19
+ $X2=0.962 $Y2=1.19
r132 49 51 4.08931 $w=3.08e-07 $l=1.1e-07 $layer=LI1_cond $X=1.105 $Y=1.19
+ $X2=1.215 $Y2=1.19
r133 47 61 6.62803 $w=2.27e-07 $l=1.81273e-07 $layer=LI1_cond $X=0.905 $Y=1.345
+ $X2=0.962 $Y2=1.19
r134 47 48 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.785
r135 46 61 6.62803 $w=2.27e-07 $l=1.55e-07 $layer=LI1_cond $X=0.962 $Y=1.035
+ $X2=0.962 $Y2=1.19
r136 45 46 9.70478 $w=2.83e-07 $l=2.4e-07 $layer=LI1_cond $X=0.962 $Y=0.795
+ $X2=0.962 $Y2=1.035
r137 44 60 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=1.895
+ $X2=0.29 $Y2=1.895
r138 43 48 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.82 $Y=1.895
+ $X2=0.905 $Y2=1.785
r139 43 44 19.1201 $w=2.18e-07 $l=3.65e-07 $layer=LI1_cond $X=0.82 $Y=1.895
+ $X2=0.455 $Y2=1.895
r140 42 58 5.18785 $w=1.8e-07 $l=1.78e-07 $layer=LI1_cond $X=0.445 $Y=0.705
+ $X2=0.267 $Y2=0.705
r141 41 45 7.27854 $w=1.8e-07 $l=1.81505e-07 $layer=LI1_cond $X=0.82 $Y=0.705
+ $X2=0.962 $Y2=0.795
r142 41 42 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=0.82 $Y=0.705
+ $X2=0.445 $Y2=0.705
r143 35 58 2.62307 $w=3.55e-07 $l=9e-08 $layer=LI1_cond $X=0.267 $Y=0.615
+ $X2=0.267 $Y2=0.705
r144 35 37 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.267 $Y=0.615
+ $X2=0.267 $Y2=0.36
r145 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.16
r146 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.985
r147 28 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=0.995
+ $X2=2.445 $Y2=1.16
r148 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.445 $Y=0.995
+ $X2=2.445 $Y2=0.56
r149 24 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.16
r150 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.985
r151 21 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.16
r152 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r153 17 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.325
+ $X2=1.885 $Y2=1.16
r154 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.885 $Y=1.325
+ $X2=1.885 $Y2=1.985
r155 14 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=0.995
+ $X2=1.585 $Y2=1.16
r156 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.585 $Y=0.995
+ $X2=1.585 $Y2=0.56
r157 10 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.325
+ $X2=1.455 $Y2=1.16
r158 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.455 $Y=1.325
+ $X2=1.455 $Y2=1.985
r159 7 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=0.995
+ $X2=1.155 $Y2=1.16
r160 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.155 $Y=0.995
+ $X2=1.155 $Y2=0.56
r161 2 60 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.485 $X2=0.29 $Y2=2
r162 1 58 182 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.7
r163 1 37 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%A2 3 7 8 10 13 15 17 20 22 24 27 31 32 35
+ 36 37 38 41 54 55
c126 35 0 3.12905e-20 $X=3.375 $Y=1.592
c127 32 0 3.88689e-19 $X=3.195 $Y=1.16
c128 8 0 6.41563e-20 $X=5.365 $Y=0.995
r129 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.285
+ $Y=1.16 $X2=6.285 $Y2=1.16
r130 52 54 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.225 $Y=1.16
+ $X2=6.285 $Y2=1.16
r131 50 52 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.945 $Y=1.16
+ $X2=6.225 $Y2=1.16
r132 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.945
+ $Y=1.16 $X2=5.945 $Y2=1.16
r133 48 50 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.795 $Y=1.16
+ $X2=5.945 $Y2=1.16
r134 47 51 6.45503 $w=6.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.605 $Y=1.39
+ $X2=5.945 $Y2=1.39
r135 46 48 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=5.605 $Y=1.16
+ $X2=5.795 $Y2=1.16
r136 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.605
+ $Y=1.16 $X2=5.605 $Y2=1.16
r137 43 46 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=5.365 $Y=1.16
+ $X2=5.605 $Y2=1.16
r138 38 55 1.4239 $w=6.28e-07 $l=7.5e-08 $layer=LI1_cond $X=6.21 $Y=1.39
+ $X2=6.285 $Y2=1.39
r139 38 51 5.03112 $w=6.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.21 $Y=1.39
+ $X2=5.945 $Y2=1.39
r140 36 47 1.61376 $w=6.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=1.39
+ $X2=5.605 $Y2=1.39
r141 36 37 11.207 $w=6.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.52 $Y=1.39
+ $X2=5.205 $Y2=1.39
r142 35 37 93.732 $w=2.23e-07 $l=1.83e-06 $layer=LI1_cond $X=3.375 $Y=1.592
+ $X2=5.205 $Y2=1.592
r143 32 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.16
+ $X2=3.195 $Y2=1.325
r144 32 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.16
+ $X2=3.195 $Y2=0.995
r145 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.16 $X2=3.195 $Y2=1.16
r146 29 35 7.21695 $w=2.25e-07 $l=2.22047e-07 $layer=LI1_cond $X=3.202 $Y=1.48
+ $X2=3.375 $Y2=1.592
r147 29 31 10.6893 $w=3.43e-07 $l=3.2e-07 $layer=LI1_cond $X=3.202 $Y=1.48
+ $X2=3.202 $Y2=1.16
r148 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.325
+ $X2=6.225 $Y2=1.16
r149 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.225 $Y=1.325
+ $X2=6.225 $Y2=1.985
r150 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=1.16
r151 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.225 $Y=0.995
+ $X2=6.225 $Y2=0.56
r152 18 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.325
+ $X2=5.795 $Y2=1.16
r153 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.795 $Y=1.325
+ $X2=5.795 $Y2=1.985
r154 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=1.16
r155 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=0.56
r156 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.365 $Y=1.325
+ $X2=5.365 $Y2=1.16
r157 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.365 $Y=1.325
+ $X2=5.365 $Y2=1.985
r158 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.365 $Y=0.995
+ $X2=5.365 $Y2=1.16
r159 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.365 $Y=0.995
+ $X2=5.365 $Y2=0.56
r160 7 41 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.215 $Y=0.56
+ $X2=3.215 $Y2=0.995
r161 3 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.205 $Y=1.985
+ $X2=3.205 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29
r72 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.455
+ $Y=1.16 $X2=4.455 $Y2=1.16
r73 35 39 31.9862 $w=2.43e-07 $l=6.8e-07 $layer=LI1_cond $X=3.775 $Y=1.187
+ $X2=4.455 $Y2=1.187
r74 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=1.16 $X2=3.775 $Y2=1.16
r75 29 39 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=4.795 $Y=1.187
+ $X2=4.455 $Y2=1.187
r76 29 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.795
+ $Y=1.16 $X2=4.795 $Y2=1.16
r77 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.935 $Y=1.295
+ $X2=4.935 $Y2=1.985
r78 22 25 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=4.935 $Y=1.142
+ $X2=4.935 $Y2=1.295
r79 22 42 27.535 $w=3.05e-07 $l=1.4e-07 $layer=POLY_cond $X=4.935 $Y=1.142
+ $X2=4.795 $Y2=1.142
r80 22 24 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.935 $Y=0.99
+ $X2=4.935 $Y2=0.56
r81 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.505 $Y=1.295
+ $X2=4.505 $Y2=1.985
r82 15 42 57.0367 $w=3.05e-07 $l=2.9e-07 $layer=POLY_cond $X=4.505 $Y=1.142
+ $X2=4.795 $Y2=1.142
r83 15 18 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=4.505 $Y=1.142
+ $X2=4.505 $Y2=1.295
r84 15 38 9.83392 $w=3.05e-07 $l=5e-08 $layer=POLY_cond $X=4.505 $Y=1.142
+ $X2=4.455 $Y2=1.142
r85 15 17 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.505 $Y=0.99
+ $X2=4.505 $Y2=0.56
r86 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.075 $Y=1.295
+ $X2=4.075 $Y2=1.985
r87 8 38 74.7378 $w=3.05e-07 $l=3.8e-07 $layer=POLY_cond $X=4.075 $Y=1.142
+ $X2=4.455 $Y2=1.142
r88 8 11 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=4.075 $Y=1.142
+ $X2=4.075 $Y2=1.295
r89 8 34 59.0035 $w=3.05e-07 $l=3e-07 $layer=POLY_cond $X=4.075 $Y=1.142
+ $X2=3.775 $Y2=1.142
r90 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.075 $Y=0.99
+ $X2=4.075 $Y2=0.56
r91 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.645 $Y=1.295
+ $X2=3.645 $Y2=1.985
r92 1 34 25.5682 $w=3.05e-07 $l=1.3e-07 $layer=POLY_cond $X=3.645 $Y=1.142
+ $X2=3.775 $Y2=1.142
r93 1 4 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=3.645 $Y=1.142
+ $X2=3.645 $Y2=1.295
r94 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.645 $Y=0.99
+ $X2=3.645 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%VPWR 1 2 3 4 5 20 24 28 32 36 39 40 42 43
+ 44 46 54 67 68 71 74 77
r117 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r118 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r122 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r123 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r124 62 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r125 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 59 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.29 $Y2=2.72
r127 59 61 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.455 $Y=2.72
+ $X2=4.83 $Y2=2.72
r128 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r129 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r130 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.43 $Y2=2.72
r132 55 57 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.91 $Y2=2.72
r133 54 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=4.29 $Y2=2.72
r134 54 57 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=3.91 $Y2=2.72
r135 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r136 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r137 50 53 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r138 50 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r139 49 52 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r140 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 47 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=0.755 $Y2=2.72
r142 47 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.885 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.43 $Y2=2.72
r144 46 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r145 44 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 42 64 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=5.75 $Y2=2.72
r147 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=6.01 $Y2=2.72
r148 41 67 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=6.67 $Y2=2.72
r149 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=2.72
+ $X2=6.01 $Y2=2.72
r150 39 61 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=2.72
+ $X2=5.15 $Y2=2.72
r152 38 64 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.75 $Y2=2.72
r153 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.72
+ $X2=5.15 $Y2=2.72
r154 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=2.635
+ $X2=6.01 $Y2=2.72
r155 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.01 $Y=2.635
+ $X2=6.01 $Y2=2.36
r156 30 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=2.635
+ $X2=5.15 $Y2=2.72
r157 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.15 $Y=2.635
+ $X2=5.15 $Y2=2.36
r158 26 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.635
+ $X2=4.29 $Y2=2.72
r159 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.29 $Y=2.635
+ $X2=4.29 $Y2=2.36
r160 22 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=2.72
r161 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=2.36
r162 18 71 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2.72
r163 18 20 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.755 $Y=2.635
+ $X2=0.755 $Y2=2.34
r164 5 36 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.485 $X2=6.01 $Y2=2.36
r165 4 32 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.485 $X2=5.15 $Y2=2.36
r166 3 28 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=1.485 $X2=4.29 $Y2=2.36
r167 2 24 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.485 $X2=3.43 $Y2=2.36
r168 1 20 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.485 $X2=0.72 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%A_223_297# 1 2 3 4 5 6 7 22 24 26 28 29 34
+ 36 40 42 44 46 55 56
c81 29 0 2.24772e-19 $X=3.095 $Y=1.99
c82 28 0 1.93847e-19 $X=4.625 $Y=1.99
r83 51 53 34.3608 $w=3.16e-07 $l=8.9e-07 $layer=LI1_cond $X=2.1 $Y=2.205
+ $X2=2.99 $Y2=2.205
r84 44 58 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=6.475 $Y=2.105
+ $X2=6.475 $Y2=1.99
r85 44 46 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=6.475 $Y=2.105
+ $X2=6.475 $Y2=2.3
r86 43 56 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.665 $Y=1.99 $X2=5.575
+ $Y2=1.99
r87 42 58 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=6.345 $Y=1.99
+ $X2=6.475 $Y2=1.99
r88 42 43 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.345 $Y=1.99
+ $X2=5.665 $Y2=1.99
r89 38 56 2.23839 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=5.575 $Y=2.105
+ $X2=5.575 $Y2=1.99
r90 38 40 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=5.575 $Y=2.105
+ $X2=5.575 $Y2=2.3
r91 37 55 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.815 $Y=1.99
+ $X2=4.72 $Y2=1.99
r92 36 56 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.485 $Y=1.99 $X2=5.575
+ $Y2=1.99
r93 36 37 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.485 $Y=1.99
+ $X2=4.815 $Y2=1.99
r94 32 55 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=4.72 $Y=2.105
+ $X2=4.72 $Y2=1.99
r95 32 34 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=4.72 $Y=2.105
+ $X2=4.72 $Y2=2.3
r96 29 53 4.97931 $w=3.16e-07 $l=2.62298e-07 $layer=LI1_cond $X=3.095 $Y=1.99
+ $X2=2.99 $Y2=2.205
r97 29 31 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.095 $Y=1.99
+ $X2=3.86 $Y2=1.99
r98 28 55 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.625 $Y=1.99
+ $X2=4.72 $Y2=1.99
r99 28 31 38.3313 $w=2.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.625 $Y=1.99
+ $X2=3.86 $Y2=1.99
r100 27 49 3.05549 $w=2.5e-07 $l=9.8e-08 $layer=LI1_cond $X=1.355 $Y=2.34
+ $X2=1.257 $Y2=2.34
r101 26 51 6.93673 $w=3.16e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.935 $Y=2.34
+ $X2=2.1 $Y2=2.205
r102 26 27 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=1.935 $Y=2.34
+ $X2=1.355 $Y2=2.34
r103 22 49 3.89731 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=1.257 $Y=2.215
+ $X2=1.257 $Y2=2.34
r104 22 24 14.5035 $w=1.93e-07 $l=2.55e-07 $layer=LI1_cond $X=1.257 $Y=2.215
+ $X2=1.257 $Y2=1.96
r105 7 58 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.485 $X2=6.44 $Y2=1.96
r106 7 46 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=6.3
+ $Y=1.485 $X2=6.44 $Y2=2.3
r107 6 40 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=5.44
+ $Y=1.485 $X2=5.58 $Y2=2.3
r108 5 55 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=4.58
+ $Y=1.485 $X2=4.72 $Y2=1.96
r109 5 34 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.58
+ $Y=1.485 $X2=4.72 $Y2=2.3
r110 4 31 600 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.485 $X2=3.86 $Y2=1.99
r111 3 53 600 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.485 $X2=2.99 $Y2=2.3
r112 2 51 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.485 $X2=2.1 $Y2=2.36
r113 1 49 600 $w=1.7e-07 $l=8.77596e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.485 $X2=1.245 $Y2=2.3
r114 1 24 600 $w=1.7e-07 $l=5.36074e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.485 $X2=1.245 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%Y 1 2 3 4 5 6 19 23 25 28 31 35 38 43 44 45
+ 46 49 55
c79 44 0 9.67612e-20 $X=2.715 $Y=0.795
c80 35 0 6.41563e-20 $X=4.72 $Y=0.76
c81 31 0 3.39132e-19 $X=3.365 $Y=0.785
r82 49 55 1.06318 $w=4.48e-07 $l=4e-08 $layer=LI1_cond $X=2.57 $Y=1.81 $X2=2.53
+ $Y2=1.81
r83 46 49 2.83704 $w=4.5e-07 $l=1.45e-07 $layer=LI1_cond $X=2.715 $Y=1.81
+ $X2=2.57 $Y2=1.81
r84 46 55 0.611329 $w=4.48e-07 $l=2.3e-08 $layer=LI1_cond $X=2.507 $Y=1.81
+ $X2=2.53 $Y2=1.81
r85 46 51 22.2471 $w=4.48e-07 $l=8.37e-07 $layer=LI1_cond $X=2.507 $Y=1.81
+ $X2=1.67 $Y2=1.81
r86 33 35 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=3.86 $Y=0.785 $X2=4.72
+ $Y2=0.785
r87 31 45 5.8804 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=3.365 $Y=0.785
+ $X2=3.255 $Y2=0.785
r88 31 33 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.365 $Y=0.785
+ $X2=3.86 $Y2=0.785
r89 30 44 7.37517 $w=1.85e-07 $l=1.45e-07 $layer=LI1_cond $X=2.86 $Y=0.795
+ $X2=2.715 $Y2=0.795
r90 30 45 21.9045 $w=1.98e-07 $l=3.95e-07 $layer=LI1_cond $X=2.86 $Y=0.795
+ $X2=3.255 $Y2=0.795
r91 28 46 4.4023 $w=2.9e-07 $l=2.25e-07 $layer=LI1_cond $X=2.715 $Y=1.585
+ $X2=2.715 $Y2=1.81
r92 27 44 0.213802 $w=2.9e-07 $l=1e-07 $layer=LI1_cond $X=2.715 $Y=0.895
+ $X2=2.715 $Y2=0.795
r93 27 28 27.4202 $w=2.88e-07 $l=6.9e-07 $layer=LI1_cond $X=2.715 $Y=0.895
+ $X2=2.715 $Y2=1.585
r94 26 43 4.74942 $w=2.1e-07 $l=1.13248e-07 $layer=LI1_cond $X=2.325 $Y=0.78
+ $X2=2.23 $Y2=0.74
r95 25 44 7.37517 $w=1.85e-07 $l=1.52315e-07 $layer=LI1_cond $X=2.57 $Y=0.78
+ $X2=2.715 $Y2=0.795
r96 25 26 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.57 $Y=0.78
+ $X2=2.325 $Y2=0.78
r97 21 43 1.70532 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.23 $Y=0.615
+ $X2=2.23 $Y2=0.74
r98 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.23 $Y=0.615
+ $X2=2.23 $Y2=0.42
r99 20 38 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.37 $Y=0.74
+ $X2=1.37 $Y2=0.535
r100 19 43 4.74942 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=2.23 $Y2=0.74
r101 19 20 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=1.465 $Y2=0.74
r102 6 55 600 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.53 $Y2=1.89
r103 5 51 600 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.485 $X2=1.67 $Y2=1.85
r104 4 35 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.58
+ $Y=0.235 $X2=4.72 $Y2=0.76
r105 3 33 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.235 $X2=3.86 $Y2=0.76
r106 2 43 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.23 $Y2=0.76
r107 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.23 $Y2=0.42
r108 1 38 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.235 $X2=1.37 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%VGND 1 2 3 4 5 18 24 28 31 37 38 40 41 43
+ 44 45 65 66 71 77
c101 40 0 1.51849e-19 $X=5.485 $Y=0
r102 76 77 8.65265 $w=6.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.22 $X2=3.085
+ $Y2=0.22
r103 73 76 0.196078 $w=6.08e-07 $l=1e-08 $layer=LI1_cond $X=2.99 $Y=0.22 $X2=3
+ $Y2=0.22
r104 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r105 70 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r106 69 73 9.01961 $w=6.08e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=0.22
+ $X2=2.99 $Y2=0.22
r107 69 71 7.67225 $w=6.08e-07 $l=3.5e-08 $layer=LI1_cond $X=2.53 $Y=0.22
+ $X2=2.495 $Y2=0.22
r108 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r109 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r110 63 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r111 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r112 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r113 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r114 57 60 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r115 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r116 56 59 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=5.29
+ $Y2=0
r117 56 77 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=3.085 $Y2=0
r118 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r119 53 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r120 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r121 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r122 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 45 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r124 43 62 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.345 $Y=0
+ $X2=6.21 $Y2=0
r125 43 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.345 $Y=0 $X2=6.475
+ $Y2=0
r126 42 65 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.67
+ $Y2=0
r127 42 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.475
+ $Y2=0
r128 40 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=0
+ $X2=5.29 $Y2=0
r129 40 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.58
+ $Y2=0
r130 39 62 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.675 $Y=0
+ $X2=6.21 $Y2=0
r131 39 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.675 $Y=0 $X2=5.58
+ $Y2=0
r132 37 52 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.61
+ $Y2=0
r133 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=0 $X2=1.8
+ $Y2=0
r134 33 52 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.105 $Y=0
+ $X2=1.61 $Y2=0
r135 31 48 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.69
+ $Y2=0
r136 31 35 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=0.912 $Y=0
+ $X2=0.912 $Y2=0.36
r137 31 33 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.912 $Y=0
+ $X2=1.105 $Y2=0
r138 26 44 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=0.085
+ $X2=6.475 $Y2=0
r139 26 28 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.475 $Y=0.085
+ $X2=6.475 $Y2=0.38
r140 22 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0
r141 22 24 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0.4
r142 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.8
+ $Y2=0
r143 21 71 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.965 $Y=0
+ $X2=2.495 $Y2=0
r144 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=0.085 $X2=1.8
+ $Y2=0
r145 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.8 $Y=0.085
+ $X2=1.8 $Y2=0.36
r146 5 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.235 $X2=6.44 $Y2=0.38
r147 4 24 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.44
+ $Y=0.235 $X2=5.58 $Y2=0.4
r148 3 76 91 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.235 $X2=3 $Y2=0.36
r149 2 18 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.235 $X2=1.8 $Y2=0.36
r150 1 35 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.235 $X2=0.9 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_4%A_658_47# 1 2 3 4 13 19 22 23 24 27
c45 1 0 1.87282e-19 $X=3.29 $Y=0.235
r46 25 27 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.01 $Y=0.735
+ $X2=6.01 $Y2=0.395
r47 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.845 $Y=0.82
+ $X2=6.01 $Y2=0.735
r48 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.845 $Y=0.82
+ $X2=5.315 $Y2=0.82
r49 20 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.185 $Y=0.735
+ $X2=5.315 $Y2=0.82
r50 20 22 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.185 $Y=0.735
+ $X2=5.185 $Y2=0.7
r51 19 30 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0.505
+ $X2=5.185 $Y2=0.38
r52 19 22 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=5.185 $Y=0.505
+ $X2=5.185 $Y2=0.7
r53 15 18 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=3.43 $Y=0.38 $X2=4.29
+ $Y2=0.38
r54 13 30 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=5.055 $Y=0.38
+ $X2=5.185 $Y2=0.38
r55 13 18 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=5.055 $Y=0.38
+ $X2=4.29 $Y2=0.38
r56 4 27 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=5.87
+ $Y=0.235 $X2=6.01 $Y2=0.395
r57 3 30 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.235 $X2=5.15 $Y2=0.36
r58 3 22 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=5.01
+ $Y=0.235 $X2=5.15 $Y2=0.7
r59 2 18 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.15
+ $Y=0.235 $X2=4.29 $Y2=0.42
r60 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.235 $X2=3.43 $Y2=0.42
.ends


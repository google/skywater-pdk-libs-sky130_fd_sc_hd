* File: sky130_fd_sc_hd__o211ai_4.spice
* Created: Tue Sep  1 19:20:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o211ai_4.pex.spice"
.subckt sky130_fd_sc_hd__o211ai_4  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_A_27_47#_M1006_d N_A1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_27_47#_M1009_d N_A1_M1009_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1019 N_A_27_47#_M1009_d N_A1_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_A2_M1005_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1005_d N_A2_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75005.1 A=0.0975 P=1.6 MULT=1
MM1018 N_A_27_47#_M1018_d N_A2_M1018_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75004.7 A=0.0975 P=1.6 MULT=1
MM1028 N_A_27_47#_M1018_d N_A2_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.09425 PD=0.93 PS=0.94 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75004.2 A=0.0975 P=1.6 MULT=1
MM1031 N_A_27_47#_M1031_d N_A1_M1031_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.09425 PD=0.96 PS=0.94 NRD=1.836 NRS=1.836 M=1 R=4.33333
+ SA=75003.2 SB=75003.8 A=0.0975 P=1.6 MULT=1
MM1002 N_A_806_47#_M1002_d N_B1_M1002_g N_A_27_47#_M1031_d VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.10075 PD=0.93 PS=0.96 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75003.7 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1026 N_A_806_47#_M1002_d N_B1_M1026_g N_A_27_47#_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1012 A_1314_47# N_B1_M1012_g N_A_27_47#_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.091 PD=0.92 PS=0.93 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1016 N_Y_M1016_d N_C1_M1016_g A_1314_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75004.9 SB=75002
+ A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1016_d N_C1_M1020_g N_A_806_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1022 N_Y_M1022_d N_C1_M1022_g N_A_806_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.8
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1022_d N_C1_M1015_g A_978_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=19.38 M=1 R=4.33333 SA=75006.2 SB=75000.8
+ A=0.0975 P=1.6 MULT=1
MM1025 A_978_47# N_B1_M1025_g N_A_27_47#_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.25675 PD=0.97 PS=2.09 NRD=19.38 NRS=0 M=1 R=4.33333 SA=75006.7
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_110_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75007
+ A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1013_d N_A1_M1013_g N_A_110_297#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75006.6 A=0.15 P=2.3 MULT=1
MM1017 N_VPWR_M1013_d N_A1_M1017_g N_A_110_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75006.2
+ A=0.15 P=2.3 MULT=1
MM1007 N_Y_M1007_d N_A2_M1007_g N_A_110_297#_M1017_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75005.7 A=0.15 P=2.3 MULT=1
MM1010 N_Y_M1007_d N_A2_M1010_g N_A_110_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75005.3 A=0.15 P=2.3 MULT=1
MM1021 N_Y_M1021_d N_A2_M1021_g N_A_110_297#_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75004.9 A=0.15 P=2.3 MULT=1
MM1027 N_Y_M1021_d N_A2_M1027_g N_A_110_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1029 N_VPWR_M1029_d N_A1_M1029_g N_A_110_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75004 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1029_d N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=3.9203 NRS=0 M=1 R=6.66667 SA=75003.7 SB=75003.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1 SB=75003.1 A=0.15
+ P=2.3 MULT=1
MM1011 N_VPWR_M1003_d N_B1_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.14
+ AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5 SB=75002.7
+ A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.9 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1000_d N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.4 SB=75001.9
+ A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_C1_M1024_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.8 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1024_d N_C1_M1030_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75006.2 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1023 N_VPWR_M1023_d N_B1_M1023_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1 AD=0.675
+ AS=0.135 PD=3.35 PS=1.27 NRD=76.8103 NRS=0 M=1 R=6.66667 SA=75006.6 SB=75000.6
+ A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.161 P=19.61
*
.include "sky130_fd_sc_hd__o211ai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a2bb2oi_4.spice.pex
* Created: Thu Aug 27 14:03:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 30 31
+ 32 35 36 38 39 50 54
c125 50 0 1.66018e-19 $X=1.31 $Y=1.16
c126 36 0 2.73979e-19 $X=3.41 $Y=1.16
c127 35 0 1.10598e-19 $X=3.41 $Y=1.16
c128 32 0 6.77964e-20 $X=1.555 $Y=1.53
c129 15 0 8.27827e-20 $X=1.31 $Y=0.995
r130 48 50 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.235 $Y=1.16
+ $X2=1.31 $Y2=1.16
r131 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.235
+ $Y=1.16 $X2=1.235 $Y2=1.16
r132 46 48 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.235 $Y2=1.16
r133 45 49 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.555 $Y=1.18
+ $X2=1.235 $Y2=1.18
r134 44 46 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.555 $Y=1.16
+ $X2=0.89 $Y2=1.16
r135 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.555
+ $Y=1.16 $X2=0.555 $Y2=1.16
r136 41 44 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.555 $Y2=1.16
r137 39 45 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.555 $Y2=1.18
r138 39 54 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.23 $Y2=1.18
r139 38 49 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=1.385 $Y=1.18
+ $X2=1.235 $Y2=1.18
r140 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.16 $X2=3.41 $Y2=1.16
r141 33 35 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.16
r142 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.41 $Y2=1.445
r143 31 32 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=1.555 $Y2=1.53
r144 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.47 $Y=1.445
+ $X2=1.555 $Y2=1.53
r145 29 38 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.47 $Y=1.285
+ $X2=1.385 $Y2=1.18
r146 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.47 $Y=1.285
+ $X2=1.47 $Y2=1.445
r147 25 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.16
r148 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.41 $Y=1.325
+ $X2=3.41 $Y2=1.985
r149 22 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.16
r150 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r151 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r152 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r153 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r154 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r155 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r156 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r157 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r158 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r159 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r160 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.985
r161 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r162 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
c65 40 0 1.66018e-19 $X=2.91 $Y=1.16
c66 1 0 1.79953e-19 $X=1.73 $Y=0.995
r67 39 41 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.91 $Y=1.16 $X2=2.99
+ $Y2=1.16
r68 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.91
+ $Y=1.16 $X2=2.91 $Y2=1.16
r69 37 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.91 $Y2=1.16
r70 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r71 34 36 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.89 $Y=1.16
+ $X2=2.15 $Y2=1.16
r72 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=1.16 $X2=1.89 $Y2=1.16
r73 31 34 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.89 $Y2=1.16
r74 29 40 46.3045 $w=1.98e-07 $l=8.35e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=2.91 $Y2=1.175
r75 29 35 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=2.075 $Y=1.175
+ $X2=1.89 $Y2=1.175
r76 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.16
r77 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.99 $Y=1.325
+ $X2=2.99 $Y2=1.985
r78 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.16
r79 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r80 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r81 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r82 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r83 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r84 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r85 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r86 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r87 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r88 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r89 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325 $X2=1.73
+ $Y2=1.985
r90 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r91 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995 $X2=1.73
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A_751_21# 1 2 3 4 5 6 19 21 24 26 28 31 33
+ 35 38 40 42 45 47 56 57 58 61 63 67 69 73 77 79 83 87 89 92 93 94 95 97 98 100
+ 107
c215 31 0 1.4428e-20 $X=4.25 $Y=1.985
c216 24 0 9.61704e-20 $X=3.83 $Y=1.985
r217 101 103 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.83 $Y=1.16
+ $X2=4.25 $Y2=1.16
r218 91 92 17.6068 $w=3.58e-07 $l=5.5e-07 $layer=LI1_cond $X=9.395 $Y=0.905
+ $X2=9.395 $Y2=1.455
r219 90 98 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=8.925 $Y=0.82
+ $X2=8.76 $Y2=0.815
r220 89 91 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=9.215 $Y=0.82
+ $X2=9.395 $Y2=0.905
r221 89 90 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.215 $Y=0.82
+ $X2=8.925 $Y2=0.82
r222 88 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.885 $Y=1.54
+ $X2=8.76 $Y2=1.54
r223 87 92 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=9.215 $Y=1.54
+ $X2=9.395 $Y2=1.455
r224 87 88 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.215 $Y=1.54
+ $X2=8.885 $Y2=1.54
r225 81 98 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.76 $Y=0.725
+ $X2=8.76 $Y2=0.815
r226 81 83 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.76 $Y=0.725
+ $X2=8.76 $Y2=0.39
r227 80 95 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0.815
+ $X2=7.92 $Y2=0.815
r228 79 98 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0.815
+ $X2=8.76 $Y2=0.815
r229 79 80 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=8.595 $Y=0.815
+ $X2=8.085 $Y2=0.815
r230 78 97 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.045 $Y=1.54
+ $X2=7.92 $Y2=1.54
r231 77 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.635 $Y=1.54
+ $X2=8.76 $Y2=1.54
r232 77 78 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.635 $Y=1.54
+ $X2=8.045 $Y2=1.54
r233 71 95 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.92 $Y=0.725
+ $X2=7.92 $Y2=0.815
r234 71 73 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=0.725
+ $X2=7.92 $Y2=0.39
r235 70 94 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0.815
+ $X2=7.08 $Y2=0.815
r236 69 95 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=0.815
+ $X2=7.92 $Y2=0.815
r237 69 70 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.755 $Y=0.815
+ $X2=7.245 $Y2=0.815
r238 65 94 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.08 $Y=0.725
+ $X2=7.08 $Y2=0.815
r239 65 67 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.08 $Y=0.725
+ $X2=7.08 $Y2=0.39
r240 64 93 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0.815
+ $X2=6.24 $Y2=0.815
r241 63 94 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0.815
+ $X2=7.08 $Y2=0.815
r242 63 64 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.915 $Y=0.815
+ $X2=6.405 $Y2=0.815
r243 59 93 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.815
r244 59 61 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.39
r245 57 93 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.075 $Y=0.82
+ $X2=6.24 $Y2=0.815
r246 57 58 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.075 $Y=0.82
+ $X2=5.725 $Y2=0.82
r247 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.64 $Y=0.905
+ $X2=5.725 $Y2=0.82
r248 55 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.64 $Y=0.905
+ $X2=5.64 $Y2=1.075
r249 54 107 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.945 $Y=1.16
+ $X2=5.09 $Y2=1.16
r250 54 105 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.945 $Y=1.16
+ $X2=4.67 $Y2=1.16
r251 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.945
+ $Y=1.16 $X2=4.945 $Y2=1.16
r252 50 105 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=4.265 $Y=1.16
+ $X2=4.67 $Y2=1.16
r253 50 103 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.265 $Y=1.16
+ $X2=4.25 $Y2=1.16
r254 49 53 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.265 $Y=1.16
+ $X2=4.945 $Y2=1.16
r255 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=1.16 $X2=4.265 $Y2=1.16
r256 47 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.555 $Y=1.16
+ $X2=5.64 $Y2=1.075
r257 47 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.555 $Y=1.16
+ $X2=4.945 $Y2=1.16
r258 43 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.16
r259 43 45 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.09 $Y=1.325
+ $X2=5.09 $Y2=1.985
r260 40 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=1.16
r261 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.09 $Y=0.995
+ $X2=5.09 $Y2=0.56
r262 36 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.16
r263 36 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.67 $Y=1.325
+ $X2=4.67 $Y2=1.985
r264 33 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=0.995
+ $X2=4.67 $Y2=1.16
r265 33 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.67 $Y=0.995
+ $X2=4.67 $Y2=0.56
r266 29 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.16
r267 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.25 $Y=1.325
+ $X2=4.25 $Y2=1.985
r268 26 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=1.16
r269 26 28 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.25 $Y=0.995
+ $X2=4.25 $Y2=0.56
r270 22 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.325
+ $X2=3.83 $Y2=1.16
r271 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.83 $Y=1.325
+ $X2=3.83 $Y2=1.985
r272 19 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.16
r273 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r274 6 100 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=8.625
+ $Y=1.485 $X2=8.76 $Y2=1.62
r275 5 97 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=7.785
+ $Y=1.485 $X2=7.92 $Y2=1.62
r276 4 83 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.625
+ $Y=0.235 $X2=8.76 $Y2=0.39
r277 3 73 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.785
+ $Y=0.235 $X2=7.92 $Y2=0.39
r278 2 67 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.945
+ $Y=0.235 $X2=7.08 $Y2=0.39
r279 1 61 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A1_N 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
r82 39 41 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.155 $Y=1.16
+ $X2=7.29 $Y2=1.16
r83 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.155
+ $Y=1.16 $X2=7.155 $Y2=1.16
r84 37 39 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=6.87 $Y=1.16
+ $X2=7.155 $Y2=1.16
r85 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.45 $Y=1.16
+ $X2=6.87 $Y2=1.16
r86 34 36 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.135 $Y=1.16
+ $X2=6.45 $Y2=1.16
r87 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.135
+ $Y=1.16 $X2=6.135 $Y2=1.16
r88 31 34 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.03 $Y=1.16
+ $X2=6.135 $Y2=1.16
r89 29 40 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.695 $Y=1.175
+ $X2=7.155 $Y2=1.175
r90 29 35 31.0545 $w=1.98e-07 $l=5.6e-07 $layer=LI1_cond $X=6.695 $Y=1.175
+ $X2=6.135 $Y2=1.175
r91 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.16
r92 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.29 $Y=1.325
+ $X2=7.29 $Y2=1.985
r93 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.16
r94 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=0.56
r95 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.16
r96 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.87 $Y=1.325
+ $X2=6.87 $Y2=1.985
r97 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=1.16
r98 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.87 $Y=0.995
+ $X2=6.87 $Y2=0.56
r99 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r101 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r103 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r104 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r105 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A2_N 1 3 6 8 10 13 15 17 20 22 24 27 29 40
+ 41
r80 39 41 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=8.855 $Y=1.16
+ $X2=8.97 $Y2=1.16
r81 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.855
+ $Y=1.16 $X2=8.855 $Y2=1.16
r82 37 39 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=8.55 $Y=1.16
+ $X2=8.855 $Y2=1.16
r83 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.13 $Y=1.16
+ $X2=8.55 $Y2=1.16
r84 34 36 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=7.835 $Y=1.16
+ $X2=8.13 $Y2=1.16
r85 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.835
+ $Y=1.16 $X2=7.835 $Y2=1.16
r86 31 34 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.71 $Y=1.16
+ $X2=7.835 $Y2=1.16
r87 29 40 43.2545 $w=1.98e-07 $l=7.8e-07 $layer=LI1_cond $X=8.075 $Y=1.175
+ $X2=8.855 $Y2=1.175
r88 29 35 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=8.075 $Y=1.175
+ $X2=7.835 $Y2=1.175
r89 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.97 $Y=1.325
+ $X2=8.97 $Y2=1.16
r90 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.97 $Y=1.325
+ $X2=8.97 $Y2=1.985
r91 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.97 $Y=0.995
+ $X2=8.97 $Y2=1.16
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.97 $Y=0.995
+ $X2=8.97 $Y2=0.56
r93 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.55 $Y=1.325
+ $X2=8.55 $Y2=1.16
r94 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.55 $Y=1.325
+ $X2=8.55 $Y2=1.985
r95 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.55 $Y=0.995
+ $X2=8.55 $Y2=1.16
r96 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.55 $Y=0.995
+ $X2=8.55 $Y2=0.56
r97 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.13 $Y=1.325
+ $X2=8.13 $Y2=1.16
r98 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.13 $Y=1.325
+ $X2=8.13 $Y2=1.985
r99 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.13 $Y=0.995
+ $X2=8.13 $Y2=1.16
r100 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.13 $Y=0.995
+ $X2=8.13 $Y2=0.56
r101 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.71 $Y=1.325
+ $X2=7.71 $Y2=1.16
r102 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.71 $Y=1.325
+ $X2=7.71 $Y2=1.985
r103 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.71 $Y=0.995
+ $X2=7.71 $Y2=1.16
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.71 $Y=0.995
+ $X2=7.71 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A_27_297# 1 2 3 4 5 6 7 24 28 29 30 34 38
+ 42 44 46 47 50 52 54 56 61 63 65 68
c96 44 0 1.25804e-19 $X=3.62 $Y=1.965
c97 42 0 1.48175e-19 $X=3.495 $Y=1.88
r98 54 70 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.295 $X2=5.3
+ $Y2=2.38
r99 54 56 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=5.3 $Y=2.295 $X2=5.3
+ $Y2=1.65
r100 53 68 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.575 $Y=2.38
+ $X2=4.455 $Y2=2.38
r101 52 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=2.38
+ $X2=5.3 $Y2=2.38
r102 52 53 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.135 $Y=2.38
+ $X2=4.575 $Y2=2.38
r103 48 68 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.295
+ $X2=4.455 $Y2=2.38
r104 48 50 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=4.455 $Y=2.295
+ $X2=4.455 $Y2=1.96
r105 46 68 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.335 $Y=2.38
+ $X2=4.455 $Y2=2.38
r106 46 47 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.335 $Y=2.38
+ $X2=3.745 $Y2=2.38
r107 45 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.62 $Y=2.295
+ $X2=3.745 $Y2=2.38
r108 44 67 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=1.965
+ $X2=3.62 $Y2=1.88
r109 44 45 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=3.62 $Y=1.965
+ $X2=3.62 $Y2=2.295
r110 43 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.905 $Y=1.88
+ $X2=2.78 $Y2=1.88
r111 42 67 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.495 $Y=1.88
+ $X2=3.62 $Y2=1.88
r112 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.495 $Y=1.88
+ $X2=2.905 $Y2=1.88
r113 39 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=1.88
+ $X2=1.94 $Y2=1.88
r114 38 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=1.88
+ $X2=2.78 $Y2=1.88
r115 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.655 $Y=1.88
+ $X2=2.065 $Y2=1.88
r116 35 61 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.215 $Y=1.88
+ $X2=1.095 $Y2=1.88
r117 34 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=1.88
+ $X2=1.94 $Y2=1.88
r118 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.815 $Y=1.88
+ $X2=1.215 $Y2=1.88
r119 31 61 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.795
+ $X2=1.095 $Y2=1.88
r120 30 59 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=1.54
r121 30 31 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=1.795
r122 28 59 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=1.095 $Y2=1.54
r123 28 29 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.975 $Y=1.54
+ $X2=0.425 $Y2=1.54
r124 24 26 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=2.33
r125 22 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.425 $Y2=1.54
r126 22 24 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.255 $Y2=1.65
r127 7 70 400 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2.33
r128 7 56 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=1.65
r129 6 50 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=1.96
r130 5 67 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=1.96
r131 4 65 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=1.96
r132 3 63 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r133 2 61 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r134 2 59 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.62
r135 1 26 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.33
r136 1 24 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 52 54 69 73 80 81 84 87 90
r144 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r145 87 88 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r146 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 81 91 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=7.13 $Y2=2.72
r148 80 81 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r149 78 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.205 $Y=2.72
+ $X2=7.08 $Y2=2.72
r150 78 80 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=7.205 $Y=2.72
+ $X2=9.43 $Y2=2.72
r151 77 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r152 77 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r153 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r154 74 87 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.365 $Y=2.72
+ $X2=6.26 $Y2=2.72
r155 74 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.365 $Y=2.72
+ $X2=6.67 $Y2=2.72
r156 73 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=7.08 $Y2=2.72
r157 73 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.955 $Y=2.72
+ $X2=6.67 $Y2=2.72
r158 72 88 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=6.21 $Y2=2.72
r159 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 69 87 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.155 $Y=2.72
+ $X2=6.26 $Y2=2.72
r161 69 71 176.476 $w=1.68e-07 $l=2.705e-06 $layer=LI1_cond $X=6.155 $Y=2.72
+ $X2=3.45 $Y2=2.72
r162 68 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r163 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r164 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r165 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r166 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r167 62 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r169 59 84 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=0.7 $Y2=2.72
r170 59 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=1.15 $Y2=2.72
r171 54 84 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.7 $Y2=2.72
r172 54 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r173 52 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r174 52 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r175 50 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=2.99 $Y2=2.72
r176 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=3.2 $Y2=2.72
r177 49 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.45 $Y2=2.72
r178 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.2 $Y2=2.72
r179 47 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r180 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.36 $Y2=2.72
r181 46 67 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.99 $Y2=2.72
r182 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.36 $Y2=2.72
r183 44 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.15 $Y2=2.72
r184 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.52 $Y2=2.72
r185 43 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=2.07 $Y2=2.72
r186 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.52 $Y2=2.72
r187 39 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=2.635
+ $X2=7.08 $Y2=2.72
r188 39 41 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.08 $Y=2.635
+ $X2=7.08 $Y2=1.96
r189 35 87 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=2.635
+ $X2=6.26 $Y2=2.72
r190 35 37 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=6.26 $Y=2.635
+ $X2=6.26 $Y2=1.96
r191 31 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.72
r192 31 33 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.3
r193 27 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.72
r194 27 29 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.36 $Y=2.635
+ $X2=2.36 $Y2=2.3
r195 23 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r196 23 25 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.3
r197 19 84 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r198 19 21 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=1.96
r199 6 41 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.945
+ $Y=1.485 $X2=7.08 $Y2=1.96
r200 5 37 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.96
r201 4 33 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=2.3
r202 3 29 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=2.3
r203 2 25 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.3
r204 1 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%Y 1 2 3 4 5 6 19 25 28 31 35 37 38 39 43
+ 45 46 50 51 57
c97 19 0 8.27827e-20 $X=2.865 $Y=0.775
r98 51 57 13.0959 $w=2.18e-07 $l=2.5e-07 $layer=LI1_cond $X=4.855 $Y=1.87
+ $X2=4.855 $Y2=1.62
r99 50 57 2.3196 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=4.855 $Y=1.615
+ $X2=4.855 $Y2=1.62
r100 41 43 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.88 $Y=0.725
+ $X2=4.88 $Y2=0.39
r101 40 46 4.10651 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=4.205 $Y=0.815
+ $X2=3.975 $Y2=0.815
r102 39 41 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.715 $Y=0.815
+ $X2=4.88 $Y2=0.725
r103 39 40 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.715 $Y=0.815
+ $X2=4.205 $Y2=0.815
r104 37 50 3.58108 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.745 $Y=1.515
+ $X2=4.855 $Y2=1.515
r105 37 38 32.1636 $w=1.98e-07 $l=5.8e-07 $layer=LI1_cond $X=4.745 $Y=1.515
+ $X2=4.165 $Y2=1.515
r106 33 38 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=4.04 $Y=1.515
+ $X2=4.165 $Y2=1.515
r107 33 47 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=4.04 $Y=1.515
+ $X2=3.83 $Y2=1.515
r108 33 35 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.04 $Y=1.615
+ $X2=4.04 $Y2=1.62
r109 29 46 2.1123 $w=3.3e-07 $l=1.1811e-07 $layer=LI1_cond $X=4.04 $Y=0.725
+ $X2=3.975 $Y2=0.815
r110 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=0.725
+ $X2=4.04 $Y2=0.39
r111 28 47 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.83 $Y=1.415 $X2=3.83
+ $Y2=1.515
r112 27 46 2.1123 $w=1.7e-07 $l=1.84594e-07 $layer=LI1_cond $X=3.83 $Y=0.905
+ $X2=3.975 $Y2=0.815
r113 27 28 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.83 $Y=0.905
+ $X2=3.83 $Y2=1.415
r114 25 46 4.10651 $w=1.8e-07 $l=2.3e-07 $layer=LI1_cond $X=3.745 $Y=0.815
+ $X2=3.975 $Y2=0.815
r115 25 45 46.2121 $w=1.78e-07 $l=7.5e-07 $layer=LI1_cond $X=3.745 $Y=0.815
+ $X2=2.995 $Y2=0.815
r116 21 24 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=1.94 $Y=0.775
+ $X2=2.78 $Y2=0.775
r117 19 45 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.865 $Y=0.775
+ $X2=2.995 $Y2=0.775
r118 19 24 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.775
+ $X2=2.78 $Y2=0.775
r119 6 57 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.62
r120 5 35 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=1.62
r121 4 43 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.39
r122 3 31 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.39
r123 2 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.73
r124 1 21 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A_1139_297# 1 2 3 4 5 18 22 23 26 28 30 31
+ 32 36 40 43 49
r67 38 40 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.185 $Y=2.295
+ $X2=9.185 $Y2=1.96
r68 37 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.465 $Y=2.38
+ $X2=8.34 $Y2=2.38
r69 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.06 $Y=2.38
+ $X2=9.185 $Y2=2.295
r70 36 37 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=9.06 $Y=2.38
+ $X2=8.465 $Y2=2.38
r71 33 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.625 $Y=2.38
+ $X2=7.5 $Y2=2.38
r72 32 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.215 $Y=2.38
+ $X2=8.34 $Y2=2.38
r73 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.215 $Y=2.38
+ $X2=7.625 $Y2=2.38
r74 31 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=2.295 $X2=7.5
+ $Y2=2.38
r75 30 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=1.625 $X2=7.5
+ $Y2=1.54
r76 30 31 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.5 $Y=1.625 $X2=7.5
+ $Y2=2.295
r77 29 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.78 $Y=1.54 $X2=6.66
+ $Y2=1.54
r78 28 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.375 $Y=1.54
+ $X2=7.5 $Y2=1.54
r79 28 29 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=7.375 $Y=1.54
+ $X2=6.78 $Y2=1.54
r80 24 43 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=1.625
+ $X2=6.66 $Y2=1.54
r81 24 26 32.4125 $w=2.38e-07 $l=6.75e-07 $layer=LI1_cond $X=6.66 $Y=1.625
+ $X2=6.66 $Y2=2.3
r82 22 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.54 $Y=1.54 $X2=6.66
+ $Y2=1.54
r83 22 23 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=6.54 $Y=1.54
+ $X2=5.985 $Y2=1.54
r84 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.82 $Y=1.65
+ $X2=5.82 $Y2=2.33
r85 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.82 $Y=1.625
+ $X2=5.985 $Y2=1.54
r86 16 18 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.82 $Y=1.625
+ $X2=5.82 $Y2=1.65
r87 5 40 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.045
+ $Y=1.485 $X2=9.18 $Y2=1.96
r88 4 49 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.205
+ $Y=1.485 $X2=8.34 $Y2=2.3
r89 3 47 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=2.3
r90 3 45 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.485 $X2=7.5 $Y2=1.62
r91 2 43 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.62
r92 2 26 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=2.3
r93 1 20 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.485 $X2=5.82 $Y2=2.33
r94 1 18 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.485 $X2=5.82 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 48
+ 52 56 60 63 64 65 66 68 69 71 72 74 75 77 78 79 81 107 108 114 119 125
r159 124 125 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.235
+ $X2=5.905 $Y2=0.235
r160 121 124 1.30821 $w=6.38e-07 $l=7e-08 $layer=LI1_cond $X=5.75 $Y=0.235
+ $X2=5.82 $Y2=0.235
r161 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r162 118 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r163 117 121 8.59681 $w=6.38e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=0.235
+ $X2=5.75 $Y2=0.235
r164 117 119 8.73487 $w=6.38e-07 $l=7.5e-08 $layer=LI1_cond $X=5.29 $Y=0.235
+ $X2=5.215 $Y2=0.235
r165 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r166 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r167 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r168 105 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r169 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r170 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r171 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r172 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r173 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r174 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r175 96 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r176 95 125 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=5.905 $Y2=0
r177 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r178 92 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r179 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r180 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r181 89 115 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=1.15 $Y2=0
r182 88 89 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r183 86 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.1
+ $Y2=0
r184 86 88 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=3.45 $Y2=0
r185 85 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r186 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r187 82 111 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r188 82 84 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r189 81 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.1
+ $Y2=0
r190 81 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=0
+ $X2=0.69 $Y2=0
r191 79 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r192 79 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r193 77 104 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.095 $Y=0
+ $X2=8.97 $Y2=0
r194 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.095 $Y=0 $X2=9.18
+ $Y2=0
r195 76 107 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.265 $Y=0
+ $X2=9.43 $Y2=0
r196 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0 $X2=9.18
+ $Y2=0
r197 74 101 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.255 $Y=0
+ $X2=8.05 $Y2=0
r198 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=0 $X2=8.34
+ $Y2=0
r199 73 104 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.425 $Y=0
+ $X2=8.97 $Y2=0
r200 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=0 $X2=8.34
+ $Y2=0
r201 71 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.415 $Y=0
+ $X2=7.13 $Y2=0
r202 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=0 $X2=7.5
+ $Y2=0
r203 70 101 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.585 $Y=0
+ $X2=8.05 $Y2=0
r204 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=0 $X2=7.5
+ $Y2=0
r205 68 95 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r206 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0 $X2=6.66
+ $Y2=0
r207 67 98 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.13 $Y2=0
r208 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.66
+ $Y2=0
r209 65 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.37
+ $Y2=0
r210 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.375 $Y=0 $X2=4.46
+ $Y2=0
r211 63 88 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.45
+ $Y2=0
r212 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0 $X2=3.62
+ $Y2=0
r213 62 91 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=4.37
+ $Y2=0
r214 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.62
+ $Y2=0
r215 58 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.18 $Y=0.085
+ $X2=9.18 $Y2=0
r216 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.18 $Y=0.085
+ $X2=9.18 $Y2=0.39
r217 54 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0
r218 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0.39
r219 50 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r220 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.39
r221 46 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0
r222 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0.39
r223 45 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=0 $X2=4.46
+ $Y2=0
r224 45 119 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.545 $Y=0
+ $X2=5.215 $Y2=0
r225 40 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r226 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.39
r227 36 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r228 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.39
r229 32 114 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r230 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.39
r231 28 111 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r232 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r233 9 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.045
+ $Y=0.235 $X2=9.18 $Y2=0.39
r234 8 56 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.205
+ $Y=0.235 $X2=8.34 $Y2=0.39
r235 7 52 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.5 $Y2=0.39
r236 6 48 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r237 5 124 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=5.165
+ $Y=0.235 $X2=5.82 $Y2=0.39
r238 4 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.39
r239 3 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.39
r240 2 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.39
r241 1 30 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2OI_4%A_109_47# 1 2 3 4 15 17 18 19 20 25
c48 20 0 1.79953e-19 $X=1.48 $Y=0.725
r49 23 25 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.36 $Y=0.365
+ $X2=3.2 $Y2=0.365
r50 21 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=0.365
+ $X2=1.48 $Y2=0.365
r51 21 23 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=1.605 $Y=0.365
+ $X2=2.36 $Y2=0.365
r52 20 30 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.48 $Y=0.725 $X2=1.48
+ $Y2=0.815
r53 19 28 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.48 $Y=0.475
+ $X2=1.48 $Y2=0.365
r54 19 20 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.48 $Y=0.475
+ $X2=1.48 $Y2=0.725
r55 17 30 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=1.48 $Y2=0.815
r56 17 18 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=0.815
+ $X2=0.845 $Y2=0.815
r57 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.845 $Y2=0.815
r58 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.725
+ $X2=0.68 $Y2=0.39
r59 4 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.39
r60 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.39
r61 2 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.73
r62 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r63 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
.ends


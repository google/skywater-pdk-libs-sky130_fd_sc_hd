* File: sky130_fd_sc_hd__nor2_1.pxi.spice
* Created: Tue Sep  1 19:17:34 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2_1%B N_B_c_29_n N_B_M1003_g N_B_M1002_g B N_B_c_31_n
+ PM_SKY130_FD_SC_HD__NOR2_1%B
x_PM_SKY130_FD_SC_HD__NOR2_1%A N_A_M1000_g N_A_c_55_n N_A_M1001_g A N_A_c_57_n
+ PM_SKY130_FD_SC_HD__NOR2_1%A
x_PM_SKY130_FD_SC_HD__NOR2_1%Y N_Y_M1003_d N_Y_M1002_s N_Y_c_88_n N_Y_c_90_n
+ N_Y_c_83_n N_Y_c_86_n N_Y_c_84_n Y PM_SKY130_FD_SC_HD__NOR2_1%Y
x_PM_SKY130_FD_SC_HD__NOR2_1%VPWR N_VPWR_M1000_d N_VPWR_c_120_n N_VPWR_c_121_n
+ VPWR N_VPWR_c_122_n N_VPWR_c_119_n VPWR PM_SKY130_FD_SC_HD__NOR2_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR2_1%VGND N_VGND_M1003_s N_VGND_M1001_d N_VGND_c_135_n
+ N_VGND_c_136_n N_VGND_c_137_n N_VGND_c_138_n VGND N_VGND_c_139_n
+ N_VGND_c_140_n PM_SKY130_FD_SC_HD__NOR2_1%VGND
cc_1 VNB N_B_c_29_n 0.0218606f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB B 0.00935867f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_B_c_31_n 0.0387673f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_c_55_n 0.0218599f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_5 VNB A 0.00908315f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_A_c_57_n 0.0418519f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_Y_c_83_n 0.00516135f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_8 VNB N_Y_c_84_n 0.00134186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VPWR_c_119_n 0.0609879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_135_n 0.0101633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_136_n 0.030355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_137_n 0.0104214f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_13 VNB N_VGND_c_138_n 0.0318347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_139_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_140_n 0.104147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VPB N_B_M1002_g 0.0255613f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_17 VPB B 0.00121238f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_18 VPB N_B_c_31_n 0.00866622f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_19 VPB N_A_M1000_g 0.0246007f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_20 VPB A 0.00119303f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_21 VPB N_A_c_57_n 0.0123812f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_22 VPB N_Y_c_83_n 0.001574f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_23 VPB N_Y_c_86_n 0.00741865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB Y 0.0306411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_VPWR_c_120_n 0.0115529f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_26 VPB N_VPWR_c_121_n 0.047482f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_27 VPB N_VPWR_c_122_n 0.0295367f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_28 VPB N_VPWR_c_119_n 0.0433341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 N_B_M1002_g N_A_M1000_g 0.0432238f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_30 N_B_c_29_n N_A_c_55_n 0.00936712f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_31 N_B_c_31_n N_A_c_57_n 0.0525909f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_32 N_B_M1002_g N_Y_c_88_n 0.0131302f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_33 B N_Y_c_88_n 6.64606e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_34 N_B_c_29_n N_Y_c_90_n 0.00545148f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_35 N_B_c_29_n N_Y_c_83_n 0.0100046f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_36 B N_Y_c_83_n 0.0188125f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_37 N_B_M1002_g N_Y_c_86_n 8.84614e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_38 B N_Y_c_86_n 0.0241802f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_39 N_B_c_31_n N_Y_c_86_n 0.00646558f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_40 N_B_c_29_n N_Y_c_84_n 0.00269062f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_41 N_B_M1002_g Y 0.0139173f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_42 N_B_M1002_g N_VPWR_c_122_n 0.00541964f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_43 N_B_M1002_g N_VPWR_c_119_n 0.0105205f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_44 N_B_c_29_n N_VGND_c_136_n 0.00342736f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_45 B N_VGND_c_136_n 0.0188825f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_46 N_B_c_31_n N_VGND_c_136_n 0.00597918f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_47 N_B_c_29_n N_VGND_c_139_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_48 N_B_c_29_n N_VGND_c_140_n 0.0104829f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_Y_c_88_n 0.0043289f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_c_55_n N_Y_c_90_n 0.00545148f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_51 N_A_M1000_g N_Y_c_83_n 0.00765851f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A_c_55_n N_Y_c_83_n 0.0052733f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_53 A N_Y_c_83_n 0.0182565f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_54 N_A_c_57_n N_Y_c_83_n 0.00361863f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_c_55_n N_Y_c_84_n 0.00341202f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A_c_57_n N_Y_c_84_n 0.00169761f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_M1000_g Y 0.00224347f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_58 N_A_M1000_g N_VPWR_c_121_n 0.00457701f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_59 A N_VPWR_c_121_n 0.0265465f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A_c_57_n N_VPWR_c_121_n 0.00744853f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_VPWR_c_122_n 0.00585385f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VPWR_c_119_n 0.011501f $X=0.83 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_c_55_n N_VGND_c_138_n 0.00344349f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_64 A N_VGND_c_138_n 0.0212807f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_VGND_c_138_n 0.00661799f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_55_n N_VGND_c_139_n 0.00541359f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_c_55_n N_VGND_c_140_n 0.0105016f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_68 N_Y_c_88_n A_109_297# 0.00415017f $X=0.605 $Y=1.58 $X2=-0.19 $Y2=-0.24
cc_69 Y N_VPWR_c_122_n 0.0192029f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_70 N_Y_M1002_s N_VPWR_c_119_n 0.00209863f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_71 Y N_VPWR_c_119_n 0.0123358f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_72 N_Y_c_90_n N_VGND_c_136_n 0.0243336f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_73 N_Y_c_90_n N_VGND_c_138_n 0.02434f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_74 N_Y_c_90_n N_VGND_c_139_n 0.0188862f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_75 N_Y_M1003_d N_VGND_c_140_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_76 N_Y_c_90_n N_VGND_c_140_n 0.0122123f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_77 A_109_297# N_VPWR_c_119_n 0.00897657f $X=0.545 $Y=1.485 $X2=0.15 $Y2=2.125

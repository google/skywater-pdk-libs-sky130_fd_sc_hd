* File: sky130_fd_sc_hd__o21ai_2.spice.pex
* Created: Thu Aug 27 14:35:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21AI_2%A1 1 3 6 10 14 15 18 19 23 24 35
c75 35 0 1.494e-19 $X=1.865 $Y=0.995
c76 18 0 1.95305e-19 $X=1.865 $Y=1.16
r77 23 24 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=0.285 $Y=1.16
+ $X2=0.285 $Y2=1.445
r78 23 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r79 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.16
+ $X2=1.865 $Y2=1.325
r80 19 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.16
+ $X2=1.865 $Y2=0.995
r81 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.16 $X2=1.865 $Y2=1.16
r82 16 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.53
+ $X2=0.285 $Y2=1.53
r83 15 18 8.94038 $w=4.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.847 $Y=1.53
+ $X2=1.847 $Y2=1.16
r84 15 16 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=1.6 $Y=1.53
+ $X2=0.45 $Y2=1.53
r85 14 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.885 $Y=0.56
+ $X2=1.885 $Y2=0.995
r86 10 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.845 $Y=1.985
+ $X2=1.845 $Y2=1.325
r87 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.485 $Y=1.305
+ $X2=0.485 $Y2=1.985
r88 1 4 22.2839 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=0.485 $Y=1.132
+ $X2=0.485 $Y2=1.305
r89 1 29 33.4517 $w=3.45e-07 $l=2e-07 $layer=POLY_cond $X=0.485 $Y=1.132
+ $X2=0.285 $Y2=1.132
r90 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.485 $Y=0.96 $X2=0.485
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%A2 1 3 6 8 10 13 15 21 22
c53 13 0 1.95305e-19 $X=1.345 $Y=1.985
r54 20 22 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.25 $Y=1.16
+ $X2=1.345 $Y2=1.16
r55 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.25
+ $Y=1.16 $X2=1.25 $Y2=1.16
r56 17 20 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.915 $Y=1.16
+ $X2=1.25 $Y2=1.16
r57 15 21 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.145 $Y=1.175
+ $X2=1.25 $Y2=1.175
r58 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=1.16
r59 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=1.985
r60 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=0.995
+ $X2=1.345 $Y2=1.16
r61 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.345 $Y=0.995
+ $X2=1.345 $Y2=0.56
r62 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=1.16
r63 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=1.985
r64 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=0.915 $Y2=1.16
r65 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.915 $Y=0.995
+ $X2=0.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%B1 1 3 6 8 10 12 15 17 18 19 22
r48 22 24 31.0968 $w=3.41e-07 $l=2.2e-07 $layer=POLY_cond $X=2.745 $Y=1.142
+ $X2=2.965 $Y2=1.142
r49 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.16 $X2=2.965 $Y2=1.16
r50 18 19 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.972 $Y=0.85
+ $X2=2.972 $Y2=1.16
r51 13 22 22.0049 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.142
r52 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.985
r53 10 22 22.0049 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=2.745 $Y=0.96
+ $X2=2.745 $Y2=1.142
r54 10 12 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.745 $Y=0.96
+ $X2=2.745 $Y2=0.56
r55 9 17 0.971436 $w=2.05e-07 $l=7.5e-08 $layer=POLY_cond $X=2.39 $Y=1.062
+ $X2=2.315 $Y2=1.062
r56 8 22 18.2091 $w=3.41e-07 $l=1.11355e-07 $layer=POLY_cond $X=2.67 $Y=1.062
+ $X2=2.745 $Y2=1.142
r57 8 9 90.5772 $w=2.05e-07 $l=2.8e-07 $layer=POLY_cond $X=2.67 $Y=1.062
+ $X2=2.39 $Y2=1.062
r58 4 17 26.2462 $w=1.5e-07 $l=1.03e-07 $layer=POLY_cond $X=2.315 $Y=1.165
+ $X2=2.315 $Y2=1.062
r59 4 6 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.315 $Y=1.165
+ $X2=2.315 $Y2=1.985
r60 1 17 26.2462 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=2.315 $Y=0.96
+ $X2=2.315 $Y2=1.062
r61 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.315 $Y=0.96 $X2=2.315
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%VPWR 1 2 3 10 12 16 18 20 22 24 32 41 45
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r57 33 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=2.72
+ $X2=2.075 $Y2=2.72
r58 33 35 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.24 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 32 44 4.59592 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=3.017 $Y2=2.72
r60 32 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.815 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r64 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 25 38 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.217 $Y2=2.72
r67 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.075 $Y2=2.72
r69 24 30 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=1.61
+ $Y2=2.72
r70 22 28 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 18 44 3.00327 $w=3.1e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=3.017 $Y2=2.72
r73 18 20 33.458 $w=3.08e-07 $l=9e-07 $layer=LI1_cond $X=2.97 $Y=2.635 $X2=2.97
+ $Y2=1.735
r74 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.72
r75 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.075 $Y=2.635
+ $X2=2.075 $Y2=2.34
r76 10 38 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.217 $Y2=2.72
r77 10 12 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=1.95
r78 3 20 300 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=1.485 $X2=2.96 $Y2=1.735
r79 2 16 600 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.485 $X2=2.075 $Y2=2.34
r80 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%A_112_297# 1 2 9 11 12 14
r19 11 14 1.386 $w=1.7e-07 $l=1.28938e-07 $layer=LI1_cond $X=1.525 $Y=2.38
+ $X2=1.62 $Y2=2.3
r20 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.525 $Y=2.38
+ $X2=0.825 $Y2=2.38
r21 7 12 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.715 $Y=2.295
+ $X2=0.825 $Y2=2.38
r22 7 9 18.0724 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=0.715 $Y=2.295
+ $X2=0.715 $Y2=1.95
r23 2 14 600 $w=1.7e-07 $l=9.05028e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.485 $X2=1.61 $Y2=2.3
r24 1 9 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=1.485 $X2=0.7 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%Y 1 2 3 10 13 14 15 16 22 30 40
c36 30 0 1.494e-19 $X=2.53 $Y=0.76
r37 30 33 45.9481 $w=2.08e-07 $l=8.7e-07 $layer=LI1_cond $X=2.54 $Y=0.76
+ $X2=2.54 $Y2=1.63
r38 16 22 2.11586 $w=1.8e-07 $l=1.17e-07 $layer=LI1_cond $X=2.527 $Y=1.875
+ $X2=2.41 $Y2=1.875
r39 16 33 6.98973 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=2.54 $Y=1.785
+ $X2=2.54 $Y2=1.63
r40 15 22 21.2576 $w=1.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.065 $Y=1.875
+ $X2=2.41 $Y2=1.875
r41 14 15 28.3434 $w=1.78e-07 $l=4.6e-07 $layer=LI1_cond $X=1.605 $Y=1.875
+ $X2=2.065 $Y2=1.875
r42 14 40 19.101 $w=1.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.605 $Y=1.875
+ $X2=1.295 $Y2=1.875
r43 13 40 7.62263 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.145 $Y=1.955
+ $X2=1.295 $Y2=1.955
r44 13 36 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=1.145 $Y=1.955
+ $X2=1.13 $Y2=1.955
r45 10 16 4.31573 $w=2.22e-07 $l=9e-08 $layer=LI1_cond $X=2.527 $Y=1.965
+ $X2=2.527 $Y2=1.875
r46 10 12 6.48936 $w=2.35e-07 $l=1.25e-07 $layer=LI1_cond $X=2.527 $Y=1.965
+ $X2=2.527 $Y2=2.09
r47 3 33 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.53 $Y2=1.63
r48 3 12 600 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.53 $Y2=2.09
r49 2 36 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.485 $X2=1.13 $Y2=1.96
r50 1 30 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.53 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%A_29_47# 1 2 3 4 15 17 18 21 23 25 26 27 29
+ 32
r73 32 35 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=2.97 $Y=0.34 $X2=2.97
+ $Y2=0.43
r74 28 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0.34
+ $X2=2.1 $Y2=0.34
r75 27 32 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=2.97 $Y2=0.34
r76 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.815 $Y=0.34
+ $X2=2.265 $Y2=0.34
r77 25 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.425 $X2=2.1
+ $Y2=0.34
r78 25 26 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.1 $Y=0.425 $X2=2.1
+ $Y2=0.715
r79 24 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=0.8
+ $X2=1.13 $Y2=0.8
r80 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.935 $Y=0.8
+ $X2=2.1 $Y2=0.715
r81 23 24 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.935 $Y=0.8
+ $X2=1.295 $Y2=0.8
r82 19 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.715
+ $X2=1.13 $Y2=0.8
r83 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.13 $Y=0.715
+ $X2=1.13 $Y2=0.4
r84 17 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0.8
+ $X2=1.13 $Y2=0.8
r85 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.965 $Y=0.8
+ $X2=0.435 $Y2=0.8
r86 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=0.715
+ $X2=0.435 $Y2=0.8
r87 13 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.27 $Y=0.715
+ $X2=0.27 $Y2=0.4
r88 4 35 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.96 $Y2=0.43
r89 3 31 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=0.235 $X2=2.1 $Y2=0.4
r90 2 21 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.235 $X2=1.13 $Y2=0.4
r91 1 15 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__O21AI_2%VGND 1 2 11 15 17 19 29 30 33 36
r52 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r53 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r56 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r57 26 29 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r58 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r59 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0 $X2=1.61
+ $Y2=0
r60 24 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.695 $Y=0 $X2=2.07
+ $Y2=0
r61 23 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r62 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r63 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r64 20 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r65 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.15
+ $Y2=0
r66 19 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.61
+ $Y2=0
r67 19 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.15
+ $Y2=0
r68 17 34 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.225 $Y=0
+ $X2=0.69 $Y2=0
r69 13 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0
r70 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.61 $Y=0.085
+ $X2=1.61 $Y2=0.38
r71 9 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r72 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.38
r73 2 15 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.42
+ $Y=0.235 $X2=1.61 $Y2=0.38
r74 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__clkinvlp_2.pex.spice
* Created: Thu Aug 27 14:12:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINVLP_2%A 3 5 7 8 10 12 15 17 18 19 20 21 26
r40 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r41 20 21 8.93773 $w=4.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.372 $Y=1.19
+ $X2=0.372 $Y2=1.53
r42 20 26 0.788623 $w=4.53e-07 $l=3e-08 $layer=LI1_cond $X=0.372 $Y=1.19
+ $X2=0.372 $Y2=1.16
r43 17 25 2.25938 $w=3.2e-07 $l=1.5e-08 $layer=POLY_cond $X=0.53 $Y=1.155
+ $X2=0.515 $Y2=1.155
r44 17 18 9.58664 $w=3.2e-07 $l=1.25e-07 $layer=POLY_cond $X=0.53 $Y=1.155
+ $X2=0.655 $Y2=1.155
r45 13 19 18.238 $w=2e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.185 $Y=1.17
+ $X2=1.15 $Y2=1.08
r46 13 15 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.185 $Y=1.17
+ $X2=1.185 $Y2=1.985
r47 10 19 18.238 $w=2e-07 $l=1.25499e-07 $layer=POLY_cond $X=1.065 $Y=0.99
+ $X2=1.15 $Y2=1.08
r48 10 12 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.065 $Y=0.99
+ $X2=1.065 $Y2=0.61
r49 9 18 9.58664 $w=1.75e-07 $l=1.57321e-07 $layer=POLY_cond $X=0.78 $Y=1.082
+ $X2=0.655 $Y2=1.155
r50 8 19 7.22026 $w=1.75e-07 $l=1.60997e-07 $layer=POLY_cond $X=0.99 $Y=1.082
+ $X2=1.15 $Y2=1.08
r51 8 9 83.9613 $w=1.75e-07 $l=2.1e-07 $layer=POLY_cond $X=0.99 $Y=1.082
+ $X2=0.78 $Y2=1.082
r52 5 18 14.7117 $w=1.5e-07 $l=1.69706e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.655 $Y2=1.155
r53 5 7 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.675 $Y=0.995
+ $X2=0.675 $Y2=0.61
r54 1 18 14.7117 $w=2.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.655 $Y=1.315
+ $X2=0.655 $Y2=1.155
r55 1 3 166.464 $w=2.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.655 $Y=1.315
+ $X2=0.655 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_2%VPWR 1 2 7 9 11 13 17 19 29
r21 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r22 23 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r23 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 20 25 4.39998 $w=1.8e-07 $l=2.78e-07 $layer=LI1_cond $X=0.555 $Y=2.715
+ $X2=0.277 $Y2=2.715
r25 20 22 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=0.555 $Y=2.715
+ $X2=1.15 $Y2=2.715
r26 19 28 4.34455 $w=1.8e-07 $l=2e-07 $layer=LI1_cond $X=1.44 $Y=2.715 $X2=1.64
+ $Y2=2.715
r27 19 22 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=1.44 $Y=2.715
+ $X2=1.15 $Y2=2.715
r28 17 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 13 16 27.2745 $w=2.98e-07 $l=7.1e-07 $layer=LI1_cond $X=1.59 $Y=1.63
+ $X2=1.59 $Y2=2.34
r31 11 28 3.04118 $w=3e-07 $l=1.1225e-07 $layer=LI1_cond $X=1.59 $Y=2.625
+ $X2=1.64 $Y2=2.715
r32 11 16 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.59 $Y=2.625
+ $X2=1.59 $Y2=2.34
r33 7 25 3.21294 $w=3.3e-07 $l=1.51456e-07 $layer=LI1_cond $X=0.39 $Y=2.625
+ $X2=0.277 $Y2=2.715
r34 7 9 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=0.39 $Y=2.625
+ $X2=0.39 $Y2=2
r35 2 16 400 $w=1.7e-07 $l=9.7857e-07 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.485 $X2=1.575 $Y2=2.34
r36 2 13 400 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.485 $X2=1.575 $Y2=1.63
r37 1 9 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.265
+ $Y=1.485 $X2=0.39 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_2%Y 1 2 7 8 9
r21 25 26 4.51417 $w=6.33e-07 $l=1.7e-07 $layer=LI1_cond $X=1.127 $Y=0.58
+ $X2=1.127 $Y2=0.75
r22 9 19 13.0158 $w=4.23e-07 $l=4.8e-07 $layer=LI1_cond $X=1.022 $Y=1.19
+ $X2=1.022 $Y2=1.67
r23 8 9 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.022 $Y=0.85
+ $X2=1.022 $Y2=1.19
r24 8 26 2.71163 $w=4.23e-07 $l=1e-07 $layer=LI1_cond $X=1.022 $Y=0.85 $X2=1.022
+ $Y2=0.75
r25 7 25 1.31851 $w=6.33e-07 $l=7e-08 $layer=LI1_cond $X=1.127 $Y=0.51 $X2=1.127
+ $Y2=0.58
r26 2 19 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=1.485 $X2=0.92 $Y2=1.67
r27 1 25 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.335 $X2=1.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINVLP_2%VGND 1 6 9 10 11 21 22
r16 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r17 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r18 18 21 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r19 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r20 11 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r21 11 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r22 9 14 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.23
+ $Y2=0
r23 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=0 $X2=0.46
+ $Y2=0
r24 8 18 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.69
+ $Y2=0
r25 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.46
+ $Y2=0
r26 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.46 $Y=0.085 $X2=0.46
+ $Y2=0
r27 4 6 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.46 $Y=0.085
+ $X2=0.46 $Y2=0.58
r28 1 6 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.335 $X2=0.46 $Y2=0.58
.ends


* NGSPICE file created from sky130_fd_sc_hd__a21boi_0.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VGND A2 a_400_47# VNB nshort w=420000u l=150000u
+  ad=3.717e+11p pd=3.45e+06u as=8.82e+10p ps=1.26e+06u
M1001 VPWR A1 a_300_369# VPB phighvt w=640000u l=150000u
+  ad=2.905e+11p pd=3.21e+06u as=3.488e+11p ps=3.65e+06u
M1002 VPWR B1_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VGND B1_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_300_369# a_27_47# Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1005 a_300_369# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=0p ps=0u
M1007 a_400_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
M1000 VPWR A a_207_413# VPB phighvt w=420000u l=150000u
+  ad=5.986e+11p pd=5e+06u as=1.218e+11p ps=1.42e+06u
M1001 a_297_47# a_27_413# a_207_413# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.092e+11p ps=1.36e+06u
M1002 VGND A a_297_47# VNB nshort w=420000u l=150000u
+  ad=3.118e+11p pd=3.34e+06u as=0p ps=0u
M1003 VPWR SLEEP a_27_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 a_207_413# a_27_413# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_207_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1006 X a_207_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1007 a_27_413# SLEEP VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o21a_4.spice.pex
* Created: Thu Aug 27 14:35:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21A_4%A_80_21# 1 2 3 10 12 15 17 19 22 24 26 29 31
+ 33 36 38 47 50 52 53 56 58 62 67 69 80
c129 62 0 1.78828e-19 $X=2.215 $Y=0.762
c130 53 0 1.69833e-19 $X=2.315 $Y=1.957
r131 77 78 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.655 $Y=1.16
+ $X2=1.765 $Y2=1.16
r132 76 77 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.655 $Y2=1.16
r133 75 76 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.225 $Y=1.16
+ $X2=1.335 $Y2=1.16
r134 74 75 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=1.16
+ $X2=1.225 $Y2=1.16
r135 73 74 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.795 $Y=1.16
+ $X2=0.905 $Y2=1.16
r136 59 67 4.19778 $w=2.42e-07 $l=1.05877e-07 $layer=LI1_cond $X=2.845 $Y=1.99
+ $X2=2.75 $Y2=1.967
r137 58 69 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=1.99
+ $X2=4.38 $Y2=1.99
r138 58 59 68.6455 $w=2.28e-07 $l=1.37e-06 $layer=LI1_cond $X=4.215 $Y=1.99
+ $X2=2.845 $Y2=1.99
r139 54 67 2.23415 $w=1.9e-07 $l=1.38e-07 $layer=LI1_cond $X=2.75 $Y=2.105
+ $X2=2.75 $Y2=1.967
r140 54 56 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.75 $Y=2.105
+ $X2=2.75 $Y2=2.3
r141 52 67 4.19778 $w=2.42e-07 $l=9.98749e-08 $layer=LI1_cond $X=2.655 $Y=1.957
+ $X2=2.75 $Y2=1.967
r142 52 53 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=2.655 $Y=1.957
+ $X2=2.315 $Y2=1.957
r143 48 62 0.301081 $w=2.15e-07 $l=1e-07 $layer=LI1_cond $X=2.315 $Y=0.762
+ $X2=2.215 $Y2=0.762
r144 48 50 32.9652 $w=2.13e-07 $l=6.15e-07 $layer=LI1_cond $X=2.315 $Y=0.762
+ $X2=2.93 $Y2=0.762
r145 47 53 7.00737 $w=2.55e-07 $l=1.67911e-07 $layer=LI1_cond $X=2.22 $Y=1.83
+ $X2=2.315 $Y2=1.957
r146 47 65 28.8947 $w=1.88e-07 $l=4.95e-07 $layer=LI1_cond $X=2.22 $Y=1.83
+ $X2=2.22 $Y2=1.335
r147 45 80 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.995 $Y=1.16
+ $X2=2.085 $Y2=1.16
r148 45 78 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.995 $Y=1.16
+ $X2=1.765 $Y2=1.16
r149 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.995
+ $Y=1.16 $X2=1.995 $Y2=1.16
r150 41 73 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.635 $Y=1.16
+ $X2=0.795 $Y2=1.16
r151 41 70 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.635 $Y=1.16
+ $X2=0.475 $Y2=1.16
r152 40 44 46.0977 $w=3.38e-07 $l=1.36e-06 $layer=LI1_cond $X=0.635 $Y=1.165
+ $X2=1.995 $Y2=1.165
r153 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.635
+ $Y=1.16 $X2=0.635 $Y2=1.16
r154 38 65 9.46595 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=2.215 $Y=1.165
+ $X2=2.215 $Y2=1.335
r155 38 62 22.3482 $w=1.98e-07 $l=4.03e-07 $layer=LI1_cond $X=2.215 $Y=1.165
+ $X2=2.215 $Y2=0.762
r156 38 44 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.115 $Y=1.165
+ $X2=1.995 $Y2=1.165
r157 34 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.325
+ $X2=2.085 $Y2=1.16
r158 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.085 $Y=1.325
+ $X2=2.085 $Y2=1.985
r159 31 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=1.16
r160 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.765 $Y=0.995
+ $X2=1.765 $Y2=0.56
r161 27 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.325
+ $X2=1.655 $Y2=1.16
r162 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.655 $Y=1.325
+ $X2=1.655 $Y2=1.985
r163 24 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=1.16
r164 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.335 $Y=0.995
+ $X2=1.335 $Y2=0.56
r165 20 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.225 $Y=1.325
+ $X2=1.225 $Y2=1.16
r166 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.225 $Y=1.325
+ $X2=1.225 $Y2=1.985
r167 17 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=1.16
r168 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.905 $Y=0.995
+ $X2=0.905 $Y2=0.56
r169 13 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.795 $Y=1.325
+ $X2=0.795 $Y2=1.16
r170 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.795 $Y=1.325
+ $X2=0.795 $Y2=1.985
r171 10 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r172 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r173 3 69 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=4.24
+ $Y=1.485 $X2=4.38 $Y2=2.02
r174 2 67 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.485 $X2=2.75 $Y2=1.96
r175 2 56 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.485 $X2=2.75 $Y2=2.3
r176 1 50 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.235 $X2=2.93 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%B1 3 5 7 10 12 14 15 21 27
c53 12 0 1.04122e-19 $X=3.145 $Y=0.995
r54 25 27 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.145 $Y2=1.16
r55 23 25 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.965 $Y=1.16
+ $X2=2.99 $Y2=1.16
r56 22 23 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.715 $Y=1.16
+ $X2=2.965 $Y2=1.16
r57 21 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.16 $X2=2.99 $Y2=1.16
r58 20 22 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.65 $Y=1.16
+ $X2=2.715 $Y2=1.16
r59 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.16 $X2=2.65 $Y2=1.16
r60 17 20 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.535 $Y=1.16
+ $X2=2.65 $Y2=1.16
r61 15 21 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.82 $Y=1.53
+ $X2=2.82 $Y2=1.16
r62 12 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=1.16
r63 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=0.56
r64 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.325
+ $X2=2.965 $Y2=1.16
r65 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.965 $Y=1.325
+ $X2=2.965 $Y2=1.985
r66 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=0.995
+ $X2=2.715 $Y2=1.16
r67 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.715 $Y=0.995
+ $X2=2.715 $Y2=0.56
r68 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=1.325
+ $X2=2.535 $Y2=1.16
r69 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.535 $Y=1.325
+ $X2=2.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%A1 3 6 10 13 17 18 20 21 22 26 29 30 31 33
c75 17 0 3.15029e-19 $X=3.6 $Y=1.16
r76 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.16
+ $X2=5.115 $Y2=1.325
r77 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.16
+ $X2=5.115 $Y2=0.995
r78 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.16 $X2=5.115 $Y2=1.16
r79 22 33 2.72052 $w=3.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.215 $Y=1.6
+ $X2=5.215 $Y2=1.495
r80 22 33 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.215 $Y=1.47
+ $X2=5.215 $Y2=1.495
r81 22 30 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.215 $Y=1.47
+ $X2=5.215 $Y2=1.16
r82 20 22 4.7933 $w=2.1e-07 $l=1.85e-07 $layer=LI1_cond $X=5.03 $Y=1.6 $X2=5.215
+ $Y2=1.6
r83 20 21 65.7532 $w=2.08e-07 $l=1.245e-06 $layer=LI1_cond $X=5.03 $Y=1.6
+ $X2=3.785 $Y2=1.6
r84 18 27 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.622 $Y=1.16
+ $X2=3.622 $Y2=1.325
r85 18 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.622 $Y=1.16
+ $X2=3.622 $Y2=0.995
r86 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.16 $X2=3.6 $Y2=1.16
r87 15 21 7.12258 $w=2.1e-07 $l=1.98681e-07 $layer=LI1_cond $X=3.632 $Y=1.495
+ $X2=3.785 $Y2=1.6
r88 15 17 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=3.632 $Y=1.495
+ $X2=3.632 $Y2=1.16
r89 13 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.025 $Y=1.985
+ $X2=5.025 $Y2=1.325
r90 10 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.025 $Y=0.56
+ $X2=5.025 $Y2=0.995
r91 6 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.735 $Y=1.985
+ $X2=3.735 $Y2=1.325
r92 3 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.655 $Y=0.56
+ $X2=3.655 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%A2 1 3 6 8 10 13 15 21 22
c47 1 0 9.88159e-20 $X=4.165 $Y=0.995
r48 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.16 $X2=4.605 $Y2=1.16
r49 19 21 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.595 $Y=1.16
+ $X2=4.605 $Y2=1.16
r50 17 19 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.165 $Y=1.16
+ $X2=4.595 $Y2=1.16
r51 15 22 0.652406 $w=5.48e-07 $l=3e-08 $layer=LI1_cond $X=4.415 $Y=1.19
+ $X2=4.415 $Y2=1.16
r52 11 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.595 $Y=1.325
+ $X2=4.595 $Y2=1.985
r54 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.595 $Y=0.995
+ $X2=4.595 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.165 $Y=1.325
+ $X2=4.165 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.165 $Y=1.325
+ $X2=4.165 $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.165 $Y=0.995
+ $X2=4.165 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.165 $Y=0.995
+ $X2=4.165 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%VPWR 1 2 3 4 5 18 22 26 28 30 33 34 36 37 39
+ 40 41 57 68 71 74
c90 39 0 1.69833e-19 $X=2.135 $Y=2.72
c91 4 0 1.12091e-19 $X=3.04 $Y=1.485
r92 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r93 70 71 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=2.54
+ $X2=3.685 $Y2=2.54
r94 66 70 1.57973 $w=5.28e-07 $l=7e-08 $layer=LI1_cond $X=3.45 $Y=2.54 $X2=3.52
+ $Y2=2.54
r95 66 68 15.7976 $w=5.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.45 $Y=2.54
+ $X2=3.015 $Y2=2.54
r96 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r97 64 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r99 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r100 61 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 60 71 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=3.685 $Y2=2.72
r103 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 57 73 5.10352 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=5.297 $Y2=2.72
r105 57 63 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.075 $Y=2.72
+ $X2=4.83 $Y2=2.72
r106 56 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 55 68 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=3.015 $Y2=2.72
r108 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 52 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r110 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r113 41 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 41 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r115 39 51 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.07 $Y2=2.72
r116 39 40 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.31 $Y2=2.72
r117 38 55 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.99 $Y2=2.72
r118 38 40 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.31 $Y2=2.72
r119 36 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=1.44 $Y2=2.72
r121 35 51 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=2.07 $Y2=2.72
r122 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.44 $Y2=2.72
r123 33 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.58 $Y2=2.72
r125 32 48 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.745 $Y=2.72
+ $X2=1.15 $Y2=2.72
r126 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=2.72
+ $X2=0.58 $Y2=2.72
r127 28 73 2.91958 $w=3.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.255 $Y=2.635
+ $X2=5.297 $Y2=2.72
r128 28 30 19.6876 $w=3.58e-07 $l=6.15e-07 $layer=LI1_cond $X=5.255 $Y=2.635
+ $X2=5.255 $Y2=2.02
r129 24 40 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.635
+ $X2=2.31 $Y2=2.72
r130 24 26 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.31 $Y=2.635
+ $X2=2.31 $Y2=2.34
r131 20 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=2.635
+ $X2=1.44 $Y2=2.72
r132 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.44 $Y=2.635
+ $X2=1.44 $Y2=1.955
r133 16 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.58 $Y=2.635
+ $X2=0.58 $Y2=2.72
r134 16 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.58 $Y=2.635
+ $X2=0.58 $Y2=1.955
r135 5 30 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=5.1
+ $Y=1.485 $X2=5.24 $Y2=2.02
r136 4 70 300 $w=1.7e-07 $l=1.08886e-06 $layer=licon1_PDIFF $count=2 $X=3.04
+ $Y=1.485 $X2=3.52 $Y2=2.36
r137 3 26 600 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=1.485 $X2=2.32 $Y2=2.34
r138 2 22 300 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=2 $X=1.3
+ $Y=1.485 $X2=1.44 $Y2=1.955
r139 1 18 300 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_PDIFF $count=2 $X=0.455
+ $Y=1.485 $X2=0.58 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%X 1 2 3 4 13 14 17 19 23 25 29 33 34 35 39 41
c51 39 0 1.01803e-19 $X=0.205 $Y=0.805
r52 39 41 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.205 $Y=0.805
+ $X2=0.205 $Y2=0.85
r53 35 39 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.205 $Y=0.72
+ $X2=0.205 $Y2=0.805
r54 35 41 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=0.205 $Y=0.87
+ $X2=0.205 $Y2=0.85
r55 33 35 14.9587 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.32 $Y2=0.72
r56 31 35 33.0701 $w=2.28e-07 $l=6.6e-07 $layer=LI1_cond $X=0.205 $Y=1.53
+ $X2=0.205 $Y2=0.87
r57 27 29 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.865 $Y=1.7
+ $X2=1.865 $Y2=1.84
r58 26 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.105 $Y=1.615
+ $X2=1.01 $Y2=1.615
r59 25 27 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.775 $Y=1.615
+ $X2=1.865 $Y2=1.7
r60 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.775 $Y=1.615
+ $X2=1.105 $Y2=1.615
r61 21 34 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=1.7 $X2=1.01
+ $Y2=1.615
r62 21 23 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=1.01 $Y=1.7 $X2=1.01
+ $Y2=1.84
r63 17 33 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.69 $Y=0.71
+ $X2=0.595 $Y2=0.71
r64 17 19 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=0.69 $Y=0.71 $X2=1.55
+ $Y2=0.71
r65 14 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.32 $Y=1.615
+ $X2=0.205 $Y2=1.53
r66 13 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.915 $Y=1.615
+ $X2=1.01 $Y2=1.615
r67 13 14 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.915 $Y=1.615
+ $X2=0.32 $Y2=1.615
r68 4 29 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=1.485 $X2=1.87 $Y2=1.84
r69 3 23 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=0.87
+ $Y=1.485 $X2=1.01 $Y2=1.84
r70 2 19 182 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.71
r71 1 17 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 60 61 67 70 73 76
c92 16 0 1.01803e-19 $X=0.26 $Y=0.085
r93 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r94 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r95 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r96 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r97 61 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r98 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r99 58 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=4.81
+ $Y2=0
r100 58 60 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=5.29 $Y2=0
r101 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r102 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r103 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r104 54 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=3.945
+ $Y2=0
r105 54 56 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=4.37 $Y2=0
r106 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=0 $X2=4.81
+ $Y2=0
r107 53 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=4.37 $Y2=0
r108 52 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r109 52 71 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.07 $Y2=0
r110 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r111 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r112 49 51 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=2.145 $Y=0
+ $X2=3.45 $Y2=0
r113 48 73 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=3.945
+ $Y2=0
r114 48 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=3.45 $Y2=0
r115 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r116 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r117 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r118 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r119 44 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.61 $Y2=0
r120 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r121 43 46 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.815 $Y=0
+ $X2=1.61 $Y2=0
r122 42 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r123 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r124 39 64 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r125 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r126 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r127 38 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.69 $Y2=0
r128 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r129 36 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r130 32 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0
r131 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0.36
r132 28 73 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0
r133 28 30 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=3.945 $Y=0.085
+ $X2=3.945 $Y2=0.36
r134 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r135 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.38
r136 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r137 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r138 16 64 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r139 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r140 5 34 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.235 $X2=4.81 $Y2=0.36
r141 4 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.73
+ $Y=0.235 $X2=3.94 $Y2=0.36
r142 3 26 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.38
r143 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.36
r144 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_4%A_475_47# 1 2 3 4 13 21 24
r39 26 27 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.44 $Y=0.37
+ $X2=3.44 $Y2=0.7
r40 24 26 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.44 $Y=0.36 $X2=3.44
+ $Y2=0.37
r41 19 21 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=4.38 $Y=0.7 $X2=5.24
+ $Y2=0.7
r42 17 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=0.7
+ $X2=3.44 $Y2=0.7
r43 17 19 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.605 $Y=0.7
+ $X2=4.38 $Y2=0.7
r44 13 26 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=0.37
+ $X2=3.44 $Y2=0.37
r45 13 15 38.8323 $w=2.28e-07 $l=7.75e-07 $layer=LI1_cond $X=3.275 $Y=0.37
+ $X2=2.5 $Y2=0.37
r46 4 21 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=5.1
+ $Y=0.235 $X2=5.24 $Y2=0.7
r47 3 19 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.24
+ $Y=0.235 $X2=4.38 $Y2=0.7
r48 2 24 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=3.22
+ $Y=0.235 $X2=3.44 $Y2=0.36
r49 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.5 $Y2=0.38
.ends


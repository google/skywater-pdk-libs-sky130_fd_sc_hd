* NGSPICE file created from sky130_fd_sc_hd__or2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
M1000 X a_35_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.4e+11p pd=5.08e+06u as=9.05e+11p ps=7.81e+06u
M1001 X a_35_297# VGND VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=7.4425e+11p ps=7.49e+06u
M1002 VPWR A a_121_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1003 VPWR a_35_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_35_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_121_297# B a_35_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1007 X a_35_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_35_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1010 VPWR a_35_297# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_35_297# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a22o_2.pex.spice
* Created: Thu Aug 27 14:02:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22O_2%B2 3 6 8 11 12 13
c27 6 0 1.14647e-19 $X=0.47 $Y=1.985
r28 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r29 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r30 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r31 8 12 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.41 $Y2=1.175
r32 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r33 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%B1 3 6 8 9 13 15
r40 17 23 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=1.13 $Y=1.075
+ $X2=1.13 $Y2=1.18
r41 14 23 10.5628 $w=2.08e-07 $l=2e-07 $layer=LI1_cond $X=0.93 $Y=1.18 $X2=1.13
+ $Y2=1.18
r42 13 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=1.325
r43 13 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=0.995
r44 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r45 9 23 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.13 $Y2=1.18
r46 8 17 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.13 $Y=0.85
+ $X2=1.13 $Y2=1.075
r47 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r48 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.56 $X2=0.85
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%A1 3 6 8 9 13 15
r38 17 21 0.716491 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=1.615 $Y=1.075
+ $X2=1.615 $Y2=1.18
r39 13 16 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.722 $Y=1.16
+ $X2=1.722 $Y2=1.325
r40 13 15 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.722 $Y=1.16
+ $X2=1.722 $Y2=0.995
r41 9 21 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=1.635 $Y=1.18 $X2=1.615
+ $Y2=1.18
r42 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r43 8 17 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.615 $Y=0.85
+ $X2=1.615 $Y2=1.075
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.985
+ $X2=1.83 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.56 $X2=1.83
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%A2 3 6 8 11 12 13
r37 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=1.325
r38 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=0.995
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.16 $X2=2.25 $Y2=1.16
r40 8 12 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=2.095 $Y=1.175
+ $X2=2.25 $Y2=1.175
r41 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.31 $Y=1.985
+ $X2=2.31 $Y2=1.325
r42 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.31 $Y=0.56 $X2=2.31
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%A_27_297# 1 2 3 4 13 15 18 20 22 25 28 30 31
+ 32 35 42 43 44 48 53 54 59
c123 59 0 2.21533e-19 $X=3.195 $Y=1.16
c124 53 0 1.14647e-19 $X=1.1 $Y=2.34
r125 58 59 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.775 $Y=1.16
+ $X2=3.195 $Y2=1.16
r126 53 54 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=2.36
+ $X2=0.935 $Y2=2.36
r127 49 58 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=2.775 $Y2=1.16
r128 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.73
+ $Y=1.16 $X2=2.73 $Y2=1.16
r129 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.73 $Y=1.455
+ $X2=2.73 $Y2=1.16
r130 45 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.73 $Y=0.905
+ $X2=2.73 $Y2=1.16
r131 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=0.82
+ $X2=2.73 $Y2=0.905
r132 43 44 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.645 $Y=0.82
+ $X2=2.145 $Y2=0.82
r133 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.735
+ $X2=2.145 $Y2=0.82
r134 41 42 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.06 $Y=0.505
+ $X2=2.06 $Y2=0.735
r135 37 40 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.06 $Y=0.38
+ $X2=1.62 $Y2=0.38
r136 35 41 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.975 $Y=0.38
+ $X2=2.06 $Y2=0.505
r137 35 40 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=1.975 $Y=0.38
+ $X2=1.62 $Y2=0.38
r138 34 51 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.26 $Y2=2.38
r139 34 54 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.935 $Y2=2.38
r140 31 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=1.54
+ $X2=2.73 $Y2=1.455
r141 31 32 144.834 $w=1.68e-07 $l=2.22e-06 $layer=LI1_cond $X=2.645 $Y=1.54
+ $X2=0.425 $Y2=1.54
r142 28 51 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=2.38
r143 28 30 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.66
r144 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.425 $Y2=1.54
r145 27 30 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.66
r146 23 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.16
r147 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.985
r148 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=0.995
+ $X2=3.195 $Y2=1.16
r149 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.195 $Y=0.995
+ $X2=3.195 $Y2=0.56
r150 16 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.325
+ $X2=2.775 $Y2=1.16
r151 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.775 $Y=1.325
+ $X2=2.775 $Y2=1.985
r152 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=0.995
+ $X2=2.775 $Y2=1.16
r153 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.775 $Y=0.995
+ $X2=2.775 $Y2=0.56
r154 4 53 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2.34
r155 3 51 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r156 3 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r157 2 40 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.42
r158 1 37 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.235 $X2=1.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%A_109_297# 1 2 7 9 11 16
r23 14 16 5.94149 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.68 $Y=1.96
+ $X2=0.825 $Y2=1.96
r24 9 18 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.105 $Y2=1.915
r25 9 11 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.105 $Y=2.035
+ $X2=2.105 $Y2=2.3
r26 7 18 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=1.98 $Y=1.915
+ $X2=2.105 $Y2=1.915
r27 7 16 55.4613 $w=2.38e-07 $l=1.155e-06 $layer=LI1_cond $X=1.98 $Y=1.915
+ $X2=0.825 $Y2=1.915
r28 2 18 600 $w=1.7e-07 $l=5.39096e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.065 $Y2=1.95
r29 2 11 600 $w=1.7e-07 $l=8.91417e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.485 $X2=2.065 $Y2=2.3
r30 1 14 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%VPWR 1 2 3 12 16 18 20 24 26 34 39 45 48 52
c55 16 0 1.18411e-19 $X=2.565 $Y=1.96
r56 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 43 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=2.72
+ $X2=2.565 $Y2=2.72
r63 40 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.73 $Y=2.72
+ $X2=2.99 $Y2=2.72
r64 39 51 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.505 $Y2=2.72
r65 39 42 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=2.99 $Y2=2.72
r66 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r67 38 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 35 45 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=1.632 $Y2=2.72
r70 35 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=2.07 $Y2=2.72
r71 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=2.72
+ $X2=2.565 $Y2=2.72
r72 34 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.4 $Y=2.72 $X2=2.07
+ $Y2=2.72
r73 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 28 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 26 45 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.632 $Y2=2.72
r77 26 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 24 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 24 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 20 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.415 $Y=1.63
+ $X2=3.415 $Y2=2.31
r81 18 51 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.415 $Y=2.635
+ $X2=3.505 $Y2=2.72
r82 18 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.415 $Y=2.635
+ $X2=3.415 $Y2=2.31
r83 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=2.635
+ $X2=2.565 $Y2=2.72
r84 14 16 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.565 $Y=2.635
+ $X2=2.565 $Y2=1.96
r85 10 45 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.72
r86 10 12 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.632 $Y=2.635
+ $X2=1.632 $Y2=2.3
r87 3 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.485 $X2=3.415 $Y2=2.31
r88 3 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.485 $X2=3.415 $Y2=1.63
r89 2 16 300 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=2 $X=2.385
+ $Y=1.485 $X2=2.565 $Y2=1.96
r90 1 12 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%X 1 2 10 13 14 30
r21 19 30 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.03 $Y=1.915
+ $X2=3.03 $Y2=1.87
r22 13 30 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.03 $Y=1.85 $X2=3.03
+ $Y2=1.87
r23 13 14 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.03 $Y=1.935
+ $X2=3.03 $Y2=2.21
r24 13 19 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.03 $Y=1.935
+ $X2=3.03 $Y2=1.915
r25 11 13 50.6043 $w=2.78e-07 $l=1.2e-06 $layer=LI1_cond $X=3.075 $Y=0.585
+ $X2=3.075 $Y2=1.785
r26 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=0.42
+ $X2=3.075 $Y2=0.585
r27 8 10 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.985 $Y=0.42 $X2=3.075
+ $Y2=0.42
r28 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=1.485 $X2=2.985 $Y2=1.96
r29 1 8 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.85
+ $Y=0.235 $X2=2.985 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_2%VGND 1 2 3 10 12 16 18 20 22 24 32 41 45
c49 16 0 1.03121e-19 $X=2.52 $Y=0.4
r50 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r51 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 36 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r53 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r54 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 33 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.52
+ $Y2=0
r56 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.99
+ $Y2=0
r57 32 44 3.40825 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.505
+ $Y2=0
r58 32 35 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=2.99
+ $Y2=0
r59 31 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r60 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r61 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r62 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r63 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r64 25 38 5.92045 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.272
+ $Y2=0
r65 25 27 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.69
+ $Y2=0
r66 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.52
+ $Y2=0
r67 24 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.07
+ $Y2=0
r68 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 18 44 3.40825 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.505 $Y2=0
r71 18 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0.4
r72 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.52 $Y2=0
r73 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.52 $Y2=0.4
r74 10 38 2.88432 $w=4.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.272 $Y2=0
r75 10 12 8.37255 $w=4.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.32 $Y2=0.4
r76 3 20 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.27
+ $Y=0.235 $X2=3.415 $Y2=0.4
r77 2 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.235 $X2=2.52 $Y2=0.4
r78 1 12 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


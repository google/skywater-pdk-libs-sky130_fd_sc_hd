* File: sky130_fd_sc_hd__o31ai_2.pex.spice
* Created: Thu Aug 27 14:40:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31AI_2%A1 3 7 11 15 17 18 19 31
c52 31 0 1.58465e-19 $X=0.91 $Y=1.16
r53 29 31 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.82 $Y=1.16 $X2=0.91
+ $Y2=1.16
r54 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.82
+ $Y=1.16 $X2=0.82 $Y2=1.16
r55 27 29 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.82 $Y2=1.16
r56 24 27 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=0.48 $Y=1.16 $X2=0.49
+ $Y2=1.16
r57 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.48
+ $Y=1.16 $X2=0.48 $Y2=1.16
r58 19 30 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=0.82 $Y2=1.19
r59 18 30 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.19
+ $X2=0.82 $Y2=1.19
r60 18 25 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.695 $Y=1.19
+ $X2=0.48 $Y2=1.19
r61 17 25 10.4574 $w=2.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.235 $Y=1.19
+ $X2=0.48 $Y2=1.19
r62 13 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=1.16
r63 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.91 $Y=1.295
+ $X2=0.91 $Y2=1.985
r64 9 31 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.91 $Y=1.025
+ $X2=0.91 $Y2=1.16
r65 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.91 $Y=1.025
+ $X2=0.91 $Y2=0.56
r66 5 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.16
r67 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.49 $Y=1.295 $X2=0.49
+ $Y2=1.985
r68 1 27 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=1.16
r69 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%A2 3 7 11 15 17 18 30
c46 18 0 2.90077e-19 $X=2.075 $Y=1.19
c47 11 0 1.01157e-19 $X=1.75 $Y=1.985
r48 28 30 38.8804 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=1.915 $Y=1.16
+ $X2=2.09 $Y2=1.16
r49 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.16 $X2=1.915 $Y2=1.16
r50 26 28 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.16
+ $X2=1.915 $Y2=1.16
r51 24 26 38.8804 $w=2.7e-07 $l=1.75e-07 $layer=POLY_cond $X=1.575 $Y=1.16
+ $X2=1.75 $Y2=1.16
r52 21 24 54.4326 $w=2.7e-07 $l=2.45e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.575 $Y2=1.16
r53 18 29 6.82929 $w=2.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.075 $Y=1.19
+ $X2=1.915 $Y2=1.19
r54 17 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.575 $Y=1.19
+ $X2=1.915 $Y2=1.19
r55 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.16 $X2=1.575 $Y2=1.16
r56 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.09 $Y=1.025
+ $X2=2.09 $Y2=1.16
r57 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.09 $Y=1.025
+ $X2=2.09 $Y2=0.56
r58 9 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.75 $Y=1.295
+ $X2=1.75 $Y2=1.16
r59 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.75 $Y=1.295
+ $X2=1.75 $Y2=1.985
r60 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.33 $Y=1.295
+ $X2=1.33 $Y2=1.16
r61 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.33 $Y=1.295 $X2=1.33
+ $Y2=1.985
r62 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.33 $Y=1.025
+ $X2=1.33 $Y2=1.16
r63 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.33 $Y=1.025
+ $X2=1.33 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%A3 3 7 11 15 17 18 30
c52 18 0 1.01157e-19 $X=2.995 $Y=1.19
c53 7 0 1.31612e-19 $X=2.71 $Y=1.985
r54 28 30 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3.04 $Y=1.16 $X2=3.13
+ $Y2=1.16
r55 26 28 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.71 $Y=1.16
+ $X2=3.04 $Y2=1.16
r56 24 26 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=2.7 $Y=1.16 $X2=2.71
+ $Y2=1.16
r57 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.16 $X2=2.7 $Y2=1.16
r58 21 24 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=2.63 $Y=1.16 $X2=2.7
+ $Y2=1.16
r59 18 25 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.995 $Y=1.19
+ $X2=2.7 $Y2=1.19
r60 18 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.16 $X2=3.04 $Y2=1.16
r61 17 25 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=1.19
+ $X2=2.7 $Y2=1.19
r62 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.16
r63 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.985
r64 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=1.16
r65 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.13 $Y=1.025
+ $X2=3.13 $Y2=0.56
r66 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.71 $Y=1.295
+ $X2=2.71 $Y2=1.16
r67 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.71 $Y=1.295 $X2=2.71
+ $Y2=1.985
r68 1 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.63 $Y=1.025
+ $X2=2.63 $Y2=1.16
r69 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.63 $Y=1.025
+ $X2=2.63 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%B1 1 3 6 8 10 12 15 17 18 19 24
r49 22 24 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.09 $Y=1.16
+ $X2=4.36 $Y2=1.16
r50 18 19 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=4.345 $Y=1.16
+ $X2=4.345 $Y2=0.85
r51 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.16 $X2=4.36 $Y2=1.16
r52 13 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=1.325
+ $X2=4.09 $Y2=1.16
r53 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.09 $Y=1.325
+ $X2=4.09 $Y2=1.985
r54 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=1.16
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=0.56
r56 9 17 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.625 $Y=1.16
+ $X2=3.55 $Y2=1.16
r57 8 22 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.015 $Y=1.16
+ $X2=4.09 $Y2=1.16
r58 8 9 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.015 $Y=1.16
+ $X2=3.625 $Y2=1.16
r59 4 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.325
+ $X2=3.55 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.55 $Y=1.325 $X2=3.55
+ $Y2=1.985
r61 1 17 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=0.995
+ $X2=3.55 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.55 $Y=0.995 $X2=3.55
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%A_27_297# 1 2 3 12 16 17 20 24 28 30
r44 26 28 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.68
r45 25 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=1.58
+ $X2=1.12 $Y2=1.58
r46 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=1.58
+ $X2=1.96 $Y2=1.665
r47 24 25 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.795 $Y=1.58
+ $X2=1.285 $Y2=1.58
r48 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.12 $Y=1.68
+ $X2=1.12 $Y2=2.36
r49 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.58
r50 18 20 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.68
r51 16 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=1.58
+ $X2=1.12 $Y2=1.58
r52 16 17 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.955 $Y=1.58
+ $X2=0.445 $Y2=1.58
r53 12 14 22.075 $w=3.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.267 $Y=1.68
+ $X2=0.267 $Y2=2.36
r54 10 17 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=1.665
+ $X2=0.445 $Y2=1.58
r55 10 12 0.486948 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=0.267 $Y=1.665
+ $X2=0.267 $Y2=1.68
r56 3 28 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.68
r57 2 22 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.36
r58 2 20 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.68
r59 1 14 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.36
r60 1 12 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%VPWR 1 2 11 15 17 19 29 30 33 36 39
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r56 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r57 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=3.84 $Y2=2.72
r58 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=4.37 $Y2=2.72
r59 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 23 26 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 22 25 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 20 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=2.72 $X2=0.7
+ $Y2=2.72
r66 20 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.84 $Y2=2.72
r68 19 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 17 34 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 17 39 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.84 $Y2=2.72
r72 13 15 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.84 $Y2=2.02
r73 9 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r74 9 11 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2
r75 2 15 300 $w=1.7e-07 $l=6.33443e-07 $layer=licon1_PDIFF $count=2 $X=3.625
+ $Y=1.485 $X2=3.84 $Y2=2.02
r76 1 11 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%A_281_297# 1 2 9 11 12 15
r19 13 15 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.92 $Y=2.295
+ $X2=2.92 $Y2=2.135
r20 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.835 $Y=2.38
+ $X2=2.92 $Y2=2.295
r21 11 12 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.835 $Y=2.38
+ $X2=1.625 $Y2=2.38
r22 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.54 $Y=2.295
+ $X2=1.625 $Y2=2.38
r23 7 9 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=2.295 $X2=1.54
+ $Y2=2.135
r24 2 15 600 $w=1.7e-07 $l=7.14318e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.485 $X2=2.92 $Y2=2.135
r25 1 9 600 $w=1.7e-07 $l=7.14318e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%Y 1 2 3 4 13 14 17 22 23 24 25 26 27 36 42
+ 49 51
r56 49 51 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=4.345 $Y=1.665
+ $X2=4.345 $Y2=1.765
r57 26 27 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=4.345 $Y=1.87
+ $X2=4.345 $Y2=2.21
r58 26 51 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=4.345 $Y=1.87
+ $X2=4.345 $Y2=1.765
r59 25 49 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.915 $Y=1.58
+ $X2=4.345 $Y2=1.58
r60 25 40 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.915 $Y=1.58
+ $X2=3.84 $Y2=1.58
r61 25 40 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.84 $Y=1.47
+ $X2=3.84 $Y2=1.495
r62 24 25 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.84 $Y=1.19 $X2=3.84
+ $Y2=1.47
r63 23 24 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.84 $Y=0.85
+ $X2=3.84 $Y2=1.19
r64 23 42 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.84 $Y=0.85
+ $X2=3.84 $Y2=0.755
r65 22 36 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.5 $Y=1.87 $X2=2.5
+ $Y2=1.68
r66 21 36 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.5 $Y=1.665
+ $X2=2.5 $Y2=1.68
r67 17 19 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.34 $Y=1.68
+ $X2=3.34 $Y2=2.36
r68 15 40 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.34 $Y=1.58 $X2=3.84
+ $Y2=1.58
r69 15 17 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.34 $Y=1.665
+ $X2=3.34 $Y2=1.68
r70 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.665 $Y=1.58
+ $X2=2.5 $Y2=1.665
r71 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=1.58
+ $X2=3.34 $Y2=1.58
r72 13 14 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.175 $Y=1.58
+ $X2=2.665 $Y2=1.58
r73 4 51 300 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=2 $X=4.165
+ $Y=1.485 $X2=4.3 $Y2=1.765
r74 3 19 400 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.485 $X2=3.34 $Y2=2.36
r75 3 17 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.485 $X2=3.34 $Y2=1.68
r76 2 36 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.5 $Y2=1.68
r77 1 42 182 $w=1.7e-07 $l=6.18223e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.84 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 32 34
+ 35 36 38 39 42
r81 42 45 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=4.345 $Y=0.34
+ $X2=4.345 $Y2=0.42
r82 37 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=0.34
+ $X2=3.34 $Y2=0.34
r83 36 42 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.175 $Y=0.34
+ $X2=4.345 $Y2=0.34
r84 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.175 $Y=0.34
+ $X2=3.505 $Y2=0.34
r85 34 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=0.425 $X2=3.34
+ $Y2=0.34
r86 34 35 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.34 $Y=0.425
+ $X2=3.34 $Y2=0.715
r87 33 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0.8
+ $X2=2.34 $Y2=0.8
r88 32 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.175 $Y=0.8
+ $X2=3.34 $Y2=0.715
r89 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.175 $Y=0.8
+ $X2=2.505 $Y2=0.8
r90 28 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.715
+ $X2=2.34 $Y2=0.8
r91 28 30 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.34 $Y=0.715
+ $X2=2.34 $Y2=0.36
r92 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0.8
+ $X2=1.12 $Y2=0.8
r93 26 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=0.8
+ $X2=2.34 $Y2=0.8
r94 26 27 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.175 $Y=0.8
+ $X2=1.285 $Y2=0.8
r95 22 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.12 $Y2=0.8
r96 22 24 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.12 $Y=0.715
+ $X2=1.12 $Y2=0.36
r97 20 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0.8
+ $X2=1.12 $Y2=0.8
r98 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.955 $Y=0.8
+ $X2=0.445 $Y2=0.8
r99 16 21 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.445 $Y2=0.8
r100 16 18 11.5244 $w=3.53e-07 $l=3.55e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.267 $Y2=0.36
r101 5 45 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.165
+ $Y=0.235 $X2=4.3 $Y2=0.42
r102 4 41 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.205
+ $Y=0.235 $X2=3.34 $Y2=0.36
r103 3 30 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=2.165
+ $Y=0.235 $X2=2.34 $Y2=0.36
r104 2 24 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.36
r105 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31AI_2%VGND 1 2 3 14 18 20 22 27 34 35 38 42 48 51
r65 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r66 42 45 8.91196 $w=5.08e-07 $l=3.8e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.71
+ $Y2=0.38
r67 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r68 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 35 49 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=2.99
+ $Y2=0
r70 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r71 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=2.84
+ $Y2=0
r72 32 34 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=3.005 $Y=0
+ $X2=4.37 $Y2=0
r73 31 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r74 31 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r75 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r76 28 42 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.71
+ $Y2=0
r77 28 30 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.53
+ $Y2=0
r78 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.84
+ $Y2=0
r79 27 30 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.53
+ $Y2=0
r80 26 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r81 26 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r82 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r83 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r84 23 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.15
+ $Y2=0
r85 22 42 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.71
+ $Y2=0
r86 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.15
+ $Y2=0
r87 20 39 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r88 20 51 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r89 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r90 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.36
r91 12 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r92 12 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.38
r93 3 18 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.235 $X2=2.84 $Y2=0.36
r94 2 45 91 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.88 $Y2=0.38
r95 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__clkinvlp_4.pxi.spice
* Created: Thu Aug 27 14:13:05 2020
* 
x_PM_SKY130_FD_SC_HD__CLKINVLP_4%A N_A_M1002_g N_A_M1001_g N_A_M1000_g
+ N_A_M1004_g N_A_M1006_g N_A_M1005_g N_A_M1003_g N_A_M1007_g A A N_A_c_36_n
+ PM_SKY130_FD_SC_HD__CLKINVLP_4%A
x_PM_SKY130_FD_SC_HD__CLKINVLP_4%VPWR N_VPWR_M1001_d N_VPWR_M1004_d
+ N_VPWR_M1007_d N_VPWR_c_101_n N_VPWR_c_102_n N_VPWR_c_103_n N_VPWR_c_104_n
+ N_VPWR_c_105_n N_VPWR_c_106_n N_VPWR_c_107_n VPWR N_VPWR_c_108_n
+ N_VPWR_c_100_n PM_SKY130_FD_SC_HD__CLKINVLP_4%VPWR
x_PM_SKY130_FD_SC_HD__CLKINVLP_4%Y N_Y_M1000_s N_Y_M1001_s N_Y_M1005_s
+ N_Y_c_141_n N_Y_c_142_n Y Y Y Y Y Y N_Y_c_158_n
+ PM_SKY130_FD_SC_HD__CLKINVLP_4%Y
x_PM_SKY130_FD_SC_HD__CLKINVLP_4%VGND N_VGND_M1002_d N_VGND_M1003_d
+ N_VGND_c_180_n N_VGND_c_181_n N_VGND_c_182_n N_VGND_c_183_n N_VGND_c_184_n
+ VGND N_VGND_c_185_n N_VGND_c_186_n PM_SKY130_FD_SC_HD__CLKINVLP_4%VGND
cc_1 VNB N_A_M1002_g 0.024296f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.51
cc_2 VNB N_A_M1000_g 0.018421f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=0.51
cc_3 VNB N_A_M1006_g 0.0202106f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.51
cc_4 VNB N_A_M1003_g 0.0282192f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=0.51
cc_5 VNB A 0.0216425f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_36_n 0.129869f $X=-0.19 $Y=-0.24 $X2=2.115 $Y2=1.16
cc_7 VNB N_VPWR_c_100_n 0.117919f $X=-0.19 $Y=-0.24 $X2=1.585 $Y2=1.16
cc_8 VNB Y 0.00353344f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.51
cc_9 VNB N_VGND_c_180_n 0.0103065f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.985
cc_10 VNB N_VGND_c_181_n 0.0162274f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=0.995
cc_11 VNB N_VGND_c_182_n 0.023902f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.325
cc_12 VNB N_VGND_c_183_n 0.0315614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_184_n 0.00513431f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.995
cc_14 VNB N_VGND_c_185_n 0.0261689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_186_n 0.187921f $X=-0.19 $Y=-0.24 $X2=2.115 $Y2=1.325
cc_16 VPB N_A_M1001_g 0.0314207f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.985
cc_17 VPB N_A_M1004_g 0.0242324f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.985
cc_18 VPB N_A_M1005_g 0.0242324f $X=-0.19 $Y=1.305 $X2=1.585 $Y2=1.985
cc_19 VPB N_A_M1007_g 0.0309724f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.985
cc_20 VPB A 0.0039889f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_21 VPB N_A_c_36_n 0.0223145f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.16
cc_22 VPB N_VPWR_c_101_n 0.0103398f $X=-0.19 $Y=1.305 $X2=0.835 $Y2=0.51
cc_23 VPB N_VPWR_c_102_n 0.0413665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_103_n 0.00278574f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.51
cc_25 VPB N_VPWR_c_104_n 0.0141676f $X=-0.19 $Y=1.305 $X2=1.585 $Y2=1.985
cc_26 VPB N_VPWR_c_105_n 0.0546532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_106_n 0.0175811f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.325
cc_28 VPB N_VPWR_c_107_n 0.00436868f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.985
cc_29 VPB N_VPWR_c_108_n 0.0178633f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_30 VPB N_VPWR_c_100_n 0.0479044f $X=-0.19 $Y=1.305 $X2=1.585 $Y2=1.16
cc_31 N_A_M1001_g N_VPWR_c_102_n 0.0219215f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_32 N_A_M1004_g N_VPWR_c_102_n 8.98363e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_33 A N_VPWR_c_102_n 0.025856f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_34 N_A_c_36_n N_VPWR_c_102_n 0.00200382f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_VPWR_c_103_n 0.00116019f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_M1004_g N_VPWR_c_103_n 0.0227105f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_37 N_A_M1005_g N_VPWR_c_103_n 0.0227105f $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_M1007_g N_VPWR_c_103_n 0.00116019f $X=2.115 $Y=1.985 $X2=0 $Y2=0
cc_39 N_A_c_36_n N_VPWR_c_103_n 0.00282284f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_40 N_A_M1005_g N_VPWR_c_105_n 0.00116019f $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_41 N_A_M1007_g N_VPWR_c_105_n 0.0247483f $X=2.115 $Y=1.985 $X2=0 $Y2=0
cc_42 N_A_M1001_g N_VPWR_c_106_n 0.00794322f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_43 N_A_M1004_g N_VPWR_c_106_n 0.00839865f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_44 N_A_M1005_g N_VPWR_c_108_n 0.00839865f $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A_M1007_g N_VPWR_c_108_n 0.00839865f $X=2.115 $Y=1.985 $X2=0 $Y2=0
cc_46 N_A_M1001_g N_VPWR_c_100_n 0.0124079f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_47 N_A_M1004_g N_VPWR_c_100_n 0.0135174f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_48 N_A_M1005_g N_VPWR_c_100_n 0.0135174f $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_49 N_A_M1007_g N_VPWR_c_100_n 0.0135174f $X=2.115 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_c_36_n N_Y_c_141_n 0.0915058f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_M1004_g N_Y_c_142_n 8.59864e-19 $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A_M1005_g N_Y_c_142_n 0.0216624f $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_53 N_A_M1007_g N_Y_c_142_n 0.0257966f $X=2.115 $Y=1.985 $X2=0 $Y2=0
cc_54 N_A_c_36_n N_Y_c_142_n 0.00597104f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_M1002_g Y 0.00174791f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_56 N_A_M1000_g Y 0.00861319f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_57 N_A_M1006_g Y 0.00494149f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_58 A Y 0.0196729f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_59 N_A_c_36_n Y 0.00243632f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_60 A Y 0.0223993f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_61 N_A_c_36_n Y 0.0135506f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_M1001_g Y 0.0289365f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_63 N_A_M1004_g Y 0.0217433f $X=1.055 $Y=1.985 $X2=0 $Y2=0
cc_64 N_A_M1005_g Y 8.58618e-19 $X=1.585 $Y=1.985 $X2=0 $Y2=0
cc_65 A Y 0.00223357f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_66 N_A_c_36_n Y 0.00530034f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_Y_c_158_n 0.0107043f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_Y_c_158_n 0.00788413f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_Y_c_158_n 0.00114752f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_70 N_A_c_36_n N_Y_c_158_n 0.00254697f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_71 A N_VGND_M1002_d 0.00242856f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_72 N_A_M1002_g N_VGND_c_181_n 0.00973267f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_VGND_c_181_n 0.00146442f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_74 A N_VGND_c_181_n 0.0232502f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_c_36_n N_VGND_c_181_n 0.00113149f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_VGND_c_182_n 0.0028519f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_VGND_c_182_n 0.0180923f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_78 N_A_c_36_n N_VGND_c_182_n 0.00752897f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_VGND_c_183_n 0.00486043f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_VGND_c_183_n 0.00357877f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_81 N_A_M1006_g N_VGND_c_183_n 0.00547467f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_VGND_c_183_n 0.00486043f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_VGND_c_186_n 0.00809891f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_VGND_c_186_n 0.00511556f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_85 N_A_M1006_g N_VGND_c_186_n 0.00973853f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VGND_c_186_n 0.00809891f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_87 A N_VGND_c_186_n 0.00163141f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_88 N_VPWR_c_100_n N_Y_M1001_s 0.00223231f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_89 N_VPWR_c_100_n N_Y_M1005_s 0.00223231f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_90 N_VPWR_c_103_n N_Y_c_141_n 0.0271408f $X=1.32 $Y=1.63 $X2=0 $Y2=0
cc_91 N_VPWR_c_103_n N_Y_c_142_n 0.0658907f $X=1.32 $Y=1.63 $X2=0 $Y2=0
cc_92 N_VPWR_c_105_n N_Y_c_142_n 0.0658907f $X=2.38 $Y=1.63 $X2=0 $Y2=0
cc_93 N_VPWR_c_108_n N_Y_c_142_n 0.0189253f $X=2.215 $Y=2.72 $X2=0 $Y2=0
cc_94 N_VPWR_c_100_n N_Y_c_142_n 0.0122674f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_95 N_VPWR_c_102_n Y 0.0732814f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_96 N_VPWR_c_103_n Y 0.0663324f $X=1.32 $Y=1.63 $X2=0 $Y2=0
cc_97 N_VPWR_c_106_n Y 0.0209707f $X=1.155 $Y=2.72 $X2=0 $Y2=0
cc_98 N_VPWR_c_100_n Y 0.0132856f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_99 N_Y_c_141_n N_VGND_c_182_n 0.0198945f $X=1.685 $Y=1.155 $X2=0 $Y2=0
cc_100 N_Y_c_158_n N_VGND_c_182_n 0.0149002f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_101 N_Y_c_158_n N_VGND_c_183_n 0.0355424f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_102 N_Y_M1000_s N_VGND_c_186_n 0.00224864f $X=0.91 $Y=0.235 $X2=0 $Y2=0
cc_103 N_Y_c_158_n N_VGND_c_186_n 0.0227618f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_104 Y A_110_47# 2.78895e-19 $X=0.605 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_105 N_Y_c_158_n A_110_47# 0.0011988f $X=1.05 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_106 N_VGND_c_186_n A_110_47# 0.00324061f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_107 N_VGND_c_186_n A_268_47# 0.00897657f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

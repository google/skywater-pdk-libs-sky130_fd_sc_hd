* File: sky130_fd_sc_hd__einvp_2.pex.spice
* Created: Thu Aug 27 14:20:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__EINVP_2%TE 3 7 9 10 11 13 14 16 18 19 20 21
c47 14 0 6.76181e-20 $X=1.29 $Y=1.035
r48 25 27 31.7105 $w=3.42e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.142
+ $X2=0.47 $Y2=1.142
r49 20 21 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r50 20 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r51 16 18 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.365 $Y=0.96
+ $X2=1.365 $Y2=0.56
r52 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.035
+ $X2=0.945 $Y2=1.035
r53 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.29 $Y=1.035
+ $X2=1.365 $Y2=0.96
r54 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.035
+ $X2=1.02 $Y2=1.035
r55 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=0.96
+ $X2=0.945 $Y2=1.035
r56 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.945 $Y=0.96
+ $X2=0.945 $Y2=0.56
r57 10 27 26.0143 $w=3.42e-07 $l=1.39549e-07 $layer=POLY_cond $X=0.545 $Y=1.035
+ $X2=0.47 $Y2=1.142
r58 9 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.945 $Y2=1.035
r59 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.545 $Y2=1.035
r60 5 27 22.0749 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.142
r61 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.165
r62 1 27 22.0749 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.47 $Y2=1.142
r63 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%A_27_47# 1 2 7 9 10 11 12 14 16 19 23 26 27
+ 29 30
c67 27 0 1.1096e-19 $X=0.875 $Y=1.16
r68 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r69 27 33 6.10785 $w=4.07e-07 $l=2.26548e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=0.687 $Y2=1.075
r70 27 29 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=1.79 $Y2=1.16
r71 25 33 1.22594 $w=3.75e-07 $l=2.5e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.075
r72 25 26 14.1366 $w=3.73e-07 $l=4.6e-07 $layer=LI1_cond $X=0.687 $Y=1.325
+ $X2=0.687 $Y2=1.785
r73 21 26 30.7936 $w=1.68e-07 $l=4.72e-07 $layer=LI1_cond $X=0.215 $Y=1.87
+ $X2=0.687 $Y2=1.87
r74 21 23 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=1.955
+ $X2=0.215 $Y2=2.165
r75 17 33 14.1484 $w=4.07e-07 $l=6.48864e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.687 $Y2=1.075
r76 17 19 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r77 15 30 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.79 $Y=1.32
+ $X2=1.79 $Y2=1.16
r78 15 16 15.2969 $w=2.1e-07 $l=1.35e-07 $layer=POLY_cond $X=1.79 $Y=1.32
+ $X2=1.655 $Y2=1.32
r79 12 16 15.2969 $w=2.1e-07 $l=2.38485e-07 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.655 $Y2=1.32
r80 12 14 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.83 $Y=1.47
+ $X2=1.83 $Y2=2.015
r81 10 16 10.1846 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=1.395
+ $X2=1.655 $Y2=1.32
r82 10 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.655 $Y=1.395
+ $X2=1.485 $Y2=1.395
r83 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.47
+ $X2=1.485 $Y2=1.395
r84 7 9 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.41 $Y=1.47 $X2=1.41
+ $Y2=2.015
r85 2 23 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r86 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%A 1 3 6 8 10 13 15 16 17 25
r39 23 25 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=2.725 $Y=1.16
+ $X2=2.98 $Y2=1.16
r40 21 23 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.305 $Y=1.16
+ $X2=2.725 $Y2=1.16
r41 15 17 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.992 $Y=1.16
+ $X2=2.992 $Y2=1.53
r42 15 16 12.5353 $w=2.83e-07 $l=3.1e-07 $layer=LI1_cond $X=2.992 $Y=1.16
+ $X2=2.992 $Y2=0.85
r43 15 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.16 $X2=2.98 $Y2=1.16
r44 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.325
+ $X2=2.725 $Y2=1.16
r45 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.725 $Y=1.325
+ $X2=2.725 $Y2=1.985
r46 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=0.995
+ $X2=2.725 $Y2=1.16
r47 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.725 $Y=0.995
+ $X2=2.725 $Y2=0.56
r48 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.325
+ $X2=2.305 $Y2=1.16
r49 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.305 $Y=1.325
+ $X2=2.305 $Y2=1.985
r50 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.995
+ $X2=2.305 $Y2=1.16
r51 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.305 $Y=0.995
+ $X2=2.305 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%VPWR 1 2 9 13 15 17 22 32 33 36 39
r45 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r49 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r53 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 23 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.695 $Y2=2.72
r58 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r60 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 17 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.695 $Y2=2.72
r62 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r63 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r66 11 13 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.02
r67 7 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r68 7 9 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.34
r69 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.545 $X2=1.62 $Y2=2.02
r70 1 9 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%A_215_309# 1 2 3 12 14 15 19 20 21 24
c40 14 0 6.76181e-20 $X=1.985 $Y=1.64
r41 22 24 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=2.992 $Y=2.295
+ $X2=2.992 $Y2=1.96
r42 20 22 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.85 $Y=2.38
+ $X2=2.992 $Y2=2.295
r43 20 21 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.85 $Y=2.38
+ $X2=2.155 $Y2=2.38
r44 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=2.295
+ $X2=2.155 $Y2=2.38
r45 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.07 $Y=2.295
+ $X2=2.07 $Y2=1.96
r46 16 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=1.725
+ $X2=2.07 $Y2=1.96
r47 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=1.64
+ $X2=2.07 $Y2=1.725
r48 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.985 $Y=1.64
+ $X2=1.285 $Y2=1.64
r49 10 15 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.165 $Y=1.725
+ $X2=1.285 $Y2=1.64
r50 10 12 11.2843 $w=2.38e-07 $l=2.35e-07 $layer=LI1_cond $X=1.165 $Y=1.725
+ $X2=1.165 $Y2=1.96
r51 3 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.8
+ $Y=1.485 $X2=2.935 $Y2=1.96
r52 2 19 300 $w=1.7e-07 $l=4.90612e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.545 $X2=2.07 $Y2=1.96
r53 1 12 300 $w=1.7e-07 $l=4.73392e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.545 $X2=1.2 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%Z 1 2 7 8 9 10 16
r18 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.515 $Y=1.53
+ $X2=2.515 $Y2=1.87
r19 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.515 $Y=1.19
+ $X2=2.515 $Y2=1.53
r20 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.515 $Y=0.85
+ $X2=2.515 $Y2=1.19
r21 7 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.515 $Y=0.85 $X2=2.515
+ $Y2=0.76
r22 2 9 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=1.485 $X2=2.515 $Y2=1.61
r23 1 16 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.515 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r53 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r54 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r55 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r56 27 39 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.59
+ $Y2=0
r57 27 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.07
+ $Y2=0
r58 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r59 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r60 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r61 23 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.695
+ $Y2=0
r62 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.15
+ $Y2=0
r63 22 39 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.59
+ $Y2=0
r64 22 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r65 17 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.695
+ $Y2=0
r66 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r67 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r68 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 11 39 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r70 11 13 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.38
r71 7 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r72 7 9 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.36
r73 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.38
r74 1 9 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.71 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__EINVP_2%A_204_47# 1 2 3 12 14 15 19 20 21
r34 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.85 $Y=0.34
+ $X2=2.18 $Y2=0.34
r35 17 19 5.76222 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.06 $Y=0.655
+ $X2=2.06 $Y2=0.535
r36 16 21 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.06 $Y=0.425
+ $X2=2.18 $Y2=0.34
r37 16 19 5.28203 $w=2.38e-07 $l=1.1e-07 $layer=LI1_cond $X=2.06 $Y=0.425
+ $X2=2.06 $Y2=0.535
r38 14 17 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.94 $Y=0.74
+ $X2=2.06 $Y2=0.655
r39 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.94 $Y=0.74 $X2=1.24
+ $Y2=0.74
r40 10 15 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=1.142 $Y=0.655
+ $X2=1.24 $Y2=0.74
r41 10 12 6.82517 $w=1.93e-07 $l=1.2e-07 $layer=LI1_cond $X=1.142 $Y=0.655
+ $X2=1.142 $Y2=0.535
r42 3 20 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.42
r43 2 19 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.235 $X2=2.095 $Y2=0.535
r44 1 12 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.535
.ends


* File: sky130_fd_sc_hd__o41ai_1.spice
* Created: Thu Aug 27 14:42:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o41ai_1.spice.pex"
.subckt sky130_fd_sc_hd__o41ai_1  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_A_109_47#_M1008_d N_B1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.203125 AS=0.169 PD=1.275 PS=1.82 NRD=57.228 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A4_M1007_g N_A_109_47#_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.203125 PD=0.92 PS=1.275 NRD=0 NRS=6.456 M=1 R=4.33333 SA=75001
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1001 N_A_109_47#_M1001_d N_A3_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_109_47#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.08775 PD=1 PS=0.92 NRD=13.836 NRS=0 M=1 R=4.33333 SA=75001.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_A_109_47#_M1009_d N_A1_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.11375 PD=1.86 PS=1 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75002.3 A=0.15
+ P=2.3 MULT=1
MM1003 A_193_297# N_A4_M1003_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=1 AD=0.3125
+ AS=0.135 PD=1.625 PS=1.27 NRD=50.7078 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 A_348_297# N_A3_M1005_g A_193_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.3125 PD=1.27 PS=1.625 NRD=15.7403 NRS=50.7078 M=1 R=6.66667 SA=75001.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1002 A_432_297# N_A2_M1002_g A_348_297# VPB PHIGHVT L=0.15 W=1 AD=0.175
+ AS=0.135 PD=1.35 PS=1.27 NRD=23.6203 NRS=15.7403 M=1 R=6.66667 SA=75001.8
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_432_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.175 PD=2.56 PS=1.35 NRD=0 NRS=23.6203 M=1 R=6.66667 SA=75002.3 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_33 VNB 0 2.99524e-19 $X=0.15 $Y=-0.085
c_55 VPB 0 1.10786e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o41ai_1.spice.SKY130_FD_SC_HD__O41AI_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a21o_1.pxi.spice
* Created: Tue Sep  1 18:52:01 2020
* 
x_PM_SKY130_FD_SC_HD__A21O_1%A_81_21# N_A_81_21#_M1005_d N_A_81_21#_M1007_s
+ N_A_81_21#_c_47_n N_A_81_21#_M1000_g N_A_81_21#_M1003_g N_A_81_21#_c_48_n
+ N_A_81_21#_c_49_n N_A_81_21#_c_56_p N_A_81_21#_c_87_p N_A_81_21#_c_53_n
+ N_A_81_21#_c_54_n N_A_81_21#_c_57_p PM_SKY130_FD_SC_HD__A21O_1%A_81_21#
x_PM_SKY130_FD_SC_HD__A21O_1%B1 N_B1_c_102_n N_B1_M1005_g N_B1_M1007_g B1
+ N_B1_c_104_n PM_SKY130_FD_SC_HD__A21O_1%B1
x_PM_SKY130_FD_SC_HD__A21O_1%A1 N_A1_c_134_n N_A1_M1002_g N_A1_M1004_g A1 A1 A1
+ N_A1_c_137_n PM_SKY130_FD_SC_HD__A21O_1%A1
x_PM_SKY130_FD_SC_HD__A21O_1%A2 N_A2_c_172_n N_A2_M1006_g N_A2_M1001_g A2
+ N_A2_c_174_n PM_SKY130_FD_SC_HD__A21O_1%A2
x_PM_SKY130_FD_SC_HD__A21O_1%X N_X_M1000_s N_X_M1003_s X X X X X X
+ PM_SKY130_FD_SC_HD__A21O_1%X
x_PM_SKY130_FD_SC_HD__A21O_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_c_209_n
+ N_VPWR_c_210_n VPWR N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n
+ N_VPWR_c_208_n N_VPWR_c_215_n N_VPWR_c_216_n PM_SKY130_FD_SC_HD__A21O_1%VPWR
x_PM_SKY130_FD_SC_HD__A21O_1%A_299_297# N_A_299_297#_M1007_d
+ N_A_299_297#_M1001_d N_A_299_297#_c_262_n N_A_299_297#_c_248_n
+ N_A_299_297#_c_250_n N_A_299_297#_c_249_n
+ PM_SKY130_FD_SC_HD__A21O_1%A_299_297#
x_PM_SKY130_FD_SC_HD__A21O_1%VGND N_VGND_M1000_d N_VGND_M1006_d N_VGND_c_268_n
+ N_VGND_c_269_n VGND N_VGND_c_270_n N_VGND_c_271_n N_VGND_c_272_n
+ N_VGND_c_273_n PM_SKY130_FD_SC_HD__A21O_1%VGND
cc_1 VNB N_A_81_21#_c_47_n 0.0231009f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_81_21#_c_48_n 0.00358448f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_3 VNB N_A_81_21#_c_49_n 0.0327653f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.16
cc_4 VNB N_B1_c_102_n 0.0202338f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_5 VNB B1 0.00232662f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_6 VNB N_B1_c_104_n 0.0295434f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=0.835
cc_7 VNB N_A1_c_134_n 0.0165967f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_8 VNB A1 0.00286183f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_9 VNB A1 0.00483389f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.325
cc_10 VNB N_A1_c_137_n 0.0195005f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.505
cc_11 VNB N_A2_c_172_n 0.0222808f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.235
cc_12 VNB A2 0.012123f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_13 VNB N_A2_c_174_n 0.0348997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB X 0.0456623f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_15 VNB N_VPWR_c_208_n 0.117919f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.615
cc_16 VNB N_VGND_c_268_n 0.0111284f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_17 VNB N_VGND_c_269_n 0.0277555f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.985
cc_18 VNB N_VGND_c_270_n 0.0289443f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.505
cc_19 VNB N_VGND_c_271_n 0.0190264f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=1.725
cc_20 VNB N_VGND_c_272_n 0.0204472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_273_n 0.16196f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_22 VPB N_A_81_21#_M1003_g 0.0254972f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_23 VPB N_A_81_21#_c_48_n 0.00266318f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_24 VPB N_A_81_21#_c_49_n 0.009457f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_25 VPB N_A_81_21#_c_53_n 0.0125781f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.725
cc_26 VPB N_A_81_21#_c_54_n 0.00788942f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=1.81
cc_27 VPB N_B1_M1007_g 0.0234061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB B1 6.39252e-19 $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_29 VPB N_B1_c_104_n 0.00890558f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=0.835
cc_30 VPB N_A1_M1004_g 0.0190957f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB A1 0.00266083f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.325
cc_32 VPB N_A1_c_137_n 0.00389059f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.505
cc_33 VPB N_A2_M1001_g 0.0261857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB A2 0.0014041f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_35 VPB N_A2_c_174_n 0.00831796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB X 0.0465418f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_37 VPB N_VPWR_c_209_n 0.00875547f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_38 VPB N_VPWR_c_210_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_211_n 0.0154228f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.16
cc_40 VPB N_VPWR_c_212_n 0.0270775f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.81
cc_41 VPB N_VPWR_c_213_n 0.015741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_208_n 0.0524378f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.615
cc_43 VPB N_VPWR_c_215_n 0.00527117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_216_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_299_297#_c_248_n 0.0104962f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_46 VPB N_A_299_297#_c_249_n 0.0269742f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.505
cc_47 N_A_81_21#_c_48_n N_B1_c_102_n 0.00406515f $X=0.695 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_48 N_A_81_21#_c_56_p N_B1_c_102_n 0.0139604f $X=1.465 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_49 N_A_81_21#_c_57_p N_B1_c_102_n 0.0112465f $X=1.62 $Y=0.635 $X2=-0.19
+ $Y2=-0.24
cc_50 N_A_81_21#_c_48_n N_B1_M1007_g 0.00459023f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_81_21#_c_48_n B1 0.0251485f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_81_21#_c_49_n B1 0.00111096f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_81_21#_c_56_p B1 0.0310103f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_54 N_A_81_21#_c_53_n B1 0.0208522f $X=1.18 $Y=1.725 $X2=0 $Y2=0
cc_55 N_A_81_21#_c_48_n N_B1_c_104_n 0.00135661f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_81_21#_c_49_n N_B1_c_104_n 0.0181897f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_81_21#_c_56_p N_B1_c_104_n 0.00615674f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_58 N_A_81_21#_c_53_n N_B1_c_104_n 0.00542681f $X=1.18 $Y=1.725 $X2=0 $Y2=0
cc_59 N_A_81_21#_c_56_p N_A1_c_134_n 0.00284278f $X=1.465 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_81_21#_c_57_p N_A1_c_134_n 0.00523586f $X=1.62 $Y=0.635 $X2=-0.19
+ $Y2=-0.24
cc_61 N_A_81_21#_c_56_p A1 0.00672348f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_62 N_A_81_21#_c_56_p N_A1_c_137_n 0.00123745f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_63 N_A_81_21#_c_57_p N_A2_c_172_n 3.9243e-19 $X=1.62 $Y=0.635 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_81_21#_c_47_n X 0.0233615f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A_81_21#_c_48_n X 0.0446331f $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_81_21#_c_48_n N_VPWR_M1003_d 6.00252e-19 $X=0.695 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_81_21#_c_53_n N_VPWR_M1003_d 0.00368555f $X=1.18 $Y=1.725 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_81_21#_M1003_g N_VPWR_c_209_n 0.0143519f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_69 N_A_81_21#_c_53_n N_VPWR_c_209_n 0.0208158f $X=1.18 $Y=1.725 $X2=0 $Y2=0
cc_70 N_A_81_21#_c_54_n N_VPWR_c_209_n 0.0434306f $X=1.21 $Y=1.81 $X2=0 $Y2=0
cc_71 N_A_81_21#_M1003_g N_VPWR_c_211_n 0.0046653f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_81_21#_c_54_n N_VPWR_c_212_n 0.0169152f $X=1.21 $Y=1.81 $X2=0 $Y2=0
cc_73 N_A_81_21#_M1007_s N_VPWR_c_208_n 0.00318026f $X=1.085 $Y=1.485 $X2=0
+ $Y2=0
cc_74 N_A_81_21#_M1003_g N_VPWR_c_208_n 0.00896841f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_75 N_A_81_21#_c_54_n N_VPWR_c_208_n 0.0102724f $X=1.21 $Y=1.81 $X2=0 $Y2=0
cc_76 N_A_81_21#_c_56_p N_A_299_297#_c_250_n 0.00339943f $X=1.465 $Y=0.735 $X2=0
+ $Y2=0
cc_77 N_A_81_21#_c_48_n N_VGND_M1000_d 8.12229e-19 $X=0.695 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_81_21#_c_56_p N_VGND_M1000_d 0.0141872f $X=1.465 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_81_21#_c_87_p N_VGND_M1000_d 0.00339863f $X=0.835 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_81_21#_c_56_p N_VGND_c_270_n 0.00257791f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_81 N_A_81_21#_c_57_p N_VGND_c_270_n 0.016407f $X=1.62 $Y=0.635 $X2=0 $Y2=0
cc_82 N_A_81_21#_c_47_n N_VGND_c_271_n 0.00574689f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_81_21#_c_87_p N_VGND_c_271_n 7.8701e-19 $X=0.835 $Y=0.735 $X2=0 $Y2=0
cc_84 N_A_81_21#_c_47_n N_VGND_c_272_n 0.0106589f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_81_21#_c_49_n N_VGND_c_272_n 7.85384e-19 $X=0.695 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_81_21#_c_56_p N_VGND_c_272_n 0.0327754f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_87 N_A_81_21#_c_87_p N_VGND_c_272_n 0.0175141f $X=0.835 $Y=0.735 $X2=0 $Y2=0
cc_88 N_A_81_21#_c_57_p N_VGND_c_272_n 0.0148485f $X=1.62 $Y=0.635 $X2=0 $Y2=0
cc_89 N_A_81_21#_M1005_d N_VGND_c_273_n 0.00221165f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_90 N_A_81_21#_c_47_n N_VGND_c_273_n 0.0127599f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_81_21#_c_56_p N_VGND_c_273_n 0.00660531f $X=1.465 $Y=0.735 $X2=0 $Y2=0
cc_92 N_A_81_21#_c_87_p N_VGND_c_273_n 0.00319797f $X=0.835 $Y=0.735 $X2=0 $Y2=0
cc_93 N_A_81_21#_c_57_p N_VGND_c_273_n 0.0115977f $X=1.62 $Y=0.635 $X2=0 $Y2=0
cc_94 N_B1_c_102_n N_A1_c_134_n 0.0238787f $X=1.42 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_95 N_B1_M1007_g N_A1_M1004_g 0.0254694f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_96 B1 A1 0.0250635f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B1_c_104_n A1 0.00196425f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_98 B1 N_A1_c_137_n 3.41095e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B1_c_104_n N_A1_c_137_n 0.0205223f $X=1.42 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_M1007_g N_VPWR_c_209_n 0.00372692f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1007_g N_VPWR_c_210_n 0.00132212f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1007_g N_VPWR_c_212_n 0.00585385f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1007_g N_VPWR_c_208_n 0.0122297f $X=1.42 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B1_M1007_g N_A_299_297#_c_250_n 0.00122267f $X=1.42 $Y=1.985 $X2=0
+ $Y2=0
cc_105 N_B1_c_102_n N_VGND_c_270_n 0.00413531f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B1_c_102_n N_VGND_c_272_n 0.0103644f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B1_c_102_n N_VGND_c_273_n 0.00706342f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A1_c_134_n N_A2_c_172_n 0.0340161f $X=1.845 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_109 A1 N_A2_c_172_n 0.00541358f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_110 N_A1_M1004_g N_A2_M1001_g 0.0291006f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_111 A1 A2 0.00139643f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_112 A1 A2 0.0243015f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_113 N_A1_c_137_n A2 2.26583e-19 $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_114 A1 N_A2_c_174_n 0.00270532f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A1_c_137_n N_A2_c_174_n 0.019498f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_M1004_g N_VPWR_c_210_n 0.010999f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A1_M1004_g N_VPWR_c_212_n 0.00486043f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A1_M1004_g N_VPWR_c_208_n 0.00831583f $X=1.845 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A1_M1004_g N_A_299_297#_c_248_n 0.0158532f $X=1.845 $Y=1.985 $X2=0
+ $Y2=0
cc_120 A1 N_A_299_297#_c_248_n 0.0283776f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_121 N_A1_c_137_n N_A_299_297#_c_248_n 0.00120793f $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_122 A1 N_A_299_297#_c_250_n 0.00480256f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_123 N_A1_c_137_n N_A_299_297#_c_250_n 3.09916e-19 $X=1.845 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A1_c_134_n N_VGND_c_270_n 0.00579368f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_125 A1 N_VGND_c_270_n 0.00781813f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_126 N_A1_c_134_n N_VGND_c_273_n 0.0107221f $X=1.845 $Y=0.995 $X2=0 $Y2=0
cc_127 A1 N_VGND_c_273_n 0.00819911f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_128 A1 A_384_47# 0.00610384f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_129 N_A2_M1001_g N_VPWR_c_210_n 0.0119226f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A2_M1001_g N_VPWR_c_213_n 0.00486043f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A2_M1001_g N_VPWR_c_208_n 0.00928036f $X=2.275 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_M1001_g N_A_299_297#_c_248_n 0.0217352f $X=2.275 $Y=1.985 $X2=0
+ $Y2=0
cc_133 A2 N_A_299_297#_c_248_n 0.0202417f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A2_c_174_n N_A_299_297#_c_248_n 0.00517789f $X=2.485 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A2_c_172_n N_VGND_c_269_n 0.00861947f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_136 A2 N_VGND_c_269_n 0.0212008f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A2_c_174_n N_VGND_c_269_n 0.00575879f $X=2.485 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A2_c_172_n N_VGND_c_270_n 0.00585385f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_172_n N_VGND_c_273_n 0.0116601f $X=2.275 $Y=0.995 $X2=0 $Y2=0
cc_140 X N_VPWR_c_211_n 0.0169196f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_141 N_X_M1003_s N_VPWR_c_208_n 0.00387432f $X=0.145 $Y=1.485 $X2=0 $Y2=0
cc_142 X N_VPWR_c_208_n 0.00988906f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_143 X N_VGND_c_271_n 0.0169196f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_144 N_X_M1000_s N_VGND_c_273_n 0.00387432f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_145 X N_VGND_c_273_n 0.00988906f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_146 N_VPWR_c_208_n N_A_299_297#_M1007_d 0.00379995f $X=2.53 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_147 N_VPWR_c_208_n N_A_299_297#_M1001_d 0.00374186f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_148 N_VPWR_c_212_n N_A_299_297#_c_262_n 0.0128833f $X=1.895 $Y=2.72 $X2=0
+ $Y2=0
cc_149 N_VPWR_c_208_n N_A_299_297#_c_262_n 0.00873917f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_150 N_VPWR_M1004_d N_A_299_297#_c_248_n 0.00362489f $X=1.92 $Y=1.485 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_210_n N_A_299_297#_c_248_n 0.016744f $X=2.06 $Y=2.02 $X2=0 $Y2=0
cc_152 N_VPWR_c_213_n N_A_299_297#_c_249_n 0.0167431f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_153 N_VPWR_c_208_n N_A_299_297#_c_249_n 0.00988906f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_154 N_VGND_c_273_n A_384_47# 0.00417598f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

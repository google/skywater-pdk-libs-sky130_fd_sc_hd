* File: sky130_fd_sc_hd__ebufn_2.spice
* Created: Tue Sep  1 19:07:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ebufn_2.pex.spice"
.subckt sky130_fd_sc_hd__ebufn_2  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.1092 PD=0.795 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_214_47#_M1008_d N_TE_B_M1008_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.07875 PD=1.36 PS=0.795 NRD=0 NRS=28.56 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_214_47#_M1005_g N_A_392_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1005_d N_A_214_47#_M1007_g N_A_392_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.125125 PD=0.92 PS=1.035 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1003 N_Z_M1003_d N_A_27_47#_M1003_g N_A_392_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.125125 PD=0.92 PS=1.035 NRD=0 NRS=10.152 M=1 R=4.33333
+ SA=75001.1 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_Z_M1003_d N_A_27_47#_M1004_g N_A_392_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.12 AS=0.1664 PD=1.015 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1010 N_A_214_47#_M1010_d N_TE_B_M1010_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.12 PD=1.8 PS=1.015 NRD=0 NRS=13.8491 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_320_309#_M1001_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.2444 PD=1.21 PS=2.4 NRD=0 NRS=0 M=1 R=6.26667 SA=75000.2
+ SB=75001.9 A=0.141 P=2.18 MULT=1
MM1011 N_VPWR_M1001_d N_TE_B_M1011_g N_A_320_309#_M1011_s VPB PHIGHVT L=0.15
+ W=0.94 AD=0.1269 AS=0.358799 PD=1.21 PS=1.69103 NRD=0 NRS=11.5245 M=1
+ R=6.26667 SA=75000.6 SB=75001.5 A=0.141 P=2.18 MULT=1
MM1000 N_A_320_309#_M1011_s N_A_27_47#_M1000_g N_Z_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.381701 AS=0.135 PD=1.79897 PS=1.27 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75001.4 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1002 N_A_320_309#_M1002_d N_A_27_47#_M1002_g N_Z_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__ebufn_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__dfrtp_4.pex.spice
* Created: Tue Sep  1 19:03:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFRTP_4%CLK 1 2 3 5 6 8 11 13 14
c40 6 0 9.23148e-20 $X=0.47 $Y=1.74
c41 1 0 2.71124e-20 $X=0.305 $Y=1.325
r42 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=1.16
+ $X2=0.265 $Y2=1.53
r43 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r44 9 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r45 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r46 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=2.135
r47 3 18 88.7086 $w=2.58e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r49 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r50 1 18 39.2009 $w=2.58e-07 $l=1.75656e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.327 $Y2=1.16
r51 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.305 $Y=1.325
+ $X2=0.305 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_27_47# 1 2 9 13 17 20 21 22 25 27 29 33 37
+ 41 42 43 46 49 50 51 52 55 61 68 71 72 77
c236 77 0 4.56546e-20 $X=6.07 $Y=1.11
c237 61 0 1.76704e-20 $X=6.11 $Y=1.19
c238 51 0 1.58851e-19 $X=5.965 $Y=1.19
c239 29 0 4.11863e-20 $X=5.845 $Y=2.275
c240 22 0 1.90473e-19 $X=2.72 $Y=1.32
r241 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.11 $X2=6.07 $Y2=1.11
r242 71 74 47.4498 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=1.095
r243 71 73 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=0.93
+ $X2=2.585 $Y2=0.765
r244 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.93 $X2=2.585 $Y2=0.93
r245 65 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r246 61 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.19
+ $X2=6.11 $Y2=1.19
r247 59 72 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.56 $Y=1.19
+ $X2=2.56 $Y2=0.93
r248 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.19
r249 55 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r250 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.19
+ $X2=0.695 $Y2=1.19
r251 52 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.19
+ $X2=2.53 $Y2=1.19
r252 51 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=6.11 $Y2=1.19
r253 51 52 4.07177 $w=1.4e-07 $l=3.29e-06 $layer=MET1_cond $X=5.965 $Y=1.19
+ $X2=2.675 $Y2=1.19
r254 50 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.19
+ $X2=0.695 $Y2=1.19
r255 49 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=2.53 $Y2=1.19
r256 49 50 1.91213 $w=1.4e-07 $l=1.545e-06 $layer=MET1_cond $X=2.385 $Y=1.19
+ $X2=0.84 $Y2=1.19
r257 48 55 30.3143 $w=2.28e-07 $l=6.05e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.19
r258 47 55 19.2909 $w=2.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.19
r259 44 46 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r260 43 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.795
r261 43 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r262 41 47 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r263 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r264 35 42 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.345 $Y2=0.72
r265 35 37 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.635
+ $X2=0.217 $Y2=0.51
r266 31 76 38.5991 $w=2.92e-07 $l=1.76125e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=5.987 $Y2=1.11
r267 31 33 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.01 $Y=0.945
+ $X2=6.01 $Y2=0.415
r268 27 76 58.4073 $w=2.92e-07 $l=3.48848e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.987 $Y2=1.11
r269 27 29 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.845 $Y=1.395
+ $X2=5.845 $Y2=2.275
r270 23 25 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.18 $Y=1.395
+ $X2=3.18 $Y2=2.275
r271 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=3.18 $Y2=1.395
r272 21 22 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.105 $Y=1.32
+ $X2=2.72 $Y2=1.32
r273 20 22 26.9401 $w=1.5e-07 $l=1.09243e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.72 $Y2=1.32
r274 20 74 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.642 $Y=1.245
+ $X2=2.642 $Y2=1.095
r275 17 73 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.64 $Y=0.415
+ $X2=2.64 $Y2=0.765
r276 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r277 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r278 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r279 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r280 2 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r281 1 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%D 3 7 9 10 15 19
c53 10 0 1.85993e-19 $X=2.09 $Y=1.3
c54 7 0 1.77283e-19 $X=2.225 $Y=2.275
r55 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.465 $X2=1.79 $Y2=1.465
r56 15 19 1.96287 $w=4.04e-07 $l=6.5e-08 $layer=LI1_cond $X=1.615 $Y=1.53
+ $X2=1.615 $Y2=1.465
r57 9 18 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.09 $Y=1.465 $X2=1.79
+ $Y2=1.465
r58 9 10 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.465
+ $X2=2.09 $Y2=1.3
r59 5 10 37.0704 $w=1.5e-07 $l=3.91727e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.09 $Y2=1.3
r60 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.225 $Y=1.63
+ $X2=2.225 $Y2=2.275
r61 1 10 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.3 $X2=2.09
+ $Y2=1.3
r62 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.165 $Y=1.3
+ $X2=2.165 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_193_47# 1 2 9 13 15 17 20 23 26 27 29 30
+ 34 35 37 38 39 40 47 49 53 65 66 70
c212 66 0 3.94709e-20 $X=6.265 $Y=1.74
c213 47 0 1.77283e-19 $X=2.99 $Y=1.87
c214 39 0 1.36782e-20 $X=5.965 $Y=1.87
c215 38 0 9.23148e-20 $X=1.245 $Y=1.87
c216 37 0 1.20979e-19 $X=2.845 $Y=1.87
c217 35 0 1.61046e-19 $X=3.095 $Y=0.9
c218 29 0 1.76704e-20 $X=5.97 $Y=1.58
c219 26 0 1.28114e-19 $X=5.59 $Y=0.87
r220 65 68 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.74
+ $X2=6.265 $Y2=1.905
r221 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.265
+ $Y=1.74 $X2=6.265 $Y2=1.74
r222 53 56 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.695 $Y=1.74
+ $X2=2.695 $Y2=1.875
r223 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.695
+ $Y=1.74 $X2=2.695 $Y2=1.74
r224 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.11 $Y=1.87
+ $X2=6.11 $Y2=1.87
r225 47 54 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=1.77
+ $X2=2.695 $Y2=1.77
r226 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=1.87
r227 43 70 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.1 $Y=1.87
+ $X2=1.1 $Y2=0.51
r228 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.1 $Y=1.87 $X2=1.1
+ $Y2=1.87
r229 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.135 $Y=1.87
+ $X2=2.99 $Y2=1.87
r230 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=6.11 $Y2=1.87
r231 39 40 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=5.965 $Y=1.87
+ $X2=3.135 $Y2=1.87
r232 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.245 $Y=1.87
+ $X2=1.1 $Y2=1.87
r233 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=2.99 $Y2=1.87
r234 37 38 1.98019 $w=1.4e-07 $l=1.6e-06 $layer=MET1_cond $X=2.845 $Y=1.87
+ $X2=1.245 $Y2=1.87
r235 35 58 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.095 $Y=0.9
+ $X2=3.095 $Y2=0.765
r236 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=0.9 $X2=3.095 $Y2=0.9
r237 31 34 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=0.875
+ $X2=3.095 $Y2=0.875
r238 29 66 5.43733 $w=3.59e-07 $l=2.995e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=6.2 $Y2=1.74
r239 29 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.675 $Y2=1.58
r240 27 60 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.59 $Y=0.87
+ $X2=5.465 $Y2=0.87
r241 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=0.87 $X2=5.59 $Y2=0.87
r242 24 30 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.675 $Y2=1.58
r243 24 26 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=5.57 $Y=1.495
+ $X2=5.57 $Y2=0.87
r244 23 47 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.99 $Y=1.575
+ $X2=2.99 $Y2=1.77
r245 22 31 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=0.875
r246 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.99 $Y=0.985
+ $X2=2.99 $Y2=1.575
r247 20 68 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.275 $Y=2.275
+ $X2=6.275 $Y2=1.905
r248 15 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.87
r249 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.465 $Y=0.705
+ $X2=5.465 $Y2=0.415
r250 13 58 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.12 $Y=0.415
+ $X2=3.12 $Y2=0.765
r251 9 56 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.685 $Y=2.275
+ $X2=2.685 $Y2=1.875
r252 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r253 1 70 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_761_289# 1 2 9 13 15 18 21 23 25 26 27 30
+ 33 36 37
c109 36 0 1.00332e-19 $X=5.145 $Y=0.835
c110 23 0 4.11863e-20 $X=5.19 $Y=1.525
r111 33 35 3.58511 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.36
+ $X2=5.19 $Y2=0.445
r112 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.58 $Y=2.005
+ $X2=5.58 $Y2=2.3
r113 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.58 $Y2=2.005
r114 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.495 $Y=1.92
+ $X2=5.275 $Y2=1.92
r115 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.19 $Y=1.835
+ $X2=5.275 $Y2=1.92
r116 24 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.61
r117 24 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.19 $Y=1.695
+ $X2=5.19 $Y2=1.835
r118 23 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=1.61
r119 23 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.19 $Y=1.525
+ $X2=5.19 $Y2=0.835
r120 21 36 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.835
r121 21 35 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=5.145 $Y=0.705
+ $X2=5.145 $Y2=0.445
r122 18 40 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.775
r123 18 39 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.942 $Y=1.61
+ $X2=3.942 $Y2=1.445
r124 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.61 $X2=3.94 $Y2=1.61
r125 15 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=5.19 $Y2=1.61
r126 15 17 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=5.105 $Y=1.61
+ $X2=3.94 $Y2=1.61
r127 13 39 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=3.95 $Y=0.445
+ $X2=3.95 $Y2=1.445
r128 9 40 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.88 $Y=2.275 $X2=3.88
+ $Y2=1.775
r129 2 30 600 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_PDIFF $count=1 $X=5.425
+ $Y=1.645 $X2=5.58 $Y2=2.3
r130 1 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.235 $X2=5.2 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%RESET_B 3 6 10 14 16 17 20 23 25 26 27 29 37
+ 39 42 57
c154 37 0 1.00332e-19 $X=4.37 $Y=0.93
c155 29 0 4.83118e-21 $X=7.19 $Y=1.165
c156 23 0 6.10372e-20 $X=4.25 $Y=0.85
c157 14 0 1.03533e-19 $X=7.235 $Y=2.275
c158 10 0 4.70414e-20 $X=7.235 $Y=0.445
r159 49 57 3.2703 $w=2.4e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=1.035
+ $X2=7.525 $Y2=1.22
r160 42 45 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=1.285
r161 42 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.12
+ $X2=7.27 $Y2=0.955
r162 37 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=1.095
r163 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.93
+ $X2=4.37 $Y2=0.765
r164 30 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.12 $X2=7.27 $Y2=1.12
r165 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.19 $Y=1.165
+ $X2=7.19 $Y2=1.165
r166 27 34 0.181159 $w=2.07e-07 $l=3e-07 $layer=MET1_cond $X=7.19 $Y=0.85
+ $X2=7.49 $Y2=0.85
r167 27 29 0.0979621 $w=2.9e-07 $l=2e-07 $layer=MET1_cond $X=7.19 $Y=0.965
+ $X2=7.19 $Y2=1.165
r168 25 27 0.10072 $w=2.07e-07 $l=1.45e-07 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=7.19 $Y2=0.85
r169 25 26 3.2797 $w=1.4e-07 $l=2.65e-06 $layer=MET1_cond $X=7.045 $Y=0.85
+ $X2=4.395 $Y2=0.85
r170 23 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=0.93 $X2=4.37 $Y2=0.93
r171 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.25 $Y=0.85
+ $X2=4.25 $Y2=0.85
r172 20 26 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.395 $Y2=0.85
r173 20 22 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=4.28 $Y=0.85
+ $X2=4.25 $Y2=0.85
r174 17 57 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.49 $Y=1.22
+ $X2=7.525 $Y2=1.22
r175 17 30 9.34413 $w=3.68e-07 $l=3e-07 $layer=LI1_cond $X=7.49 $Y=1.22 $X2=7.19
+ $Y2=1.22
r176 16 49 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=7.525 $Y=0.85
+ $X2=7.525 $Y2=1.035
r177 16 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.49 $Y=0.85
+ $X2=7.49 $Y2=0.85
r178 14 45 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=7.235 $Y=2.275
+ $X2=7.235 $Y2=1.285
r179 10 44 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.235 $Y=0.445
+ $X2=7.235 $Y2=0.955
r180 6 40 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=4.365 $Y=2.275
+ $X2=4.365 $Y2=1.095
r181 3 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_543_47# 1 2 9 11 13 15 16 20 25 27 28 29
+ 34 35
c126 35 0 6.10372e-20 $X=4.85 $Y=1.17
c127 29 0 1.61046e-19 $X=3.6 $Y=1.27
c128 11 0 1.36782e-20 $X=5.275 $Y=1.495
c129 9 0 1.28114e-19 $X=4.97 $Y=0.555
r130 34 37 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.85 $Y=1.17 $X2=4.85
+ $Y2=1.27
r131 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.17 $X2=4.85 $Y2=1.17
r132 30 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.33 $Y=1.27
+ $X2=3.515 $Y2=1.27
r133 29 32 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.27
+ $X2=3.515 $Y2=1.27
r134 28 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=4.85 $Y2=1.27
r135 28 29 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.765 $Y=1.27
+ $X2=3.6 $Y2=1.27
r136 27 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=1.185
+ $X2=3.515 $Y2=1.27
r137 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.515 $Y=0.475
+ $X2=3.515 $Y2=1.185
r138 24 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=1.27
r139 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.33 $Y=1.355
+ $X2=3.33 $Y2=2.135
r140 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=3.515 $Y2=0.475
r141 20 22 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.43 $Y=0.39
+ $X2=2.91 $Y2=0.39
r142 16 25 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=3.33 $Y2=2.135
r143 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.245 $Y=2.3
+ $X2=2.9 $Y2=2.3
r144 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=5.35 $Y=1.57
+ $X2=5.35 $Y2=2.065
r145 12 35 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=5.045 $Y=1.495
+ $X2=4.88 $Y2=1.17
r146 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.35 $Y2=1.57
r147 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.275 $Y=1.495
+ $X2=5.045 $Y2=1.495
r148 7 35 39.2931 $w=2.55e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.88 $Y2=1.17
r149 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.97 $Y=1.005
+ $X2=4.97 $Y2=0.555
r150 2 18 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.065 $X2=2.9 $Y2=2.33
r151 1 22 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.91 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_1283_21# 1 2 9 13 15 17 20 22 24 27 29 31
+ 34 36 38 41 45 49 50 51 54 56 57 58 59 60 61 67 72 78 86
c202 86 0 1.79991e-19 $X=9.89 $Y=1.16
c203 78 0 6.15427e-20 $X=6.695 $Y=0.98
c204 72 0 1.94811e-19 $X=7.15 $Y=0.78
c205 60 0 1.99375e-19 $X=8.075 $Y=1.295
c206 13 0 2.35828e-20 $X=6.695 $Y=2.275
r207 83 84 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=9.05 $Y=1.16
+ $X2=9.47 $Y2=1.16
r208 68 86 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=9.68 $Y=1.16
+ $X2=9.89 $Y2=1.16
r209 68 84 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=9.68 $Y=1.16
+ $X2=9.47 $Y2=1.16
r210 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.68
+ $Y=1.16 $X2=9.68 $Y2=1.16
r211 65 83 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=8.66 $Y=1.16
+ $X2=9.05 $Y2=1.16
r212 65 80 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.66 $Y=1.16 $X2=8.63
+ $Y2=1.16
r213 64 67 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=8.66 $Y=1.18
+ $X2=9.68 $Y2=1.18
r214 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.66
+ $Y=1.16 $X2=8.66 $Y2=1.16
r215 62 76 3.45218 $w=2.1e-07 $l=1.73e-07 $layer=LI1_cond $X=8.16 $Y=1.18
+ $X2=7.987 $Y2=1.18
r216 62 64 26.4069 $w=2.08e-07 $l=5e-07 $layer=LI1_cond $X=8.16 $Y=1.18 $X2=8.66
+ $Y2=1.18
r217 60 76 7.13508 $w=3.34e-07 $l=1.52791e-07 $layer=LI1_cond $X=8.075 $Y=1.295
+ $X2=7.987 $Y2=1.18
r218 60 61 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.075 $Y=1.295
+ $X2=8.075 $Y2=1.915
r219 59 76 13.1497 $w=3.34e-07 $l=3.65951e-07 $layer=LI1_cond $X=7.975 $Y=0.82
+ $X2=7.987 $Y2=1.18
r220 58 75 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.38
r221 58 59 12.7849 $w=3.18e-07 $l=3.55e-07 $layer=LI1_cond $X=7.975 $Y=0.465
+ $X2=7.975 $Y2=0.82
r222 56 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=2
+ $X2=8.075 $Y2=1.915
r223 56 57 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.99 $Y=2 $X2=7.53
+ $Y2=2
r224 52 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.53 $Y2=2
r225 52 54 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=2.085
+ $X2=7.445 $Y2=2.21
r226 50 75 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.975 $Y2=0.38
r227 50 51 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.815 $Y=0.38
+ $X2=7.235 $Y2=0.38
r228 49 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.695
+ $X2=7.15 $Y2=0.78
r229 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.235 $Y2=0.38
r230 48 49 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=7.15 $Y=0.465
+ $X2=7.15 $Y2=0.695
r231 46 78 17.8171 $w=2.57e-07 $l=9.5e-08 $layer=POLY_cond $X=6.79 $Y=0.98
+ $X2=6.695 $Y2=0.98
r232 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=0.98 $X2=6.79 $Y2=0.98
r233 43 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.815 $Y=0.78
+ $X2=7.15 $Y2=0.78
r234 43 45 6.02413 $w=2.18e-07 $l=1.15e-07 $layer=LI1_cond $X=6.815 $Y=0.865
+ $X2=6.815 $Y2=0.98
r235 39 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.89 $Y=1.325
+ $X2=9.89 $Y2=1.16
r236 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.89 $Y=1.325
+ $X2=9.89 $Y2=1.985
r237 36 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.89 $Y=0.995
+ $X2=9.89 $Y2=1.16
r238 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.89 $Y=0.995
+ $X2=9.89 $Y2=0.56
r239 32 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.47 $Y=1.325
+ $X2=9.47 $Y2=1.16
r240 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.47 $Y=1.325
+ $X2=9.47 $Y2=1.985
r241 29 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.47 $Y=0.995
+ $X2=9.47 $Y2=1.16
r242 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.47 $Y=0.995
+ $X2=9.47 $Y2=0.56
r243 25 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.325
+ $X2=9.05 $Y2=1.16
r244 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.05 $Y=1.325
+ $X2=9.05 $Y2=1.985
r245 22 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=0.995
+ $X2=9.05 $Y2=1.16
r246 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.05 $Y=0.995
+ $X2=9.05 $Y2=0.56
r247 18 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.325
+ $X2=8.63 $Y2=1.16
r248 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.63 $Y=1.325
+ $X2=8.63 $Y2=1.985
r249 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=1.16
r250 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.63 $Y=0.995
+ $X2=8.63 $Y2=0.56
r251 11 78 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=0.98
r252 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=6.695 $Y=1.145
+ $X2=6.695 $Y2=2.275
r253 7 78 38.4475 $w=2.57e-07 $l=2.75409e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.695 $Y2=0.98
r254 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.49 $Y=0.815
+ $X2=6.49 $Y2=0.445
r255 2 54 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=2.065 $X2=7.445 $Y2=2.21
r256 1 75 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=7.765
+ $Y=0.235 $X2=7.9 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_1108_47# 1 2 9 13 15 19 24 25 26 29 30
c103 25 0 2.04429e-20 $X=6.685 $Y=1.745
c104 24 0 1.60161e-19 $X=6.45 $Y=1.315
c105 19 0 1.03533e-19 $X=6.6 $Y=2.295
c106 15 0 4.70414e-20 $X=6.365 $Y=0.395
c107 13 0 1.79199e-19 $X=7.69 $Y=0.445
r108 30 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.66
+ $X2=7.655 $Y2=1.495
r109 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.655
+ $Y=1.66 $X2=7.655 $Y2=1.66
r110 27 32 3.26844 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.77 $Y=1.66 $X2=6.6
+ $Y2=1.66
r111 27 29 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=6.77 $Y=1.66
+ $X2=7.655 $Y2=1.66
r112 25 32 5.45986 $w=2.62e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.6 $Y2=1.66
r113 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.685 $Y=1.745
+ $X2=6.685 $Y2=2.125
r114 24 32 17.5667 $w=2.62e-07 $l=4.13249e-07 $layer=LI1_cond $X=6.45 $Y=1.315
+ $X2=6.6 $Y2=1.66
r115 23 24 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.45 $Y=0.535
+ $X2=6.45 $Y2=1.315
r116 19 26 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.685 $Y2=2.125
r117 19 21 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=6.6 $Y=2.295
+ $X2=6.065 $Y2=2.295
r118 15 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=6.45 $Y2=0.535
r119 15 17 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.365 $Y=0.395
+ $X2=5.75 $Y2=0.395
r120 13 34 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=7.69 $Y=0.445
+ $X2=7.69 $Y2=1.495
r121 7 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=1.66
r122 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.655 $Y=1.825
+ $X2=7.655 $Y2=2.275
r123 2 21 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=2.065 $X2=6.065 $Y2=2.335
r124 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.235 $X2=5.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 62 65 66 68 69 71 72 74 75 77 78 80 81 82 84 89 98 119 120 123 126 129
c169 54 0 1.79991e-19 $X=8.42 $Y=2
c170 9 0 7.44113e-20 $X=9.965 $Y=1.485
r171 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r172 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r173 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r174 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r175 117 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r176 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r177 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r178 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r179 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r180 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r181 108 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r182 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r183 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r184 105 130 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.29 $Y2=2.72
r185 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r186 102 129 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=5.14 $Y2=2.72
r187 102 104 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.325 $Y=2.72
+ $X2=6.67 $Y2=2.72
r188 101 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r189 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r190 98 129 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.14 $Y2=2.72
r191 98 100 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r192 97 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r193 97 127 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.07 $Y2=2.72
r194 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r195 94 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=1.975 $Y2=2.72
r196 94 96 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=2.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r197 93 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r198 93 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r199 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r200 90 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r201 90 92 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r202 89 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.975 $Y2=2.72
r203 89 92 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r204 84 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r205 84 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r206 82 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r207 82 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r208 80 116 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.015 $Y=2.72
+ $X2=9.89 $Y2=2.72
r209 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.015 $Y=2.72
+ $X2=10.1 $Y2=2.72
r210 79 119 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.185 $Y=2.72
+ $X2=10.35 $Y2=2.72
r211 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.185 $Y=2.72
+ $X2=10.1 $Y2=2.72
r212 77 113 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=9.175 $Y=2.72
+ $X2=8.97 $Y2=2.72
r213 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.175 $Y=2.72
+ $X2=9.26 $Y2=2.72
r214 76 116 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=9.345 $Y=2.72
+ $X2=9.89 $Y2=2.72
r215 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=2.72
+ $X2=9.26 $Y2=2.72
r216 74 110 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.335 $Y=2.72
+ $X2=8.05 $Y2=2.72
r217 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=2.72
+ $X2=8.42 $Y2=2.72
r218 73 113 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.505 $Y=2.72
+ $X2=8.97 $Y2=2.72
r219 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=2.72
+ $X2=8.42 $Y2=2.72
r220 71 107 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r221 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.875 $Y2=2.72
r222 70 110 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=8.05 $Y2=2.72
r223 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=7.875 $Y2=2.72
r224 68 104 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.67 $Y2=2.72
r225 68 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.065 $Y2=2.72
r226 67 107 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.59 $Y2=2.72
r227 67 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.19 $Y=2.72
+ $X2=7.065 $Y2=2.72
r228 65 96 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.99 $Y=2.72 $X2=3.91
+ $Y2=2.72
r229 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=2.72
+ $X2=4.155 $Y2=2.72
r230 64 100 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.83 $Y2=2.72
r231 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.72
+ $X2=4.155 $Y2=2.72
r232 60 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.1 $Y=2.635
+ $X2=10.1 $Y2=2.72
r233 60 62 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=10.1 $Y=2.635
+ $X2=10.1 $Y2=1.96
r234 56 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=2.635
+ $X2=9.26 $Y2=2.72
r235 56 58 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=9.26 $Y=2.635
+ $X2=9.26 $Y2=1.96
r236 52 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=2.635
+ $X2=8.42 $Y2=2.72
r237 52 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.42 $Y=2.635
+ $X2=8.42 $Y2=2
r238 48 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.72
r239 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.34
r240 44 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.72
r241 44 46 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2.34
r242 40 129 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.72
r243 40 42 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.14 $Y=2.635
+ $X2=5.14 $Y2=2.34
r244 36 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.72
r245 36 38 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.155 $Y=2.635
+ $X2=4.155 $Y2=2.29
r246 32 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.72
r247 32 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=2.635
+ $X2=1.975 $Y2=2.34
r248 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r249 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r250 9 62 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.965
+ $Y=1.485 $X2=10.1 $Y2=1.96
r251 8 58 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=9.125
+ $Y=1.485 $X2=9.26 $Y2=1.96
r252 7 54 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=1.485 $X2=8.42 $Y2=2
r253 6 50 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=7.73
+ $Y=2.065 $X2=7.875 $Y2=2.34
r254 5 46 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=2.065 $X2=7.025 $Y2=2.34
r255 4 42 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=1.645 $X2=5.14 $Y2=2.34
r256 3 38 600 $w=1.7e-07 $l=3.09233e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=2.065 $X2=4.155 $Y2=2.29
r257 2 34 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.065 $X2=2.015 $Y2=2.34
r258 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_448_47# 1 2 8 9 11
c34 8 0 6.94938e-20 $X=2.13 $Y=1.835
r35 9 11 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.215 $Y=0.39
+ $X2=2.375 $Y2=0.39
r36 8 14 22.5629 $w=2.72e-07 $l=5.35635e-07 $layer=LI1_cond $X=2.13 $Y=1.835
+ $X2=2.282 $Y2=2.3
r37 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.215 $Y2=0.39
r38 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.13 $Y=0.475
+ $X2=2.13 $Y2=1.835
r39 2 14 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.065 $X2=2.435 $Y2=2.3
r40 1 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%A_651_413# 1 2 9 11 12 15
c36 12 0 1.58851e-19 $X=3.755 $Y=1.95
r37 13 15 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.575 $Y=2.035
+ $X2=4.575 $Y2=2.21
r38 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=4.575 $Y2=2.035
r39 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.49 $Y=1.95
+ $X2=3.755 $Y2=1.95
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.755 $Y2=1.95
r41 7 9 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.67 $Y=2.035
+ $X2=3.67 $Y2=2.21
r42 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.065 $X2=4.575 $Y2=2.21
r43 1 9 600 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.065 $X2=3.67 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%Q 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 41 42 43 44 50 51
c79 35 0 7.44058e-20 $X=10.03 $Y=0.82
c80 33 0 7.44113e-20 $X=10.03 $Y=1.54
r81 44 51 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=1.54
+ $X2=10.235 $Y2=1.455
r82 44 51 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=10.235 $Y=1.45
+ $X2=10.235 $Y2=1.455
r83 43 44 7.30818 $w=4.08e-07 $l=2.6e-07 $layer=LI1_cond $X=10.235 $Y=1.19
+ $X2=10.235 $Y2=1.45
r84 42 50 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=0.82
+ $X2=10.235 $Y2=0.905
r85 42 43 7.58926 $w=4.08e-07 $l=2.7e-07 $layer=LI1_cond $X=10.235 $Y=0.92
+ $X2=10.235 $Y2=1.19
r86 42 50 0.421625 $w=4.08e-07 $l=1.5e-08 $layer=LI1_cond $X=10.235 $Y=0.92
+ $X2=10.235 $Y2=0.905
r87 36 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.845 $Y=0.82
+ $X2=9.68 $Y2=0.82
r88 35 42 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=10.03 $Y=0.82
+ $X2=10.235 $Y2=0.82
r89 35 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=10.03 $Y=0.82
+ $X2=9.845 $Y2=0.82
r90 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.805 $Y=1.54
+ $X2=9.68 $Y2=1.54
r91 33 44 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=10.03 $Y=1.54
+ $X2=10.235 $Y2=1.54
r92 33 34 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.03 $Y=1.54
+ $X2=9.805 $Y2=1.54
r93 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.68 $Y=1.625
+ $X2=9.68 $Y2=1.54
r94 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.68 $Y=1.625
+ $X2=9.68 $Y2=2.3
r95 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.68 $Y=0.735
+ $X2=9.68 $Y2=0.82
r96 25 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.68 $Y=0.735
+ $X2=9.68 $Y2=0.39
r97 24 38 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.005 $Y=1.54
+ $X2=8.86 $Y2=1.54
r98 23 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.555 $Y=1.54
+ $X2=9.68 $Y2=1.54
r99 23 24 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=9.555 $Y=1.54
+ $X2=9.005 $Y2=1.54
r100 21 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.515 $Y=0.82
+ $X2=9.68 $Y2=0.82
r101 21 22 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.515 $Y=0.82
+ $X2=9.005 $Y2=0.82
r102 17 38 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=1.625
+ $X2=8.86 $Y2=1.54
r103 17 19 26.8241 $w=2.88e-07 $l=6.75e-07 $layer=LI1_cond $X=8.86 $Y=1.625
+ $X2=8.86 $Y2=2.3
r104 13 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.84 $Y=0.735
+ $X2=9.005 $Y2=0.82
r105 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=8.84 $Y=0.735
+ $X2=8.84 $Y2=0.39
r106 4 41 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=1.485 $X2=9.68 $Y2=1.62
r107 4 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.545
+ $Y=1.485 $X2=9.68 $Y2=2.3
r108 3 38 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.485 $X2=8.84 $Y2=1.62
r109 3 19 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.485 $X2=8.84 $Y2=2.3
r110 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.545
+ $Y=0.235 $X2=9.68 $Y2=0.39
r111 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.705
+ $Y=0.235 $X2=8.84 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFRTP_4%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 50
+ 53 54 56 57 59 60 62 63 65 66 67 69 100 101 104 107
c167 101 0 2.26487e-19 $X=10.35 $Y=0
c168 7 0 7.44058e-20 $X=9.965 $Y=0.235
r169 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r170 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r171 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r172 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r173 98 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r174 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r175 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r176 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r177 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r178 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r179 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r180 88 91 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r181 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r182 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r183 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r184 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r185 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r186 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r187 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r188 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r189 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r190 77 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r191 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=4.37
+ $Y2=0
r192 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r193 74 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.71 $Y2=0
r194 74 76 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.07 $Y2=0
r195 69 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r196 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r197 67 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r198 67 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r199 65 97 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.015 $Y=0
+ $X2=9.89 $Y2=0
r200 65 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.015 $Y=0 $X2=10.1
+ $Y2=0
r201 64 100 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=10.35 $Y2=0
r202 64 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.185 $Y=0 $X2=10.1
+ $Y2=0
r203 62 94 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=9.175 $Y=0
+ $X2=8.97 $Y2=0
r204 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.26
+ $Y2=0
r205 61 97 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=9.345 $Y=0
+ $X2=9.89 $Y2=0
r206 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=0 $X2=9.26
+ $Y2=0
r207 59 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.335 $Y=0
+ $X2=8.05 $Y2=0
r208 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0 $X2=8.42
+ $Y2=0
r209 58 94 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.505 $Y=0
+ $X2=8.97 $Y2=0
r210 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.42
+ $Y2=0
r211 56 85 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.67
+ $Y2=0
r212 56 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.8
+ $Y2=0
r213 55 88 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.895 $Y=0
+ $X2=7.13 $Y2=0
r214 55 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.8
+ $Y2=0
r215 53 79 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r216 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.64
+ $Y2=0
r217 52 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.83
+ $Y2=0
r218 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=0 $X2=4.64
+ $Y2=0
r219 48 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.1 $Y=0.085
+ $X2=10.1 $Y2=0
r220 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.1 $Y=0.085
+ $X2=10.1 $Y2=0.39
r221 44 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0
r222 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0.39
r223 40 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r224 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.39
r225 36 57 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0
r226 36 38 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0.36
r227 32 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0
r228 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.64 $Y=0.085
+ $X2=4.64 $Y2=0.38
r229 28 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r230 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.36
r231 27 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r232 26 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=0
+ $X2=1.71 $Y2=0
r233 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=0.845
+ $Y2=0
r234 22 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r235 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r236 7 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.965
+ $Y=0.235 $X2=10.1 $Y2=0.39
r237 6 46 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.125
+ $Y=0.235 $X2=9.26 $Y2=0.39
r238 5 42 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=8.295
+ $Y=0.235 $X2=8.42 $Y2=0.39
r239 4 38 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.81 $Y2=0.36
r240 3 34 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.64 $Y2=0.38
r241 2 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.71 $Y2=0.36
r242 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o311ai_2.spice.SKY130_FD_SC_HD__O311AI_2.pxi
* Created: Thu Aug 27 14:39:33 2020
* 
x_PM_SKY130_FD_SC_HD__O311AI_2%A1 N_A1_M1002_g N_A1_M1003_g N_A1_M1019_g
+ N_A1_M1016_g A1 A1 N_A1_c_96_n N_A1_c_97_n PM_SKY130_FD_SC_HD__O311AI_2%A1
x_PM_SKY130_FD_SC_HD__O311AI_2%A2 N_A2_M1006_g N_A2_M1009_g N_A2_M1010_g
+ N_A2_M1018_g A2 A2 N_A2_c_137_n PM_SKY130_FD_SC_HD__O311AI_2%A2
x_PM_SKY130_FD_SC_HD__O311AI_2%A3 N_A3_M1013_g N_A3_M1000_g N_A3_M1014_g
+ N_A3_M1001_g N_A3_c_186_n A3 A3 N_A3_c_187_n N_A3_c_188_n
+ PM_SKY130_FD_SC_HD__O311AI_2%A3
x_PM_SKY130_FD_SC_HD__O311AI_2%B1 N_B1_M1005_g N_B1_M1011_g N_B1_M1008_g
+ N_B1_M1015_g B1 B1 N_B1_c_234_n N_B1_c_235_n PM_SKY130_FD_SC_HD__O311AI_2%B1
x_PM_SKY130_FD_SC_HD__O311AI_2%C1 N_C1_M1004_g N_C1_M1007_g N_C1_M1012_g
+ N_C1_M1017_g C1 C1 N_C1_c_279_n N_C1_c_280_n PM_SKY130_FD_SC_HD__O311AI_2%C1
x_PM_SKY130_FD_SC_HD__O311AI_2%A_51_297# N_A_51_297#_M1002_s N_A_51_297#_M1019_s
+ N_A_51_297#_M1010_d N_A_51_297#_c_317_n N_A_51_297#_c_322_n
+ N_A_51_297#_c_318_n N_A_51_297#_c_337_p N_A_51_297#_c_319_n
+ N_A_51_297#_c_320_n N_A_51_297#_c_321_n PM_SKY130_FD_SC_HD__O311AI_2%A_51_297#
x_PM_SKY130_FD_SC_HD__O311AI_2%VPWR N_VPWR_M1002_d N_VPWR_M1011_s N_VPWR_M1004_s
+ N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n
+ VPWR N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_354_n N_VPWR_c_363_n
+ N_VPWR_c_364_n PM_SKY130_FD_SC_HD__O311AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O311AI_2%A_301_297# N_A_301_297#_M1006_s
+ N_A_301_297#_M1000_s N_A_301_297#_c_425_n N_A_301_297#_c_424_n
+ N_A_301_297#_c_428_n N_A_301_297#_c_432_n
+ PM_SKY130_FD_SC_HD__O311AI_2%A_301_297#
x_PM_SKY130_FD_SC_HD__O311AI_2%Y N_Y_M1007_d N_Y_M1017_d N_Y_M1000_d N_Y_M1001_d
+ N_Y_M1015_d N_Y_M1012_d N_Y_c_462_n N_Y_c_454_n N_Y_c_500_n N_Y_c_468_n
+ N_Y_c_504_n N_Y_c_455_n N_Y_c_456_n N_Y_c_450_n Y Y Y Y Y Y Y N_Y_c_453_n
+ N_Y_c_460_n PM_SKY130_FD_SC_HD__O311AI_2%Y
x_PM_SKY130_FD_SC_HD__O311AI_2%A_55_47# N_A_55_47#_M1003_d N_A_55_47#_M1016_d
+ N_A_55_47#_M1018_s N_A_55_47#_M1014_d N_A_55_47#_M1008_d N_A_55_47#_c_534_n
+ N_A_55_47#_c_570_p N_A_55_47#_c_540_n N_A_55_47#_c_583_p N_A_55_47#_c_547_n
+ N_A_55_47#_c_573_p N_A_55_47#_c_529_n N_A_55_47#_c_530_n N_A_55_47#_c_531_n
+ N_A_55_47#_c_532_n N_A_55_47#_c_533_n PM_SKY130_FD_SC_HD__O311AI_2%A_55_47#
x_PM_SKY130_FD_SC_HD__O311AI_2%VGND N_VGND_M1003_s N_VGND_M1009_d N_VGND_M1013_s
+ N_VGND_c_597_n N_VGND_c_598_n VGND N_VGND_c_599_n N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n N_VGND_c_605_n
+ PM_SKY130_FD_SC_HD__O311AI_2%VGND
x_PM_SKY130_FD_SC_HD__O311AI_2%A_729_47# N_A_729_47#_M1005_s N_A_729_47#_M1007_s
+ N_A_729_47#_c_677_n PM_SKY130_FD_SC_HD__O311AI_2%A_729_47#
cc_1 VNB N_A1_M1002_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.985
cc_2 VNB N_A1_M1003_g 0.0240758f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.56
cc_3 VNB N_A1_M1019_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_4 VNB N_A1_M1016_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_5 VNB N_A1_c_96_n 0.016487f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.16
cc_6 VNB N_A1_c_97_n 0.0406106f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.16
cc_7 VNB N_A2_M1006_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.985
cc_8 VNB N_A2_M1009_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.56
cc_9 VNB N_A2_M1010_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_10 VNB N_A2_M1018_g 0.0175231f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_11 VNB A2 0.00495458f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_12 VNB N_A2_c_137_n 0.0353237f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.16
cc_13 VNB N_A3_M1013_g 0.0209052f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.985
cc_14 VNB N_A3_M1000_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.56
cc_15 VNB N_A3_M1014_g 0.0209052f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_16 VNB N_A3_M1001_g 4.60355e-19 $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_17 VNB N_A3_c_186_n 0.0160247f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_A3_c_187_n 0.0259544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A3_c_188_n 0.0318984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B1_M1005_g 0.0177503f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.985
cc_21 VNB N_B1_M1011_g 4.6156e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.56
cc_22 VNB N_B1_M1008_g 0.0216741f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_23 VNB N_B1_M1015_g 5.5242e-19 $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_24 VNB N_B1_c_234_n 0.00297107f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.16
cc_25 VNB N_B1_c_235_n 0.0640843f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.16
cc_26 VNB N_C1_M1004_g 4.55087e-19 $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.985
cc_27 VNB N_C1_M1007_g 0.0217573f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.56
cc_28 VNB N_C1_M1012_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_29 VNB N_C1_M1017_g 0.0242935f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_30 VNB C1 0.0114934f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_31 VNB N_C1_c_279_n 0.0275777f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_32 VNB N_C1_c_280_n 0.0318124f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.16
cc_33 VNB N_VPWR_c_354_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_450_n 0.0134713f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.185
cc_35 VNB Y 0.0057336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB Y 0.0188522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_453_n 0.0026753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_55_47#_c_529_n 0.00257306f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.185
cc_39 VNB N_A_55_47#_c_530_n 0.0333437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_55_47#_c_531_n 0.00222126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_55_47#_c_532_n 0.00143487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_55_47#_c_533_n 0.00199231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_597_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.56
cc_44 VNB N_VGND_c_598_n 3.01556e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_45 VNB N_VGND_c_599_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_600_n 0.0685078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_601_n 0.299434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_602_n 0.021824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_603_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_604_n 0.0110169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_605_n 0.0146419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_729_47#_c_677_n 0.0093693f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.985
cc_53 VPB N_A1_M1002_g 0.0271545f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_54 VPB N_A1_M1019_g 0.0195548f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_55 VPB N_A1_c_96_n 0.00713673f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_56 VPB N_A2_M1006_g 0.019782f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_57 VPB N_A2_M1010_g 0.0273817f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_58 VPB A2 0.005487f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_59 VPB N_A3_M1000_g 0.0273817f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.56
cc_60 VPB N_A3_M1001_g 0.0198668f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.56
cc_61 VPB A3 0.00809882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B1_M1011_g 0.0228236f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.56
cc_63 VPB N_B1_M1015_g 0.0242859f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.56
cc_64 VPB N_B1_c_234_n 0.00746483f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.16
cc_65 VPB N_C1_M1004_g 0.0201298f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.985
cc_66 VPB N_C1_M1012_g 0.0271411f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_67 VPB C1 0.00652041f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_68 VPB N_A_51_297#_c_317_n 0.0338711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_51_297#_c_318_n 0.0147035f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.56
cc_70 VPB N_A_51_297#_c_319_n 0.00481323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_51_297#_c_320_n 0.0038648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_51_297#_c_321_n 0.00239282f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_73 VPB N_VPWR_c_355_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.56
cc_74 VPB N_VPWR_c_356_n 0.00179753f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_75 VPB N_VPWR_c_357_n 4.18394e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_358_n 0.0156295f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_77 VPB N_VPWR_c_359_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.16
cc_78 VPB N_VPWR_c_360_n 0.064509f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_361_n 0.0181828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_354_n 0.0486665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_363_n 0.0221032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_364_n 0.0103759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_301_297#_c_424_n 0.0109117f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=1.985
cc_84 VPB N_Y_c_454_n 0.00364642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_Y_c_455_n 0.00159718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Y_c_456_n 0.0143437f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.185
cc_87 VPB Y 0.0038648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB Y 0.00209956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB Y 0.00134401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_460_n 0.0347398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 N_A1_M1019_g N_A2_M1006_g 0.0282041f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A1_M1016_g N_A2_M1009_g 0.0251782f $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_93 N_A1_c_96_n A2 0.0230876f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_c_97_n A2 8.99031e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A1_c_96_n N_A2_c_137_n 2.70316e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_c_97_n N_A2_c_137_n 0.0181851f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A1_M1002_g N_A_51_297#_c_322_n 0.0170415f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A1_M1019_g N_A_51_297#_c_322_n 0.0156313f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A1_c_96_n N_A_51_297#_c_322_n 0.0411931f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_c_97_n N_A_51_297#_c_322_n 6.15477e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_96_n N_A_51_297#_c_318_n 0.0323661f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_c_97_n N_A_51_297#_c_318_n 2.05204e-19 $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A1_M1002_g N_VPWR_c_355_n 0.0123094f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A1_M1019_g N_VPWR_c_355_n 0.0116083f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A1_M1019_g N_VPWR_c_360_n 0.0046653f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A1_M1002_g N_VPWR_c_354_n 0.00905913f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A1_M1019_g N_VPWR_c_354_n 0.00799591f $X=1.01 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A1_M1002_g N_VPWR_c_363_n 0.0046653f $X=0.59 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A1_M1003_g N_A_55_47#_c_534_n 0.0130573f $X=0.61 $Y=0.56 $X2=0 $Y2=0
cc_110 N_A1_M1016_g N_A_55_47#_c_534_n 0.0125178f $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A1_c_96_n N_A_55_47#_c_534_n 0.0390078f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_c_97_n N_A_55_47#_c_534_n 0.00212133f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A1_c_96_n N_A_55_47#_c_530_n 0.0335801f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A1_c_97_n N_A_55_47#_c_530_n 0.00111409f $X=1.03 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A1_M1003_g N_VGND_c_597_n 0.00856801f $X=0.61 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A1_M1016_g N_VGND_c_597_n 0.00685342f $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A1_M1016_g N_VGND_c_598_n 5.54209e-19 $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_118 N_A1_M1016_g N_VGND_c_599_n 0.00341689f $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A1_M1003_g N_VGND_c_601_n 0.00513114f $X=0.61 $Y=0.56 $X2=0 $Y2=0
cc_120 N_A1_M1016_g N_VGND_c_601_n 0.00405445f $X=1.03 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A1_M1003_g N_VGND_c_602_n 0.00341689f $X=0.61 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A2_M1018_g N_A3_M1013_g 0.0251781f $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_123 A2 N_A3_c_186_n 0.00210498f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A2_c_137_n N_A3_c_186_n 0.0163247f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_125 A2 A3 0.0230853f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_126 N_A2_M1006_g N_A_51_297#_c_319_n 0.0156313f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A2_M1010_g N_A_51_297#_c_319_n 0.0145015f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_128 A2 N_A_51_297#_c_319_n 0.0573518f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_129 N_A2_c_137_n N_A_51_297#_c_319_n 6.6998e-19 $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_130 A2 N_A_51_297#_c_321_n 0.00224209f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_131 N_A2_M1006_g N_VPWR_c_355_n 0.00130728f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A2_M1006_g N_VPWR_c_360_n 0.00539841f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A2_M1010_g N_VPWR_c_360_n 0.00357835f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A2_M1006_g N_VPWR_c_354_n 0.00969144f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A2_M1010_g N_VPWR_c_354_n 0.0066022f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A2_M1006_g N_A_301_297#_c_425_n 0.0045641f $X=1.43 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A2_M1010_g N_A_301_297#_c_425_n 0.0103247f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A2_M1010_g N_A_301_297#_c_424_n 0.0101161f $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A2_M1006_g N_A_301_297#_c_428_n 0.00202057f $X=1.43 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A2_M1010_g N_A_301_297#_c_428_n 7.04098e-19 $X=1.85 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A2_M1010_g N_Y_c_454_n 7.60605e-19 $X=1.85 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A2_M1009_g N_A_55_47#_c_540_n 0.0125777f $X=1.45 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A2_M1018_g N_A_55_47#_c_540_n 0.0125777f $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_144 A2 N_A_55_47#_c_540_n 0.0408564f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A2_c_137_n N_A_55_47#_c_540_n 0.00212133f $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_146 A2 N_A_55_47#_c_531_n 0.00388473f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A2_c_137_n N_A_55_47#_c_531_n 2.09233e-19 $X=1.87 $Y=1.16 $X2=0 $Y2=0
cc_148 A2 N_A_55_47#_c_532_n 0.0132419f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A2_M1009_g N_VGND_c_597_n 5.54209e-19 $X=1.45 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A2_M1009_g N_VGND_c_598_n 0.00685342f $X=1.45 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A2_M1018_g N_VGND_c_598_n 0.00684321f $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A2_M1009_g N_VGND_c_599_n 0.00341689f $X=1.45 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A2_M1009_g N_VGND_c_601_n 0.00405445f $X=1.45 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A2_M1018_g N_VGND_c_601_n 0.00405445f $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A2_M1018_g N_VGND_c_604_n 0.00341689f $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A2_M1018_g N_VGND_c_605_n 5.71356e-19 $X=1.87 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A3_M1014_g N_B1_M1005_g 0.0252561f $X=3.15 $Y=0.56 $X2=0 $Y2=0
cc_158 N_A3_M1001_g N_B1_M1011_g 0.0281127f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_159 A3 N_B1_c_234_n 0.0154797f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A3_c_188_n N_B1_c_234_n 0.00265179f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A3_c_188_n N_B1_c_235_n 0.0183137f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A3_M1000_g N_A_51_297#_c_319_n 7.60605e-19 $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A3_c_186_n N_A_51_297#_c_319_n 3.22569e-19 $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A3_M1001_g N_VPWR_c_356_n 0.00136224f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A3_M1000_g N_VPWR_c_360_n 0.00357835f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A3_M1001_g N_VPWR_c_360_n 0.00539841f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A3_M1000_g N_VPWR_c_354_n 0.0066022f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A3_M1001_g N_VPWR_c_354_n 0.00969144f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A3_M1000_g N_A_301_297#_c_424_n 0.0108202f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A3_M1001_g N_A_301_297#_c_424_n 0.00202057f $X=3.21 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A3_M1000_g N_A_301_297#_c_432_n 0.0103247f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A3_M1001_g N_A_301_297#_c_432_n 0.0045641f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A3_M1000_g N_Y_c_462_n 0.0145015f $X=2.79 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A3_M1001_g N_Y_c_462_n 0.0174971f $X=3.21 $Y=1.985 $X2=0 $Y2=0
cc_175 A3 N_Y_c_462_n 0.027079f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A3_c_188_n N_Y_c_462_n 6.11033e-19 $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_177 A3 N_Y_c_454_n 0.0209598f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A3_c_187_n N_Y_c_454_n 0.00183712f $X=2.715 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A3_M1013_g N_A_55_47#_c_547_n 0.0177692f $X=2.29 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A3_M1014_g N_A_55_47#_c_547_n 0.0168817f $X=3.15 $Y=0.56 $X2=0 $Y2=0
cc_181 A3 N_A_55_47#_c_547_n 0.0511266f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A3_c_187_n N_A_55_47#_c_547_n 0.013084f $X=2.715 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A3_c_188_n N_A_55_47#_c_533_n 2.77978e-19 $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A3_M1013_g N_VGND_c_598_n 5.53786e-19 $X=2.29 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A3_M1014_g N_VGND_c_600_n 0.00341689f $X=3.15 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A3_M1013_g N_VGND_c_601_n 0.0040385f $X=2.29 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A3_M1014_g N_VGND_c_601_n 0.0040385f $X=3.15 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A3_M1013_g N_VGND_c_604_n 0.00341689f $X=2.29 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A3_M1013_g N_VGND_c_605_n 0.00814926f $X=2.29 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A3_M1014_g N_VGND_c_605_n 0.0093743f $X=3.15 $Y=0.56 $X2=0 $Y2=0
cc_191 N_B1_M1015_g N_C1_M1004_g 0.0186128f $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B1_c_235_n N_C1_c_279_n 0.0186128f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B1_M1011_g N_VPWR_c_356_n 0.0127148f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_194 N_B1_M1015_g N_VPWR_c_356_n 0.0119337f $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_M1015_g N_VPWR_c_357_n 5.82599e-19 $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1015_g N_VPWR_c_358_n 0.0046653f $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_M1011_g N_VPWR_c_360_n 0.0046653f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_198 N_B1_M1011_g N_VPWR_c_354_n 0.00799591f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B1_M1015_g N_VPWR_c_354_n 0.0083134f $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_M1011_g N_Y_c_468_n 0.0176306f $X=3.63 $Y=1.985 $X2=0 $Y2=0
cc_201 N_B1_M1015_g N_Y_c_468_n 0.0222094f $X=4.39 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B1_c_234_n N_Y_c_468_n 0.0612929f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B1_c_235_n N_Y_c_468_n 0.00292457f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B1_c_234_n N_Y_c_455_n 0.011615f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B1_M1008_g Y 0.0037137f $X=3.99 $Y=0.56 $X2=0 $Y2=0
cc_206 N_B1_c_234_n Y 0.0217486f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B1_c_235_n Y 0.00843505f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B1_M1005_g N_A_55_47#_c_529_n 0.0125926f $X=3.57 $Y=0.56 $X2=0 $Y2=0
cc_209 N_B1_M1008_g N_A_55_47#_c_529_n 0.00994985f $X=3.99 $Y=0.56 $X2=0 $Y2=0
cc_210 N_B1_c_234_n N_A_55_47#_c_529_n 0.0607972f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B1_c_235_n N_A_55_47#_c_529_n 0.0101665f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_212 N_B1_c_234_n N_A_55_47#_c_533_n 0.00646562f $X=4 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B1_M1005_g N_VGND_c_600_n 0.00413993f $X=3.57 $Y=0.56 $X2=0 $Y2=0
cc_214 N_B1_M1008_g N_VGND_c_600_n 0.00357877f $X=3.99 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B1_M1005_g N_VGND_c_601_n 0.00578258f $X=3.57 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B1_M1008_g N_VGND_c_601_n 0.00660224f $X=3.99 $Y=0.56 $X2=0 $Y2=0
cc_217 N_B1_M1005_g N_VGND_c_605_n 0.00127196f $X=3.57 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B1_M1005_g N_A_729_47#_c_677_n 0.00304023f $X=3.57 $Y=0.56 $X2=0 $Y2=0
cc_219 N_B1_M1008_g N_A_729_47#_c_677_n 0.0120413f $X=3.99 $Y=0.56 $X2=0 $Y2=0
cc_220 N_B1_c_235_n N_A_729_47#_c_677_n 0.00263842f $X=4.39 $Y=1.16 $X2=0 $Y2=0
cc_221 N_C1_M1004_g N_VPWR_c_356_n 5.94824e-19 $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_222 N_C1_M1004_g N_VPWR_c_357_n 0.0108501f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_223 N_C1_M1012_g N_VPWR_c_357_n 0.0123094f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_224 N_C1_M1004_g N_VPWR_c_358_n 0.0046653f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_225 N_C1_M1012_g N_VPWR_c_361_n 0.0046653f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_226 N_C1_M1004_g N_VPWR_c_354_n 0.0083134f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_227 N_C1_M1012_g N_VPWR_c_354_n 0.00907261f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_228 N_C1_M1004_g N_Y_c_456_n 0.0121922f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_229 N_C1_M1012_g N_Y_c_456_n 0.0170699f $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_230 C1 N_Y_c_456_n 0.0611835f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_231 N_C1_c_279_n N_Y_c_456_n 6.15477e-19 $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_232 N_C1_c_280_n N_Y_c_456_n 0.0019356f $X=5.59 $Y=1.16 $X2=0 $Y2=0
cc_233 N_C1_M1007_g N_Y_c_450_n 0.0106243f $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_234 N_C1_M1017_g N_Y_c_450_n 0.0139502f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_235 C1 N_Y_c_450_n 0.0579902f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_236 N_C1_c_279_n N_Y_c_450_n 0.00212133f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_237 N_C1_c_280_n N_Y_c_450_n 0.00552704f $X=5.59 $Y=1.16 $X2=0 $Y2=0
cc_238 N_C1_M1004_g Y 0.00603173f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_239 N_C1_M1007_g Y 0.00534223f $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_240 N_C1_M1012_g Y 8.71561e-19 $X=5.37 $Y=1.985 $X2=0 $Y2=0
cc_241 N_C1_M1017_g Y 6.70696e-19 $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_242 C1 Y 0.0207724f $X=5.665 $Y=1.105 $X2=0 $Y2=0
cc_243 N_C1_c_279_n Y 0.00989091f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_244 N_C1_M1004_g Y 0.00666195f $X=4.95 $Y=1.985 $X2=0 $Y2=0
cc_245 N_C1_M1007_g N_Y_c_453_n 6.84149e-19 $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_246 N_C1_M1007_g N_VGND_c_600_n 0.00357877f $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_247 N_C1_M1017_g N_VGND_c_600_n 0.00413993f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_248 N_C1_M1007_g N_VGND_c_601_n 0.00660224f $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_249 N_C1_M1017_g N_VGND_c_601_n 0.0068458f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_250 N_C1_M1007_g N_A_729_47#_c_677_n 0.0120405f $X=4.97 $Y=0.56 $X2=0 $Y2=0
cc_251 N_C1_M1017_g N_A_729_47#_c_677_n 0.00316853f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A_51_297#_c_322_n N_VPWR_M1002_d 0.00315342f $X=1.135 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_253 N_A_51_297#_c_322_n N_VPWR_c_355_n 0.017435f $X=1.135 $Y=1.605 $X2=0
+ $Y2=0
cc_254 N_A_51_297#_c_337_p N_VPWR_c_360_n 0.0113958f $X=1.22 $Y=1.815 $X2=0
+ $Y2=0
cc_255 N_A_51_297#_M1002_s N_VPWR_c_354_n 0.00387172f $X=0.255 $Y=1.485 $X2=0
+ $Y2=0
cc_256 N_A_51_297#_M1019_s N_VPWR_c_354_n 0.00570907f $X=1.085 $Y=1.485 $X2=0
+ $Y2=0
cc_257 N_A_51_297#_M1010_d N_VPWR_c_354_n 0.00210147f $X=1.925 $Y=1.485 $X2=0
+ $Y2=0
cc_258 N_A_51_297#_c_317_n N_VPWR_c_354_n 0.0145574f $X=0.38 $Y=1.815 $X2=0
+ $Y2=0
cc_259 N_A_51_297#_c_337_p N_VPWR_c_354_n 0.00646998f $X=1.22 $Y=1.815 $X2=0
+ $Y2=0
cc_260 N_A_51_297#_c_317_n N_VPWR_c_363_n 0.0266045f $X=0.38 $Y=1.815 $X2=0
+ $Y2=0
cc_261 N_A_51_297#_c_319_n N_A_301_297#_M1006_s 0.00315342f $X=1.975 $Y=1.605
+ $X2=-0.19 $Y2=1.305
cc_262 N_A_51_297#_c_319_n N_A_301_297#_c_425_n 0.0171917f $X=1.975 $Y=1.605
+ $X2=0 $Y2=0
cc_263 N_A_51_297#_M1010_d N_A_301_297#_c_424_n 0.00480843f $X=1.925 $Y=1.485
+ $X2=0 $Y2=0
cc_264 N_A_51_297#_c_319_n N_A_301_297#_c_424_n 0.0030597f $X=1.975 $Y=1.605
+ $X2=0 $Y2=0
cc_265 N_A_51_297#_c_320_n N_A_301_297#_c_424_n 0.0184655f $X=2.1 $Y=1.725 $X2=0
+ $Y2=0
cc_266 N_A_51_297#_c_319_n N_Y_c_454_n 0.0207751f $X=1.975 $Y=1.605 $X2=0 $Y2=0
cc_267 N_A_51_297#_c_320_n Y 0.0294591f $X=2.1 $Y=1.725 $X2=0 $Y2=0
cc_268 N_A_51_297#_c_319_n N_A_55_47#_c_547_n 0.00123599f $X=1.975 $Y=1.605
+ $X2=0 $Y2=0
cc_269 N_A_51_297#_c_321_n N_A_55_47#_c_531_n 0.00404483f $X=1.22 $Y=1.605 $X2=0
+ $Y2=0
cc_270 N_A_51_297#_c_319_n N_A_55_47#_c_532_n 2.24764e-19 $X=1.975 $Y=1.605
+ $X2=0 $Y2=0
cc_271 N_VPWR_c_354_n N_A_301_297#_M1006_s 0.00215201f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_272 N_VPWR_c_354_n N_A_301_297#_M1000_s 0.00215201f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_360_n N_A_301_297#_c_424_n 0.0807156f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_354_n N_A_301_297#_c_424_n 0.0494971f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_360_n N_A_301_297#_c_428_n 0.0188514f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_354_n N_A_301_297#_c_428_n 0.0122326f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_354_n N_Y_M1000_d 0.00210147f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_354_n N_Y_M1001_d 0.00570907f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_354_n N_Y_M1015_d 0.00684166f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_354_n N_Y_M1012_d 0.00387172f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_360_n N_Y_c_500_n 0.0113958f $X=3.675 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_354_n N_Y_c_500_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_M1011_s N_Y_c_468_n 0.0129956f $X=3.705 $Y=1.485 $X2=0 $Y2=0
cc_284 N_VPWR_c_356_n N_Y_c_468_n 0.0457545f $X=4.18 $Y=2.02 $X2=0 $Y2=0
cc_285 N_VPWR_c_358_n N_Y_c_504_n 0.0212407f $X=4.995 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_354_n N_Y_c_504_n 0.0118616f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_M1004_s N_Y_c_456_n 0.00312111f $X=5.025 $Y=1.485 $X2=0 $Y2=0
cc_288 N_VPWR_c_357_n N_Y_c_456_n 0.017435f $X=5.16 $Y=2.02 $X2=0 $Y2=0
cc_289 N_VPWR_c_361_n N_Y_c_460_n 0.0280384f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_c_354_n N_Y_c_460_n 0.0153277f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_291 N_A_301_297#_c_424_n N_Y_M1000_d 0.00480843f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_292 N_A_301_297#_M1000_s N_Y_c_462_n 0.00312111f $X=2.865 $Y=1.485 $X2=0
+ $Y2=0
cc_293 N_A_301_297#_c_424_n N_Y_c_462_n 0.0030597f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_294 N_A_301_297#_c_432_n N_Y_c_462_n 0.0171917f $X=3 $Y=2.02 $X2=0 $Y2=0
cc_295 N_A_301_297#_c_424_n Y 0.0184655f $X=2.835 $Y=2.38 $X2=0 $Y2=0
cc_296 N_Y_c_462_n N_A_55_47#_c_547_n 0.00368425f $X=3.335 $Y=1.605 $X2=0 $Y2=0
cc_297 N_Y_c_453_n N_A_55_47#_c_529_n 0.0213627f $X=4.735 $Y=0.885 $X2=0 $Y2=0
cc_298 N_Y_c_462_n N_A_55_47#_c_533_n 0.00103922f $X=3.335 $Y=1.605 $X2=0 $Y2=0
cc_299 N_Y_c_455_n N_A_55_47#_c_533_n 9.19224e-19 $X=3.42 $Y=1.605 $X2=0 $Y2=0
cc_300 N_Y_c_450_n N_VGND_c_600_n 0.00236914f $X=5.515 $Y=0.77 $X2=0 $Y2=0
cc_301 Y N_VGND_c_600_n 0.0264549f $X=5.665 $Y=0.425 $X2=0 $Y2=0
cc_302 N_Y_M1007_d N_VGND_c_601_n 0.00226545f $X=4.615 $Y=0.235 $X2=0 $Y2=0
cc_303 N_Y_M1017_d N_VGND_c_601_n 0.00229009f $X=5.465 $Y=0.235 $X2=0 $Y2=0
cc_304 N_Y_c_450_n N_VGND_c_601_n 0.00497798f $X=5.515 $Y=0.77 $X2=0 $Y2=0
cc_305 Y N_VGND_c_601_n 0.0145283f $X=5.665 $Y=0.425 $X2=0 $Y2=0
cc_306 N_Y_c_450_n N_A_729_47#_M1007_s 0.0030829f $X=5.515 $Y=0.77 $X2=0 $Y2=0
cc_307 N_Y_M1007_d N_A_729_47#_c_677_n 0.00576876f $X=4.615 $Y=0.235 $X2=0 $Y2=0
cc_308 N_Y_c_450_n N_A_729_47#_c_677_n 0.0220062f $X=5.515 $Y=0.77 $X2=0 $Y2=0
cc_309 N_Y_c_453_n N_A_729_47#_c_677_n 0.0239232f $X=4.735 $Y=0.885 $X2=0 $Y2=0
cc_310 N_A_55_47#_c_534_n N_VGND_M1003_s 0.00307912f $X=1.155 $Y=0.77 $X2=-0.19
+ $Y2=-0.24
cc_311 N_A_55_47#_c_540_n N_VGND_M1009_d 0.00307912f $X=1.995 $Y=0.77 $X2=0
+ $Y2=0
cc_312 N_A_55_47#_c_547_n N_VGND_M1013_s 0.0155957f $X=3.275 $Y=0.77 $X2=0 $Y2=0
cc_313 N_A_55_47#_c_534_n N_VGND_c_597_n 0.0163853f $X=1.155 $Y=0.77 $X2=0 $Y2=0
cc_314 N_A_55_47#_c_540_n N_VGND_c_598_n 0.0163853f $X=1.995 $Y=0.77 $X2=0 $Y2=0
cc_315 N_A_55_47#_c_534_n N_VGND_c_599_n 0.00235985f $X=1.155 $Y=0.77 $X2=0
+ $Y2=0
cc_316 N_A_55_47#_c_570_p N_VGND_c_599_n 0.0113346f $X=1.24 $Y=0.655 $X2=0 $Y2=0
cc_317 N_A_55_47#_c_540_n N_VGND_c_599_n 0.00235985f $X=1.995 $Y=0.77 $X2=0
+ $Y2=0
cc_318 N_A_55_47#_c_547_n N_VGND_c_600_n 0.00235985f $X=3.275 $Y=0.77 $X2=0
+ $Y2=0
cc_319 N_A_55_47#_c_573_p N_VGND_c_600_n 0.0113346f $X=3.36 $Y=0.655 $X2=0 $Y2=0
cc_320 N_A_55_47#_c_529_n N_VGND_c_600_n 0.00236914f $X=4.2 $Y=0.76 $X2=0 $Y2=0
cc_321 N_A_55_47#_M1003_d N_VGND_c_601_n 0.00229009f $X=0.275 $Y=0.235 $X2=0
+ $Y2=0
cc_322 N_A_55_47#_M1016_d N_VGND_c_601_n 0.00254582f $X=1.105 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_55_47#_M1018_s N_VGND_c_601_n 0.00254582f $X=1.945 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_A_55_47#_M1014_d N_VGND_c_601_n 0.00254582f $X=3.225 $Y=0.235 $X2=0
+ $Y2=0
cc_325 N_A_55_47#_M1008_d N_VGND_c_601_n 0.00226545f $X=4.065 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_55_47#_c_534_n N_VGND_c_601_n 0.00985588f $X=1.155 $Y=0.77 $X2=0
+ $Y2=0
cc_327 N_A_55_47#_c_570_p N_VGND_c_601_n 0.00645703f $X=1.24 $Y=0.655 $X2=0
+ $Y2=0
cc_328 N_A_55_47#_c_540_n N_VGND_c_601_n 0.00984999f $X=1.995 $Y=0.77 $X2=0
+ $Y2=0
cc_329 N_A_55_47#_c_583_p N_VGND_c_601_n 0.00645703f $X=2.08 $Y=0.655 $X2=0
+ $Y2=0
cc_330 N_A_55_47#_c_547_n N_VGND_c_601_n 0.0117336f $X=3.275 $Y=0.77 $X2=0 $Y2=0
cc_331 N_A_55_47#_c_573_p N_VGND_c_601_n 0.00645703f $X=3.36 $Y=0.655 $X2=0
+ $Y2=0
cc_332 N_A_55_47#_c_529_n N_VGND_c_601_n 0.00564817f $X=4.2 $Y=0.76 $X2=0 $Y2=0
cc_333 N_A_55_47#_c_530_n N_VGND_c_601_n 0.015297f $X=0.4 $Y=0.56 $X2=0 $Y2=0
cc_334 N_A_55_47#_c_534_n N_VGND_c_602_n 0.00235985f $X=1.155 $Y=0.77 $X2=0
+ $Y2=0
cc_335 N_A_55_47#_c_530_n N_VGND_c_602_n 0.0278806f $X=0.4 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A_55_47#_c_540_n N_VGND_c_604_n 0.00235985f $X=1.995 $Y=0.77 $X2=0
+ $Y2=0
cc_337 N_A_55_47#_c_583_p N_VGND_c_604_n 0.0113346f $X=2.08 $Y=0.655 $X2=0 $Y2=0
cc_338 N_A_55_47#_c_547_n N_VGND_c_604_n 0.00235985f $X=3.275 $Y=0.77 $X2=0
+ $Y2=0
cc_339 N_A_55_47#_c_547_n N_VGND_c_605_n 0.0507112f $X=3.275 $Y=0.77 $X2=0 $Y2=0
cc_340 N_A_55_47#_c_529_n N_A_729_47#_M1005_s 0.0030829f $X=4.2 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_341 N_A_55_47#_M1008_d N_A_729_47#_c_677_n 0.00553375f $X=4.065 $Y=0.235
+ $X2=0 $Y2=0
cc_342 N_A_55_47#_c_529_n N_A_729_47#_c_677_n 0.0425011f $X=4.2 $Y=0.76 $X2=0
+ $Y2=0
cc_343 N_VGND_c_601_n N_A_729_47#_M1005_s 0.00215227f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_344 N_VGND_c_601_n N_A_729_47#_M1007_s 0.00215227f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_c_600_n N_A_729_47#_c_677_n 0.101352f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_601_n N_A_729_47#_c_677_n 0.0629356f $X=5.75 $Y=0 $X2=0 $Y2=0

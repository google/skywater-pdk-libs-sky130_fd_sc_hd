* File: sky130_fd_sc_hd__a2111o_4.pxi.spice
* Created: Thu Aug 27 13:58:44 2020
* 
x_PM_SKY130_FD_SC_HD__A2111O_4%D1 N_D1_M1005_g N_D1_c_115_n N_D1_M1000_g
+ N_D1_M1018_g N_D1_c_116_n N_D1_M1001_g D1 D1 N_D1_c_118_n
+ PM_SKY130_FD_SC_HD__A2111O_4%D1
x_PM_SKY130_FD_SC_HD__A2111O_4%C1 N_C1_M1006_g N_C1_c_154_n N_C1_M1015_g
+ N_C1_M1024_g N_C1_c_155_n N_C1_M1016_g C1 C1 C1
+ PM_SKY130_FD_SC_HD__A2111O_4%C1
x_PM_SKY130_FD_SC_HD__A2111O_4%B1 N_B1_c_203_n N_B1_M1008_g N_B1_M1004_g
+ N_B1_M1014_g N_B1_c_204_n N_B1_M1019_g B1 B1 N_B1_c_205_n
+ PM_SKY130_FD_SC_HD__A2111O_4%B1
x_PM_SKY130_FD_SC_HD__A2111O_4%A1 N_A1_c_251_n N_A1_M1010_g N_A1_M1002_g
+ N_A1_c_252_n N_A1_M1026_g N_A1_M1017_g A1 A1 N_A1_c_254_n
+ PM_SKY130_FD_SC_HD__A2111O_4%A1
x_PM_SKY130_FD_SC_HD__A2111O_4%A2 N_A2_c_296_n N_A2_M1011_g N_A2_M1003_g
+ N_A2_c_297_n N_A2_M1022_g N_A2_M1023_g A2 A2 N_A2_c_298_n N_A2_c_299_n A2
+ PM_SKY130_FD_SC_HD__A2111O_4%A2
x_PM_SKY130_FD_SC_HD__A2111O_4%A_44_47# N_A_44_47#_M1000_s N_A_44_47#_M1001_s
+ N_A_44_47#_M1016_s N_A_44_47#_M1019_d N_A_44_47#_M1026_s N_A_44_47#_M1005_d
+ N_A_44_47#_c_338_n N_A_44_47#_M1009_g N_A_44_47#_M1007_g N_A_44_47#_c_339_n
+ N_A_44_47#_M1012_g N_A_44_47#_M1013_g N_A_44_47#_c_340_n N_A_44_47#_M1020_g
+ N_A_44_47#_M1025_g N_A_44_47#_c_341_n N_A_44_47#_M1021_g N_A_44_47#_M1027_g
+ N_A_44_47#_c_342_n N_A_44_47#_c_343_n N_A_44_47#_c_365_n N_A_44_47#_c_344_n
+ N_A_44_47#_c_484_p N_A_44_47#_c_372_n N_A_44_47#_c_496_p N_A_44_47#_c_378_n
+ N_A_44_47#_c_487_p N_A_44_47#_c_345_n N_A_44_47#_c_346_n N_A_44_47#_c_355_n
+ N_A_44_47#_c_356_n N_A_44_47#_c_347_n N_A_44_47#_c_348_n N_A_44_47#_c_426_p
+ N_A_44_47#_c_375_n N_A_44_47#_c_377_n N_A_44_47#_c_349_n
+ PM_SKY130_FD_SC_HD__A2111O_4%A_44_47#
x_PM_SKY130_FD_SC_HD__A2111O_4%A_30_297# N_A_30_297#_M1005_s N_A_30_297#_M1018_s
+ N_A_30_297#_M1024_s N_A_30_297#_c_521_n N_A_30_297#_c_529_n
+ N_A_30_297#_c_522_n N_A_30_297#_c_523_n N_A_30_297#_c_524_n
+ N_A_30_297#_c_525_n N_A_30_297#_c_551_p PM_SKY130_FD_SC_HD__A2111O_4%A_30_297#
x_PM_SKY130_FD_SC_HD__A2111O_4%A_285_297# N_A_285_297#_M1006_d
+ N_A_285_297#_M1004_s N_A_285_297#_c_562_n N_A_285_297#_c_559_n
+ N_A_285_297#_c_560_n N_A_285_297#_c_561_n
+ PM_SKY130_FD_SC_HD__A2111O_4%A_285_297#
x_PM_SKY130_FD_SC_HD__A2111O_4%A_477_297# N_A_477_297#_M1004_d
+ N_A_477_297#_M1014_d N_A_477_297#_M1017_s N_A_477_297#_M1003_d
+ N_A_477_297#_c_595_n N_A_477_297#_c_602_n N_A_477_297#_c_596_n
+ N_A_477_297#_c_605_n N_A_477_297#_c_607_n N_A_477_297#_c_610_n
+ N_A_477_297#_c_597_n N_A_477_297#_c_598_n N_A_477_297#_c_599_n
+ N_A_477_297#_c_623_n PM_SKY130_FD_SC_HD__A2111O_4%A_477_297#
x_PM_SKY130_FD_SC_HD__A2111O_4%VPWR N_VPWR_M1002_d N_VPWR_M1003_s N_VPWR_M1023_s
+ N_VPWR_M1013_s N_VPWR_M1027_s N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n
+ N_VPWR_c_662_n N_VPWR_c_663_n N_VPWR_c_664_n N_VPWR_c_665_n VPWR
+ N_VPWR_c_666_n N_VPWR_c_667_n N_VPWR_c_668_n N_VPWR_c_669_n N_VPWR_c_670_n
+ N_VPWR_c_671_n N_VPWR_c_672_n N_VPWR_c_673_n N_VPWR_c_658_n
+ PM_SKY130_FD_SC_HD__A2111O_4%VPWR
x_PM_SKY130_FD_SC_HD__A2111O_4%X N_X_M1009_d N_X_M1020_d N_X_M1007_d N_X_M1025_d
+ N_X_c_827_p N_X_c_809_n N_X_c_783_n N_X_c_787_n N_X_c_777_n N_X_c_778_n
+ N_X_c_830_p N_X_c_813_n N_X_c_797_n N_X_c_779_n N_X_c_801_n N_X_c_780_n X X X
+ N_X_c_775_n N_X_c_781_n X PM_SKY130_FD_SC_HD__A2111O_4%X
x_PM_SKY130_FD_SC_HD__A2111O_4%VGND N_VGND_M1000_d N_VGND_M1015_d N_VGND_M1008_s
+ N_VGND_M1011_d N_VGND_M1022_d N_VGND_M1012_s N_VGND_M1021_s N_VGND_c_839_n
+ N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n
+ N_VGND_c_845_n VGND N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n
+ N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n
+ N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n N_VGND_c_858_n
+ PM_SKY130_FD_SC_HD__A2111O_4%VGND
x_PM_SKY130_FD_SC_HD__A2111O_4%A_770_47# N_A_770_47#_M1010_d N_A_770_47#_M1011_s
+ N_A_770_47#_c_974_n N_A_770_47#_c_993_n PM_SKY130_FD_SC_HD__A2111O_4%A_770_47#
cc_1 VNB N_D1_c_115_n 0.0209206f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_2 VNB N_D1_c_116_n 0.0161053f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB D1 0.0177638f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_D1_c_118_n 0.0604475f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_5 VNB N_C1_c_154_n 0.0165962f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.995
cc_6 VNB N_C1_c_155_n 0.0566914f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_7 VNB C1 0.0178525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_c_203_n 0.0214978f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_9 VNB N_B1_c_204_n 0.0883873f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_10 VNB N_B1_c_205_n 0.00770357f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_11 VNB N_A1_c_251_n 0.0164509f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_12 VNB N_A1_c_252_n 0.0220764f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.325
cc_13 VNB A1 0.00144351f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_14 VNB N_A1_c_254_n 0.0472495f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.16
cc_15 VNB N_A2_c_296_n 0.0211871f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_16 VNB N_A2_c_297_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.325
cc_17 VNB N_A2_c_298_n 0.00771343f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_18 VNB N_A2_c_299_n 0.0465417f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_19 VNB N_A_44_47#_c_338_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_20 VNB N_A_44_47#_c_339_n 0.0160063f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_21 VNB N_A_44_47#_c_340_n 0.0160024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_44_47#_c_341_n 0.0184169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_44_47#_c_342_n 0.0146667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_44_47#_c_343_n 9.95532e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_44_47#_c_344_n 0.00743543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_44_47#_c_345_n 0.00828684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_44_47#_c_346_n 0.00209911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_44_47#_c_347_n 4.52616e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_44_47#_c_348_n 0.00376107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_44_47#_c_349_n 0.0671388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_658_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_775_n 0.00789458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB X 0.0247392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_839_n 4.06069e-19 $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_35 VNB N_VGND_c_840_n 0.00207523f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_841_n 0.00495694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_842_n 3.08203e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_843_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_844_n 0.0105624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_845_n 0.0119016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_846_n 0.0133254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_847_n 0.0343441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_848_n 0.0120336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_849_n 0.0121761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_850_n 0.0114125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_851_n 0.0216742f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_852_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_853_n 0.0125382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_854_n 0.017302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_855_n 0.00516648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_856_n 0.00436447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_857_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_858_n 0.376913f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_770_47#_c_974_n 0.00850366f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.56
cc_55 VPB N_D1_M1005_g 0.0213135f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_56 VPB N_D1_M1018_g 0.0183803f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_57 VPB D1 0.0143026f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_58 VPB N_D1_c_118_n 0.0156114f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_59 VPB N_C1_M1006_g 0.0190953f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_60 VPB N_C1_M1024_g 0.0257893f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_61 VPB N_C1_c_155_n 0.00828698f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_62 VPB N_B1_M1004_g 0.025792f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.56
cc_63 VPB N_B1_M1014_g 0.0213002f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.985
cc_64 VPB N_B1_c_204_n 0.0218635f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_65 VPB N_A1_M1002_g 0.0198672f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.56
cc_66 VPB N_A1_M1017_g 0.0241397f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_67 VPB N_A1_c_254_n 0.0117131f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.16
cc_68 VPB N_A2_M1003_g 0.0240916f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.56
cc_69 VPB N_A2_M1023_g 0.0183397f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_70 VPB N_A2_c_299_n 0.00459586f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_71 VPB N_A_44_47#_M1007_g 0.0178715f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_72 VPB N_A_44_47#_M1013_g 0.0183387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_44_47#_M1025_g 0.0183253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_44_47#_M1027_g 0.0211356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_44_47#_c_345_n 0.00318233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_44_47#_c_355_n 0.021905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_44_47#_c_356_n 5.01553e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_44_47#_c_347_n 0.00129437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_44_47#_c_349_n 0.0109578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_30_297#_c_521_n 0.019062f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_81 VPB N_A_30_297#_c_522_n 0.00745908f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_82 VPB N_A_30_297#_c_523_n 0.00218211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_30_297#_c_524_n 0.00185888f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_84 VPB N_A_30_297#_c_525_n 0.00486432f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_85 VPB N_A_285_297#_c_559_n 0.0155311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_285_297#_c_560_n 0.00229485f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_87 VPB N_A_285_297#_c_561_n 0.00181605f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_88 VPB N_A_477_297#_c_595_n 0.00478541f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_89 VPB N_A_477_297#_c_596_n 0.00184411f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_477_297#_c_597_n 0.00565166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_477_297#_c_598_n 0.00670759f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.53
cc_92 VPB N_A_477_297#_c_599_n 7.45409e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_659_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_660_n 0.0147821f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_95 VPB N_VPWR_c_661_n 0.00489721f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_96 VPB N_VPWR_c_662_n 3.08203e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_663_n 3.0911e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_664_n 0.0106587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_665_n 0.0293229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_666_n 0.0908597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_667_n 0.0121874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_668_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_669_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_670_n 0.00436664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_671_n 0.00516774f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_672_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_673_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_658_n 0.056562f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_X_c_777_n 0.00336484f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_110 VPB N_X_c_778_n 0.00174166f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.16
cc_111 VPB N_X_c_779_n 0.0016327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_X_c_780_n 0.00158547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_X_c_781_n 0.00854386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB X 0.00808214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 N_D1_M1018_g N_C1_M1006_g 0.0110356f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_116 N_D1_c_116_n N_C1_c_154_n 0.0237277f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_117 N_D1_c_118_n N_C1_c_155_n 0.020847f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_118 N_D1_c_116_n C1 7.45681e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_119 N_D1_c_118_n C1 0.00571939f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_120 N_D1_M1005_g N_A_44_47#_c_343_n 0.016299f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_121 N_D1_c_115_n N_A_44_47#_c_343_n 0.010679f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_122 N_D1_M1018_g N_A_44_47#_c_343_n 0.0113575f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_123 N_D1_c_116_n N_A_44_47#_c_343_n 0.00295823f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_124 D1 N_A_44_47#_c_343_n 0.043706f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_125 N_D1_c_118_n N_A_44_47#_c_343_n 0.0228904f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_126 N_D1_c_116_n N_A_44_47#_c_365_n 0.01521f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_127 N_D1_c_115_n N_A_44_47#_c_344_n 0.013731f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_128 D1 N_A_44_47#_c_344_n 0.0157043f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_129 N_D1_c_118_n N_A_44_47#_c_344_n 0.00527592f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_130 D1 N_A_30_297#_M1005_s 0.00368016f $X=0.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_131 D1 N_A_30_297#_c_521_n 0.0223083f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_132 N_D1_c_118_n N_A_30_297#_c_521_n 0.00104271f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_133 N_D1_M1005_g N_A_30_297#_c_529_n 0.0115032f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_134 N_D1_M1018_g N_A_30_297#_c_529_n 0.0115032f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_135 N_D1_M1018_g N_A_30_297#_c_523_n 2.13358e-19 $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_136 N_D1_M1005_g N_VPWR_c_666_n 0.00357877f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_137 N_D1_M1018_g N_VPWR_c_666_n 0.00357877f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_138 N_D1_M1005_g N_VPWR_c_658_n 0.00622544f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_139 N_D1_M1018_g N_VPWR_c_658_n 0.00530427f $X=0.92 $Y=1.985 $X2=0 $Y2=0
cc_140 N_D1_c_115_n N_VGND_c_839_n 0.00810303f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_141 N_D1_c_116_n N_VGND_c_839_n 0.00654948f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_142 N_D1_c_116_n N_VGND_c_846_n 0.00353537f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_143 N_D1_c_115_n N_VGND_c_851_n 0.00353537f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_144 N_D1_c_115_n N_VGND_c_858_n 0.00511674f $X=0.56 $Y=0.995 $X2=0 $Y2=0
cc_145 N_D1_c_116_n N_VGND_c_858_n 0.00413843f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_146 N_C1_c_155_n N_B1_c_203_n 0.0200876f $X=1.885 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_147 C1 N_B1_c_203_n 0.0032803f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_148 N_C1_c_155_n N_B1_c_204_n 0.0153055f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_149 C1 N_B1_c_205_n 0.0275405f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_150 N_C1_c_155_n N_A_44_47#_c_343_n 0.00124417f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_151 C1 N_A_44_47#_c_343_n 0.0252463f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_152 C1 N_A_44_47#_c_365_n 0.00363231f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_153 N_C1_c_154_n N_A_44_47#_c_372_n 0.0126854f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_154 N_C1_c_155_n N_A_44_47#_c_372_n 0.0136867f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_155 C1 N_A_44_47#_c_372_n 0.0443804f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_156 N_C1_c_155_n N_A_44_47#_c_375_n 3.27228e-19 $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_157 C1 N_A_44_47#_c_375_n 0.0167451f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_158 C1 N_A_44_47#_c_377_n 0.0189301f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_159 N_C1_M1006_g N_A_30_297#_c_523_n 2.12903e-19 $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_160 C1 N_A_30_297#_c_523_n 0.0165566f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_161 N_C1_M1006_g N_A_30_297#_c_524_n 0.0115032f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_162 N_C1_M1024_g N_A_30_297#_c_524_n 0.00955545f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_163 N_C1_M1006_g N_A_285_297#_c_562_n 0.00537055f $X=1.35 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_C1_M1024_g N_A_285_297#_c_562_n 0.0111682f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_165 N_C1_M1024_g N_A_285_297#_c_559_n 0.011287f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_166 N_C1_c_155_n N_A_285_297#_c_559_n 0.00416365f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_167 C1 N_A_285_297#_c_559_n 0.0417221f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_168 N_C1_M1006_g N_A_285_297#_c_560_n 0.00242244f $X=1.35 $Y=1.985 $X2=0
+ $Y2=0
cc_169 N_C1_M1024_g N_A_285_297#_c_560_n 0.00108107f $X=1.78 $Y=1.985 $X2=0
+ $Y2=0
cc_170 N_C1_c_155_n N_A_285_297#_c_560_n 0.00270934f $X=1.885 $Y=0.995 $X2=0
+ $Y2=0
cc_171 C1 N_A_285_297#_c_560_n 0.0274556f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_172 N_C1_M1006_g N_VPWR_c_666_n 0.00357877f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_173 N_C1_M1024_g N_VPWR_c_666_n 0.00357877f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_174 N_C1_M1006_g N_VPWR_c_658_n 0.00530427f $X=1.35 $Y=1.985 $X2=0 $Y2=0
cc_175 N_C1_M1024_g N_VPWR_c_658_n 0.00657863f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_176 N_C1_c_154_n N_VGND_c_839_n 5.20137e-19 $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_177 N_C1_c_154_n N_VGND_c_840_n 0.00163938f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_178 N_C1_c_155_n N_VGND_c_840_n 0.00658563f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_179 N_C1_c_154_n N_VGND_c_846_n 0.00422112f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C1_c_155_n N_VGND_c_853_n 0.00337001f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_181 N_C1_c_155_n N_VGND_c_854_n 5.00863e-19 $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_182 N_C1_c_154_n N_VGND_c_858_n 0.00569962f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C1_c_155_n N_VGND_c_858_n 0.00408452f $X=1.885 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B1_c_204_n N_A1_c_251_n 0.0120745f $X=3.34 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_185 N_B1_M1014_g N_A1_M1002_g 0.0224164f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_186 N_B1_M1014_g N_A1_c_254_n 2.67212e-19 $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B1_c_204_n N_A1_c_254_n 0.0120745f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_188 N_B1_c_203_n N_A_44_47#_c_378_n 0.0166956f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_204_n N_A_44_47#_c_378_n 0.0208082f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_205_n N_A_44_47#_c_378_n 0.0592706f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B1_M1014_g N_A_44_47#_c_345_n 0.00265494f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B1_c_204_n N_A_44_47#_c_345_n 0.00610402f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B1_c_205_n N_A_44_47#_c_345_n 0.0212272f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B1_M1014_g N_A_44_47#_c_356_n 0.00201573f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_195 N_B1_M1004_g N_A_30_297#_c_524_n 3.51118e-19 $X=2.72 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B1_M1004_g N_A_285_297#_c_559_n 0.012627f $X=2.72 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B1_c_204_n N_A_285_297#_c_559_n 0.00993607f $X=3.34 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_B1_c_205_n N_A_285_297#_c_559_n 0.0289465f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_M1014_g N_A_285_297#_c_561_n 0.0109782f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_200 N_B1_c_204_n N_A_285_297#_c_561_n 0.00241745f $X=3.34 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_B1_c_205_n N_A_285_297#_c_561_n 0.0212768f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_M1004_g N_A_477_297#_c_595_n 0.00715486f $X=2.72 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_B1_M1014_g N_A_477_297#_c_595_n 4.62664e-19 $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_B1_M1004_g N_A_477_297#_c_602_n 0.00835057f $X=2.72 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_B1_M1014_g N_A_477_297#_c_602_n 0.0143317f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B1_M1004_g N_A_477_297#_c_596_n 0.00111862f $X=2.72 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_B1_M1014_g N_A_477_297#_c_605_n 0.00219939f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_B1_c_204_n N_A_477_297#_c_605_n 0.0033085f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_209 N_B1_M1014_g N_A_477_297#_c_607_n 0.00399765f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_B1_M1014_g N_VPWR_c_659_n 9.56281e-19 $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B1_M1004_g N_VPWR_c_666_n 0.00357835f $X=2.72 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B1_M1014_g N_VPWR_c_666_n 0.00357877f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_VPWR_c_658_n 0.00666848f $X=2.72 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B1_M1014_g N_VPWR_c_658_n 0.00582751f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B1_c_203_n N_VGND_c_840_n 4.88702e-19 $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_204_n N_VGND_c_847_n 0.00337001f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_203_n N_VGND_c_853_n 0.00351072f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_203_n N_VGND_c_854_n 0.00804168f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_204_n N_VGND_c_854_n 0.00931815f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_c_203_n N_VGND_c_858_n 0.00421026f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_204_n N_VGND_c_858_n 0.00395417f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_222 A1 N_A2_c_298_n 0.0168838f $X=4.295 $Y=1.105 $X2=0 $Y2=0
cc_223 N_A1_c_254_n N_A2_c_298_n 8.96772e-19 $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A1_c_254_n N_A2_c_299_n 0.00952502f $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A1_c_251_n N_A_44_47#_c_345_n 0.00833994f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A1_M1002_g N_A_44_47#_c_345_n 0.00284841f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_227 A1 N_A_44_47#_c_345_n 0.01593f $X=4.295 $Y=1.105 $X2=0 $Y2=0
cc_228 N_A1_c_251_n N_A_44_47#_c_346_n 0.0120659f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A1_c_252_n N_A_44_47#_c_346_n 0.00816381f $X=4.205 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A1_M1002_g N_A_44_47#_c_355_n 0.013926f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_M1017_g N_A_44_47#_c_355_n 0.0129956f $X=4.245 $Y=1.985 $X2=0 $Y2=0
cc_232 A1 N_A_44_47#_c_355_n 0.0479065f $X=4.295 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A1_c_254_n N_A_44_47#_c_355_n 0.00861179f $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A1_M1002_g N_A_285_297#_c_561_n 8.974e-19 $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A1_M1002_g N_A_477_297#_c_602_n 0.00187224f $X=3.815 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A1_M1002_g N_A_477_297#_c_607_n 0.00617058f $X=3.815 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A1_M1002_g N_A_477_297#_c_610_n 0.013967f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A1_M1017_g N_A_477_297#_c_610_n 0.0106678f $X=4.245 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A1_M1002_g N_VPWR_c_659_n 0.00947128f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A1_M1017_g N_VPWR_c_659_n 0.00876929f $X=4.245 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A1_M1017_g N_VPWR_c_660_n 0.00364083f $X=4.245 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A1_M1017_g N_VPWR_c_661_n 0.00235472f $X=4.245 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A1_M1002_g N_VPWR_c_666_n 0.00364083f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A1_M1002_g N_VPWR_c_658_n 0.00485174f $X=3.815 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A1_M1017_g N_VPWR_c_658_n 0.00569274f $X=4.245 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A1_c_252_n N_VGND_c_841_n 0.00223149f $X=4.205 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A1_c_251_n N_VGND_c_847_n 0.00357877f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A1_c_252_n N_VGND_c_847_n 0.00357877f $X=4.205 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A1_c_251_n N_VGND_c_854_n 0.0011428f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A1_c_251_n N_VGND_c_858_n 0.00531636f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_252_n N_VGND_c_858_n 0.00657863f $X=4.205 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_251_n N_A_770_47#_c_974_n 0.00246548f $X=3.775 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A1_c_252_n N_A_770_47#_c_974_n 0.0111389f $X=4.205 $Y=0.995 $X2=0 $Y2=0
cc_254 A1 N_A_770_47#_c_974_n 0.0269595f $X=4.295 $Y=1.105 $X2=0 $Y2=0
cc_255 N_A1_c_254_n N_A_770_47#_c_974_n 0.00728549f $X=4.33 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A2_c_297_n N_A_44_47#_c_338_n 0.0223562f $X=5.615 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A2_M1023_g N_A_44_47#_M1007_g 0.0223562f $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A2_M1003_g N_A_44_47#_c_355_n 0.013045f $X=5.185 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A2_M1023_g N_A_44_47#_c_355_n 0.0167206f $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A2_c_298_n N_A_44_47#_c_355_n 0.0692718f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A2_c_299_n N_A_44_47#_c_355_n 0.00580038f $X=5.615 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A2_c_298_n N_A_44_47#_c_347_n 0.00228883f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A2_c_299_n N_A_44_47#_c_347_n 0.00415512f $X=5.615 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A2_c_298_n N_A_44_47#_c_348_n 0.0150658f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A2_c_299_n N_A_44_47#_c_348_n 0.00153605f $X=5.615 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A2_c_299_n N_A_44_47#_c_349_n 0.0223562f $X=5.615 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A2_M1003_g N_A_477_297#_c_597_n 0.00537856f $X=5.185 $Y=1.985 $X2=0
+ $Y2=0
cc_268 N_A2_M1003_g N_A_477_297#_c_598_n 0.0131142f $X=5.185 $Y=1.985 $X2=0
+ $Y2=0
cc_269 N_A2_M1003_g N_VPWR_c_661_n 0.00789963f $X=5.185 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A2_M1023_g N_VPWR_c_661_n 5.08869e-19 $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A2_M1003_g N_VPWR_c_662_n 5.76051e-19 $X=5.185 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A2_M1023_g N_VPWR_c_662_n 0.0117678f $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A2_M1003_g N_VPWR_c_667_n 0.00349488f $X=5.185 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A2_M1023_g N_VPWR_c_667_n 0.00486043f $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A2_M1003_g N_VPWR_c_658_n 0.00414757f $X=5.185 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A2_M1023_g N_VPWR_c_658_n 0.00822531f $X=5.615 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A2_c_296_n N_VGND_c_841_n 0.00758646f $X=5.185 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_297_n N_VGND_c_841_n 5.03136e-19 $X=5.615 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A2_c_296_n N_VGND_c_842_n 5.16359e-19 $X=5.185 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A2_c_297_n N_VGND_c_842_n 0.00776186f $X=5.615 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A2_c_296_n N_VGND_c_848_n 0.00337001f $X=5.185 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A2_c_297_n N_VGND_c_848_n 0.00486043f $X=5.615 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A2_c_296_n N_VGND_c_858_n 0.00393206f $X=5.185 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A2_c_297_n N_VGND_c_858_n 0.00822531f $X=5.615 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A2_c_296_n N_A_770_47#_c_974_n 0.0137822f $X=5.185 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A2_c_298_n N_A_770_47#_c_974_n 0.0373661f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A2_c_299_n N_A_770_47#_c_974_n 0.0054498f $X=5.615 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_44_47#_M1005_d N_A_30_297#_c_529_n 0.0033237f $X=0.565 $Y=1.485 $X2=0
+ $Y2=0
cc_289 N_A_44_47#_c_343_n N_A_30_297#_c_529_n 0.0159977f $X=0.705 $Y=1.67 $X2=0
+ $Y2=0
cc_290 N_A_44_47#_c_343_n N_A_30_297#_c_523_n 0.0262497f $X=0.705 $Y=1.67 $X2=0
+ $Y2=0
cc_291 N_A_44_47#_c_378_n N_A_285_297#_c_559_n 0.00416363f $X=3.465 $Y=0.71
+ $X2=0 $Y2=0
cc_292 N_A_44_47#_c_356_n N_A_285_297#_c_561_n 0.00827877f $X=3.655 $Y=1.535
+ $X2=0 $Y2=0
cc_293 N_A_44_47#_c_355_n N_A_477_297#_M1014_d 2.88223e-19 $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_294 N_A_44_47#_c_356_n N_A_477_297#_M1014_d 0.00455159f $X=3.655 $Y=1.535
+ $X2=0 $Y2=0
cc_295 N_A_44_47#_c_355_n N_A_477_297#_M1017_s 0.00277723f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_296 N_A_44_47#_c_355_n N_A_477_297#_M1003_d 0.00176773f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_297 N_A_44_47#_c_356_n N_A_477_297#_c_605_n 0.0166616f $X=3.655 $Y=1.535
+ $X2=0 $Y2=0
cc_298 N_A_44_47#_c_355_n N_A_477_297#_c_610_n 0.0349353f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_299 N_A_44_47#_c_356_n N_A_477_297#_c_610_n 3.73915e-19 $X=3.655 $Y=1.535
+ $X2=0 $Y2=0
cc_300 N_A_44_47#_c_355_n N_A_477_297#_c_598_n 0.0424858f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_301 N_A_44_47#_c_355_n N_A_477_297#_c_599_n 0.0202428f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_302 N_A_44_47#_c_355_n N_A_477_297#_c_623_n 0.0135413f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_303 N_A_44_47#_c_355_n N_VPWR_M1002_d 0.00177204f $X=5.795 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_304 N_A_44_47#_c_355_n N_VPWR_M1003_s 0.00278251f $X=5.795 $Y=1.535 $X2=0
+ $Y2=0
cc_305 N_A_44_47#_c_355_n N_VPWR_M1023_s 0.00181991f $X=5.795 $Y=1.535 $X2=0
+ $Y2=0
cc_306 N_A_44_47#_M1007_g N_VPWR_c_662_n 0.0119835f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_307 N_A_44_47#_M1013_g N_VPWR_c_662_n 6.32953e-19 $X=6.475 $Y=1.985 $X2=0
+ $Y2=0
cc_308 N_A_44_47#_c_355_n N_VPWR_c_662_n 0.0161254f $X=5.795 $Y=1.535 $X2=0
+ $Y2=0
cc_309 N_A_44_47#_c_426_p N_VPWR_c_662_n 5.32959e-19 $X=7.155 $Y=1.16 $X2=0
+ $Y2=0
cc_310 N_A_44_47#_M1007_g N_VPWR_c_663_n 6.08906e-19 $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_311 N_A_44_47#_M1013_g N_VPWR_c_663_n 0.0101993f $X=6.475 $Y=1.985 $X2=0
+ $Y2=0
cc_312 N_A_44_47#_M1025_g N_VPWR_c_663_n 0.0101993f $X=6.905 $Y=1.985 $X2=0
+ $Y2=0
cc_313 N_A_44_47#_M1027_g N_VPWR_c_663_n 6.08906e-19 $X=7.335 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_44_47#_M1025_g N_VPWR_c_665_n 6.31539e-19 $X=6.905 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_44_47#_M1027_g N_VPWR_c_665_n 0.0120712f $X=7.335 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_A_44_47#_M1007_g N_VPWR_c_668_n 0.00486043f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_A_44_47#_M1013_g N_VPWR_c_668_n 0.00486043f $X=6.475 $Y=1.985 $X2=0
+ $Y2=0
cc_318 N_A_44_47#_M1025_g N_VPWR_c_669_n 0.00486043f $X=6.905 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A_44_47#_M1027_g N_VPWR_c_669_n 0.00486043f $X=7.335 $Y=1.985 $X2=0
+ $Y2=0
cc_320 N_A_44_47#_M1005_d N_VPWR_c_658_n 0.00224864f $X=0.565 $Y=1.485 $X2=0
+ $Y2=0
cc_321 N_A_44_47#_M1007_g N_VPWR_c_658_n 0.00822531f $X=6.045 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_44_47#_M1013_g N_VPWR_c_658_n 0.00822531f $X=6.475 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_44_47#_M1025_g N_VPWR_c_658_n 0.00822531f $X=6.905 $Y=1.985 $X2=0
+ $Y2=0
cc_324 N_A_44_47#_M1027_g N_VPWR_c_658_n 0.00822531f $X=7.335 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_44_47#_c_339_n N_X_c_783_n 0.0117723f $X=6.475 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_44_47#_c_340_n N_X_c_783_n 0.0121753f $X=6.905 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_44_47#_c_426_p N_X_c_783_n 0.0270033f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_44_47#_c_349_n N_X_c_783_n 0.00230068f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_44_47#_c_426_p N_X_c_787_n 0.00958922f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_44_47#_c_349_n N_X_c_787_n 0.00240202f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_44_47#_M1013_g N_X_c_777_n 0.0165553f $X=6.475 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_44_47#_M1025_g N_X_c_777_n 0.0169607f $X=6.905 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A_44_47#_c_426_p N_X_c_777_n 0.0395183f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_44_47#_c_349_n N_X_c_777_n 0.00241175f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_44_47#_M1007_g N_X_c_778_n 8.36081e-19 $X=6.045 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_44_47#_c_355_n N_X_c_778_n 0.00700994f $X=5.795 $Y=1.535 $X2=0 $Y2=0
cc_337 N_A_44_47#_c_426_p N_X_c_778_n 0.0126488f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_338 N_A_44_47#_c_349_n N_X_c_778_n 0.00250185f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_44_47#_c_341_n N_X_c_797_n 0.0145984f $X=7.335 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_44_47#_c_426_p N_X_c_797_n 0.00386393f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_44_47#_M1027_g N_X_c_779_n 0.0172025f $X=7.335 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_44_47#_c_426_p N_X_c_779_n 0.00593347f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_44_47#_c_426_p N_X_c_801_n 0.00958922f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_44_47#_c_349_n N_X_c_801_n 0.00240202f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A_44_47#_c_426_p N_X_c_780_n 0.0126488f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_44_47#_c_349_n N_X_c_780_n 0.00250185f $X=7.335 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_44_47#_c_341_n X 0.0255817f $X=7.335 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A_44_47#_c_426_p X 0.0137867f $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A_44_47#_c_343_n N_VGND_M1000_d 4.86796e-19 $X=0.705 $Y=1.67 $X2=-0.19
+ $Y2=-0.24
cc_350 N_A_44_47#_c_344_n N_VGND_M1000_d 0.00213605f $X=0.87 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_351 N_A_44_47#_c_372_n N_VGND_M1015_d 0.00390197f $X=2.015 $Y=0.71 $X2=0
+ $Y2=0
cc_352 N_A_44_47#_c_378_n N_VGND_M1008_s 0.0181381f $X=3.465 $Y=0.71 $X2=0 $Y2=0
cc_353 N_A_44_47#_c_344_n N_VGND_c_839_n 0.0160114f $X=0.87 $Y=0.72 $X2=0 $Y2=0
cc_354 N_A_44_47#_c_372_n N_VGND_c_840_n 0.0173796f $X=2.015 $Y=0.71 $X2=0 $Y2=0
cc_355 N_A_44_47#_c_346_n N_VGND_c_841_n 0.0138867f $X=4.415 $Y=0.36 $X2=0 $Y2=0
cc_356 N_A_44_47#_c_338_n N_VGND_c_842_n 0.00712615f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_44_47#_c_339_n N_VGND_c_842_n 5.18376e-19 $X=6.475 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_44_47#_c_348_n N_VGND_c_842_n 0.00572833f $X=5.975 $Y=1.16 $X2=0
+ $Y2=0
cc_359 N_A_44_47#_c_426_p N_VGND_c_842_n 5.2302e-19 $X=7.155 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A_44_47#_c_338_n N_VGND_c_843_n 4.98572e-19 $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_361 N_A_44_47#_c_339_n N_VGND_c_843_n 0.00627457f $X=6.475 $Y=0.995 $X2=0
+ $Y2=0
cc_362 N_A_44_47#_c_340_n N_VGND_c_843_n 0.00627457f $X=6.905 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A_44_47#_c_341_n N_VGND_c_843_n 4.98572e-19 $X=7.335 $Y=0.995 $X2=0
+ $Y2=0
cc_364 N_A_44_47#_c_340_n N_VGND_c_845_n 5.0423e-19 $X=6.905 $Y=0.995 $X2=0
+ $Y2=0
cc_365 N_A_44_47#_c_341_n N_VGND_c_845_n 0.00752096f $X=7.335 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_44_47#_c_365_n N_VGND_c_846_n 0.00247598f $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_367 N_A_44_47#_c_484_p N_VGND_c_846_n 0.0136939f $X=1.205 $Y=0.42 $X2=0 $Y2=0
cc_368 N_A_44_47#_c_372_n N_VGND_c_846_n 0.00278633f $X=2.015 $Y=0.71 $X2=0
+ $Y2=0
cc_369 N_A_44_47#_c_378_n N_VGND_c_847_n 0.00257076f $X=3.465 $Y=0.71 $X2=0
+ $Y2=0
cc_370 N_A_44_47#_c_487_p N_VGND_c_847_n 0.012699f $X=3.56 $Y=0.445 $X2=0 $Y2=0
cc_371 N_A_44_47#_c_346_n N_VGND_c_847_n 0.0526223f $X=4.415 $Y=0.36 $X2=0 $Y2=0
cc_372 N_A_44_47#_c_338_n N_VGND_c_849_n 0.00486043f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_44_47#_c_339_n N_VGND_c_849_n 0.00353537f $X=6.475 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A_44_47#_c_340_n N_VGND_c_850_n 0.00353537f $X=6.905 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_A_44_47#_c_341_n N_VGND_c_850_n 0.00353537f $X=7.335 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_44_47#_c_342_n N_VGND_c_851_n 0.0170956f $X=0.345 $Y=0.42 $X2=0 $Y2=0
cc_377 N_A_44_47#_c_344_n N_VGND_c_851_n 0.00250404f $X=0.87 $Y=0.72 $X2=0 $Y2=0
cc_378 N_A_44_47#_c_372_n N_VGND_c_853_n 0.00262929f $X=2.015 $Y=0.71 $X2=0
+ $Y2=0
cc_379 N_A_44_47#_c_496_p N_VGND_c_853_n 0.0153733f $X=2.1 $Y=0.42 $X2=0 $Y2=0
cc_380 N_A_44_47#_c_378_n N_VGND_c_853_n 0.00271564f $X=3.465 $Y=0.71 $X2=0
+ $Y2=0
cc_381 N_A_44_47#_c_378_n N_VGND_c_854_n 0.0574448f $X=3.465 $Y=0.71 $X2=0 $Y2=0
cc_382 N_A_44_47#_M1000_s N_VGND_c_858_n 0.00229835f $X=0.22 $Y=0.235 $X2=0
+ $Y2=0
cc_383 N_A_44_47#_M1001_s N_VGND_c_858_n 0.00234465f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_384 N_A_44_47#_M1016_s N_VGND_c_858_n 0.00302097f $X=1.96 $Y=0.235 $X2=0
+ $Y2=0
cc_385 N_A_44_47#_M1019_d N_VGND_c_858_n 0.00243723f $X=3.415 $Y=0.235 $X2=0
+ $Y2=0
cc_386 N_A_44_47#_M1026_s N_VGND_c_858_n 0.00225742f $X=4.28 $Y=0.235 $X2=0
+ $Y2=0
cc_387 N_A_44_47#_c_338_n N_VGND_c_858_n 0.00822531f $X=6.045 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_A_44_47#_c_339_n N_VGND_c_858_n 0.00411309f $X=6.475 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_A_44_47#_c_340_n N_VGND_c_858_n 0.00411309f $X=6.905 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A_44_47#_c_341_n N_VGND_c_858_n 0.00411309f $X=7.335 $Y=0.995 $X2=0
+ $Y2=0
cc_391 N_A_44_47#_c_342_n N_VGND_c_858_n 0.00979174f $X=0.345 $Y=0.42 $X2=0
+ $Y2=0
cc_392 N_A_44_47#_c_365_n N_VGND_c_858_n 0.00417883f $X=1.11 $Y=0.72 $X2=0 $Y2=0
cc_393 N_A_44_47#_c_344_n N_VGND_c_858_n 0.00568091f $X=0.87 $Y=0.72 $X2=0 $Y2=0
cc_394 N_A_44_47#_c_484_p N_VGND_c_858_n 0.00873251f $X=1.205 $Y=0.42 $X2=0
+ $Y2=0
cc_395 N_A_44_47#_c_372_n N_VGND_c_858_n 0.0100254f $X=2.015 $Y=0.71 $X2=0 $Y2=0
cc_396 N_A_44_47#_c_496_p N_VGND_c_858_n 0.00853098f $X=2.1 $Y=0.42 $X2=0 $Y2=0
cc_397 N_A_44_47#_c_378_n N_VGND_c_858_n 0.0128404f $X=3.465 $Y=0.71 $X2=0 $Y2=0
cc_398 N_A_44_47#_c_487_p N_VGND_c_858_n 0.00731723f $X=3.56 $Y=0.445 $X2=0
+ $Y2=0
cc_399 N_A_44_47#_c_346_n N_VGND_c_858_n 0.0332109f $X=4.415 $Y=0.36 $X2=0 $Y2=0
cc_400 N_A_44_47#_c_346_n N_A_770_47#_M1010_d 0.00323484f $X=4.415 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_401 N_A_44_47#_M1026_s N_A_770_47#_c_974_n 0.0062344f $X=4.28 $Y=0.235 $X2=0
+ $Y2=0
cc_402 N_A_44_47#_c_346_n N_A_770_47#_c_974_n 0.0399725f $X=4.415 $Y=0.36 $X2=0
+ $Y2=0
cc_403 N_A_44_47#_c_355_n N_A_770_47#_c_974_n 0.00518284f $X=5.795 $Y=1.535
+ $X2=0 $Y2=0
cc_404 N_A_30_297#_c_524_n N_A_285_297#_M1006_d 0.0033237f $X=1.9 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_405 N_A_30_297#_c_524_n N_A_285_297#_c_562_n 0.0159794f $X=1.9 $Y=2.38 $X2=0
+ $Y2=0
cc_406 N_A_30_297#_M1024_s N_A_285_297#_c_559_n 0.00277342f $X=1.855 $Y=1.485
+ $X2=0 $Y2=0
cc_407 N_A_30_297#_c_524_n N_A_285_297#_c_559_n 0.00267072f $X=1.9 $Y=2.38 $X2=0
+ $Y2=0
cc_408 N_A_30_297#_c_525_n N_A_285_297#_c_559_n 0.0202075f $X=1.99 $Y=1.96 $X2=0
+ $Y2=0
cc_409 N_A_30_297#_c_523_n N_A_285_297#_c_560_n 0.00827545f $X=1.135 $Y=1.62
+ $X2=0 $Y2=0
cc_410 N_A_30_297#_c_525_n N_A_477_297#_c_595_n 0.0392482f $X=1.99 $Y=1.96 $X2=0
+ $Y2=0
cc_411 N_A_30_297#_c_524_n N_A_477_297#_c_596_n 0.0152916f $X=1.9 $Y=2.38 $X2=0
+ $Y2=0
cc_412 N_A_30_297#_c_529_n N_VPWR_c_666_n 0.0361203f $X=1.04 $Y=2.38 $X2=0 $Y2=0
cc_413 N_A_30_297#_c_522_n N_VPWR_c_666_n 0.0179012f $X=0.37 $Y=2.38 $X2=0 $Y2=0
cc_414 N_A_30_297#_c_524_n N_VPWR_c_666_n 0.0540284f $X=1.9 $Y=2.38 $X2=0 $Y2=0
cc_415 N_A_30_297#_c_551_p N_VPWR_c_666_n 0.0125248f $X=1.135 $Y=2.3 $X2=0 $Y2=0
cc_416 N_A_30_297#_M1005_s N_VPWR_c_658_n 0.00213422f $X=0.15 $Y=1.485 $X2=0
+ $Y2=0
cc_417 N_A_30_297#_M1018_s N_VPWR_c_658_n 0.00223239f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_418 N_A_30_297#_M1024_s N_VPWR_c_658_n 0.00209323f $X=1.855 $Y=1.485 $X2=0
+ $Y2=0
cc_419 N_A_30_297#_c_529_n N_VPWR_c_658_n 0.0234424f $X=1.04 $Y=2.38 $X2=0 $Y2=0
cc_420 N_A_30_297#_c_522_n N_VPWR_c_658_n 0.010004f $X=0.37 $Y=2.38 $X2=0 $Y2=0
cc_421 N_A_30_297#_c_524_n N_VPWR_c_658_n 0.0334515f $X=1.9 $Y=2.38 $X2=0 $Y2=0
cc_422 N_A_30_297#_c_551_p N_VPWR_c_658_n 0.00730678f $X=1.135 $Y=2.3 $X2=0
+ $Y2=0
cc_423 N_A_285_297#_c_559_n N_A_477_297#_M1004_d 0.00277342f $X=2.845 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_424 N_A_285_297#_c_559_n N_A_477_297#_c_595_n 0.0223717f $X=2.845 $Y=1.54
+ $X2=0 $Y2=0
cc_425 N_A_285_297#_M1004_s N_A_477_297#_c_602_n 0.0033237f $X=2.795 $Y=1.485
+ $X2=0 $Y2=0
cc_426 N_A_285_297#_c_559_n N_A_477_297#_c_602_n 0.00256303f $X=2.845 $Y=1.54
+ $X2=0 $Y2=0
cc_427 N_A_285_297#_c_561_n N_A_477_297#_c_602_n 0.0143067f $X=2.935 $Y=1.62
+ $X2=0 $Y2=0
cc_428 N_A_285_297#_c_561_n N_A_477_297#_c_605_n 0.0133012f $X=2.935 $Y=1.62
+ $X2=0 $Y2=0
cc_429 N_A_285_297#_c_561_n N_A_477_297#_c_607_n 0.00809064f $X=2.935 $Y=1.62
+ $X2=0 $Y2=0
cc_430 N_A_285_297#_M1006_d N_VPWR_c_658_n 0.00224864f $X=1.425 $Y=1.485 $X2=0
+ $Y2=0
cc_431 N_A_285_297#_M1004_s N_VPWR_c_658_n 0.00224864f $X=2.795 $Y=1.485 $X2=0
+ $Y2=0
cc_432 N_A_477_297#_c_610_n N_VPWR_M1002_d 0.00337663f $X=4.365 $Y=1.895
+ $X2=-0.19 $Y2=1.305
cc_433 N_A_477_297#_c_598_n N_VPWR_M1003_s 0.00547849f $X=5.31 $Y=1.895 $X2=0
+ $Y2=0
cc_434 N_A_477_297#_c_602_n N_VPWR_c_659_n 0.0117125f $X=3.32 $Y=2.38 $X2=0
+ $Y2=0
cc_435 N_A_477_297#_c_607_n N_VPWR_c_659_n 0.00839072f $X=3.485 $Y=2.24 $X2=0
+ $Y2=0
cc_436 N_A_477_297#_c_610_n N_VPWR_c_659_n 0.0166041f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_437 N_A_477_297#_c_610_n N_VPWR_c_660_n 0.00202688f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_438 N_A_477_297#_c_597_n N_VPWR_c_660_n 0.0134005f $X=4.455 $Y=2.25 $X2=0
+ $Y2=0
cc_439 N_A_477_297#_c_598_n N_VPWR_c_660_n 0.00276164f $X=5.31 $Y=1.895 $X2=0
+ $Y2=0
cc_440 N_A_477_297#_c_597_n N_VPWR_c_661_n 0.0125846f $X=4.455 $Y=2.25 $X2=0
+ $Y2=0
cc_441 N_A_477_297#_c_598_n N_VPWR_c_661_n 0.0149001f $X=5.31 $Y=1.895 $X2=0
+ $Y2=0
cc_442 N_A_477_297#_c_602_n N_VPWR_c_666_n 0.0586986f $X=3.32 $Y=2.38 $X2=0
+ $Y2=0
cc_443 N_A_477_297#_c_596_n N_VPWR_c_666_n 0.021548f $X=2.675 $Y=2.38 $X2=0
+ $Y2=0
cc_444 N_A_477_297#_c_610_n N_VPWR_c_666_n 0.00260213f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_445 N_A_477_297#_c_598_n N_VPWR_c_667_n 0.001998f $X=5.31 $Y=1.895 $X2=0
+ $Y2=0
cc_446 N_A_477_297#_c_623_n N_VPWR_c_667_n 0.0122637f $X=5.4 $Y=1.96 $X2=0 $Y2=0
cc_447 N_A_477_297#_M1004_d N_VPWR_c_658_n 0.00210122f $X=2.385 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_477_297#_M1014_d N_VPWR_c_658_n 0.00460897f $X=3.225 $Y=1.485 $X2=0
+ $Y2=0
cc_449 N_A_477_297#_M1017_s N_VPWR_c_658_n 0.00234332f $X=4.32 $Y=1.485 $X2=0
+ $Y2=0
cc_450 N_A_477_297#_M1003_d N_VPWR_c_658_n 0.00403008f $X=5.26 $Y=1.485 $X2=0
+ $Y2=0
cc_451 N_A_477_297#_c_602_n N_VPWR_c_658_n 0.035492f $X=3.32 $Y=2.38 $X2=0 $Y2=0
cc_452 N_A_477_297#_c_596_n N_VPWR_c_658_n 0.0127592f $X=2.675 $Y=2.38 $X2=0
+ $Y2=0
cc_453 N_A_477_297#_c_610_n N_VPWR_c_658_n 0.0102815f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_454 N_A_477_297#_c_597_n N_VPWR_c_658_n 0.00966008f $X=4.455 $Y=2.25 $X2=0
+ $Y2=0
cc_455 N_A_477_297#_c_598_n N_VPWR_c_658_n 0.0102699f $X=5.31 $Y=1.895 $X2=0
+ $Y2=0
cc_456 N_A_477_297#_c_623_n N_VPWR_c_658_n 0.0070449f $X=5.4 $Y=1.96 $X2=0 $Y2=0
cc_457 N_VPWR_c_658_n N_X_M1007_d 0.00535672f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_658_n N_X_M1025_d 0.00535672f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_668_n N_X_c_809_n 0.0124538f $X=6.525 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_658_n N_X_c_809_n 0.00724021f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_461 N_VPWR_M1013_s N_X_c_777_n 0.00178571f $X=6.55 $Y=1.485 $X2=0 $Y2=0
cc_462 N_VPWR_c_663_n N_X_c_777_n 0.0175375f $X=6.69 $Y=1.97 $X2=0 $Y2=0
cc_463 N_VPWR_c_669_n N_X_c_813_n 0.0124538f $X=7.385 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_658_n N_X_c_813_n 0.00724021f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_M1027_s N_X_c_779_n 2.33864e-19 $X=7.41 $Y=1.485 $X2=0 $Y2=0
cc_466 N_VPWR_c_665_n N_X_c_779_n 0.00362085f $X=7.55 $Y=1.97 $X2=0 $Y2=0
cc_467 N_VPWR_M1027_s N_X_c_781_n 0.00275297f $X=7.41 $Y=1.485 $X2=0 $Y2=0
cc_468 N_VPWR_c_665_n N_X_c_781_n 0.0203341f $X=7.55 $Y=1.97 $X2=0 $Y2=0
cc_469 N_X_c_783_n N_VGND_M1012_s 0.00365795f $X=7.025 $Y=0.72 $X2=0 $Y2=0
cc_470 N_X_c_797_n N_VGND_M1021_s 6.61764e-19 $X=7.49 $Y=0.72 $X2=0 $Y2=0
cc_471 N_X_c_775_n N_VGND_M1021_s 0.00276922f $X=7.612 $Y=0.805 $X2=0 $Y2=0
cc_472 X N_VGND_M1021_s 0.00128565f $X=7.61 $Y=0.85 $X2=0 $Y2=0
cc_473 N_X_c_783_n N_VGND_c_843_n 0.014476f $X=7.025 $Y=0.72 $X2=0 $Y2=0
cc_474 N_X_c_775_n N_VGND_c_844_n 4.07212e-19 $X=7.612 $Y=0.805 $X2=0 $Y2=0
cc_475 N_X_c_797_n N_VGND_c_845_n 0.00339507f $X=7.49 $Y=0.72 $X2=0 $Y2=0
cc_476 N_X_c_775_n N_VGND_c_845_n 0.0190055f $X=7.612 $Y=0.805 $X2=0 $Y2=0
cc_477 N_X_c_827_p N_VGND_c_849_n 0.0122747f $X=6.26 $Y=0.42 $X2=0 $Y2=0
cc_478 N_X_c_783_n N_VGND_c_849_n 0.00247598f $X=7.025 $Y=0.72 $X2=0 $Y2=0
cc_479 N_X_c_783_n N_VGND_c_850_n 0.00247598f $X=7.025 $Y=0.72 $X2=0 $Y2=0
cc_480 N_X_c_830_p N_VGND_c_850_n 0.0122747f $X=7.12 $Y=0.42 $X2=0 $Y2=0
cc_481 N_X_c_797_n N_VGND_c_850_n 0.00247598f $X=7.49 $Y=0.72 $X2=0 $Y2=0
cc_482 N_X_M1009_d N_VGND_c_858_n 0.00394701f $X=6.12 $Y=0.235 $X2=0 $Y2=0
cc_483 N_X_M1020_d N_VGND_c_858_n 0.00253729f $X=6.98 $Y=0.235 $X2=0 $Y2=0
cc_484 N_X_c_827_p N_VGND_c_858_n 0.00720049f $X=6.26 $Y=0.42 $X2=0 $Y2=0
cc_485 N_X_c_783_n N_VGND_c_858_n 0.00986428f $X=7.025 $Y=0.72 $X2=0 $Y2=0
cc_486 N_X_c_830_p N_VGND_c_858_n 0.00720049f $X=7.12 $Y=0.42 $X2=0 $Y2=0
cc_487 N_X_c_797_n N_VGND_c_858_n 0.0046298f $X=7.49 $Y=0.72 $X2=0 $Y2=0
cc_488 N_X_c_775_n N_VGND_c_858_n 0.00177799f $X=7.612 $Y=0.805 $X2=0 $Y2=0
cc_489 N_VGND_c_858_n N_A_770_47#_M1010_d 0.00224864f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_490 N_VGND_c_858_n N_A_770_47#_M1011_s 0.00395122f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_M1011_d N_A_770_47#_c_974_n 0.00594858f $X=4.83 $Y=0.235 $X2=0
+ $Y2=0
cc_492 N_VGND_c_841_n N_A_770_47#_c_974_n 0.0208104f $X=4.975 $Y=0.36 $X2=0
+ $Y2=0
cc_493 N_VGND_c_847_n N_A_770_47#_c_974_n 0.00418723f $X=4.805 $Y=0 $X2=0 $Y2=0
cc_494 N_VGND_c_848_n N_A_770_47#_c_974_n 0.00256355f $X=5.665 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_858_n N_A_770_47#_c_974_n 0.013632f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_848_n N_A_770_47#_c_993_n 0.0120665f $X=5.665 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_858_n N_A_770_47#_c_993_n 0.0070024f $X=7.59 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor4_2.pxi.spice
* Created: Tue Sep  1 19:19:01 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4_2%A N_A_c_72_n N_A_M1004_g N_A_M1001_g N_A_c_73_n
+ N_A_M1007_g N_A_M1015_g A N_A_c_75_n PM_SKY130_FD_SC_HD__NOR4_2%A
x_PM_SKY130_FD_SC_HD__NOR4_2%B N_B_c_112_n N_B_M1002_g N_B_M1010_g N_B_c_113_n
+ N_B_M1006_g N_B_M1012_g B N_B_c_115_n PM_SKY130_FD_SC_HD__NOR4_2%B
x_PM_SKY130_FD_SC_HD__NOR4_2%C N_C_c_156_n N_C_M1008_g N_C_M1000_g N_C_c_157_n
+ N_C_M1014_g N_C_M1003_g C N_C_c_158_n N_C_c_159_n PM_SKY130_FD_SC_HD__NOR4_2%C
x_PM_SKY130_FD_SC_HD__NOR4_2%D N_D_c_197_n N_D_M1009_g N_D_M1005_g N_D_c_198_n
+ N_D_M1011_g N_D_M1013_g D N_D_c_199_n N_D_c_200_n PM_SKY130_FD_SC_HD__NOR4_2%D
x_PM_SKY130_FD_SC_HD__NOR4_2%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1015_s
+ N_A_27_297#_M1012_d N_A_27_297#_c_240_n N_A_27_297#_c_259_p
+ N_A_27_297#_c_241_n N_A_27_297#_c_260_p N_A_27_297#_c_242_n
+ N_A_27_297#_c_243_n N_A_27_297#_c_244_n PM_SKY130_FD_SC_HD__NOR4_2%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR4_2%VPWR N_VPWR_M1001_d N_VPWR_c_277_n VPWR
+ N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_276_n N_VPWR_c_281_n
+ PM_SKY130_FD_SC_HD__NOR4_2%VPWR
x_PM_SKY130_FD_SC_HD__NOR4_2%A_281_297# N_A_281_297#_M1010_s
+ N_A_281_297#_M1000_s N_A_281_297#_c_327_n N_A_281_297#_c_323_n
+ N_A_281_297#_c_335_n N_A_281_297#_c_340_p
+ PM_SKY130_FD_SC_HD__NOR4_2%A_281_297#
x_PM_SKY130_FD_SC_HD__NOR4_2%A_475_297# N_A_475_297#_M1000_d
+ N_A_475_297#_M1003_d N_A_475_297#_M1013_d N_A_475_297#_c_342_n
+ N_A_475_297#_c_343_n N_A_475_297#_c_360_n N_A_475_297#_c_344_n
+ N_A_475_297#_c_374_p N_A_475_297#_c_345_n
+ PM_SKY130_FD_SC_HD__NOR4_2%A_475_297#
x_PM_SKY130_FD_SC_HD__NOR4_2%Y N_Y_M1004_s N_Y_M1002_d N_Y_M1008_d N_Y_M1009_s
+ N_Y_M1005_s N_Y_c_390_n N_Y_c_377_n N_Y_c_378_n N_Y_c_398_n N_Y_c_379_n
+ N_Y_c_412_n N_Y_c_380_n N_Y_c_415_n N_Y_c_387_n N_Y_c_381_n N_Y_c_382_n
+ N_Y_c_383_n N_Y_c_384_n N_Y_c_388_n Y N_Y_c_386_n PM_SKY130_FD_SC_HD__NOR4_2%Y
x_PM_SKY130_FD_SC_HD__NOR4_2%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_M1006_s
+ N_VGND_M1008_s N_VGND_M1014_s N_VGND_M1011_d N_VGND_c_486_n N_VGND_c_487_n
+ N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n
+ N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n VGND N_VGND_c_496_n
+ N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n PM_SKY130_FD_SC_HD__NOR4_2%VGND
cc_1 VNB N_A_c_72_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_73_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB A 0.0140266f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_4 VNB N_A_c_75_n 0.0382849f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_5 VNB N_B_c_112_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_113_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_7 VNB B 0.00791736f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_B_c_115_n 0.0369647f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_9 VNB N_C_c_156_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_C_c_157_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_11 VNB N_C_c_158_n 0.0167322f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_12 VNB N_C_c_159_n 0.0382791f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_13 VNB N_D_c_197_n 0.0160105f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_D_c_198_n 0.0191824f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_15 VNB N_D_c_199_n 0.00449738f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_16 VNB N_D_c_200_n 0.0332279f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_17 VNB N_VPWR_c_276_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_18 VNB N_Y_c_377_n 0.00338427f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_19 VNB N_Y_c_378_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_20 VNB N_Y_c_379_n 0.0158955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_380_n 0.00317397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_381_n 0.00152735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_382_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_383_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_384_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.02266f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_386_n 0.0109627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_486_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_29 VNB N_VGND_c_487_n 0.0351006f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_30 VNB N_VGND_c_488_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_489_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_490_n 0.0135581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_491_n 0.0181289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_492_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_493_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_494_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_495_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_496_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_497_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_498_n 0.0264442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_499_n 0.237811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_A_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_43 VPB N_A_M1015_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_44 VPB N_A_c_75_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_45 VPB N_B_M1010_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_46 VPB N_B_M1012_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_47 VPB N_B_c_115_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_48 VPB N_C_M1000_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_49 VPB N_C_M1003_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_50 VPB N_C_c_159_n 0.00480973f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_51 VPB N_D_M1005_g 0.0188145f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_52 VPB N_D_M1013_g 0.0219473f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_53 VPB N_D_c_200_n 0.00422661f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_54 VPB N_A_27_297#_c_240_n 0.00402354f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_55 VPB N_A_27_297#_c_241_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_297#_c_242_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_57 VPB N_A_27_297#_c_243_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_297#_c_244_n 0.003591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_277_n 0.00516508f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_60 VPB N_VPWR_c_278_n 0.0180608f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_61 VPB N_VPWR_c_279_n 0.0936174f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_62 VPB N_VPWR_c_276_n 0.0553414f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_63 VPB N_VPWR_c_281_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_281_297#_c_323_n 0.0128761f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.325
cc_65 VPB N_A_475_297#_c_342_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_66 VPB N_A_475_297#_c_343_n 0.00323111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_475_297#_c_344_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_475_297#_c_345_n 0.00268836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_387_n 0.0175146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_388_n 0.00225182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB Y 0.00855033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 N_A_c_73_n N_B_c_112_n 0.0194931f $X=0.91 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_73 N_A_M1015_g N_B_M1010_g 0.0194931f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_74 A B 0.0185436f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_75_n B 0.00160637f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_76 A N_B_c_115_n 2.03927e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_B_c_115_n 0.0194931f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_78 A N_A_27_297#_c_240_n 0.0175673f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_A_27_297#_c_241_n 0.0134951f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_80 N_A_M1015_g N_A_27_297#_c_241_n 0.0134675f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_81 A N_A_27_297#_c_241_n 0.0396361f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_75_n N_A_27_297#_c_241_n 0.00211509f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1001_g N_VPWR_c_277_n 0.00302074f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_M1015_g N_VPWR_c_277_n 0.00302074f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_VPWR_c_278_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1015_g N_VPWR_c_279_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VPWR_c_276_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_88 N_A_M1015_g N_VPWR_c_276_n 0.010464f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_89 N_A_c_72_n N_Y_c_390_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_c_73_n N_Y_c_390_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_73_n N_Y_c_377_n 0.00890517f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_92 A N_Y_c_377_n 0.00688575f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_c_72_n N_Y_c_378_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_c_73_n N_Y_c_378_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_95 A N_Y_c_378_n 0.0266272f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_75_n N_Y_c_378_n 0.00230339f $X=0.91 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_c_73_n N_Y_c_398_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_c_72_n N_VGND_c_487_n 0.00366968f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_99 A N_VGND_c_487_n 0.0140538f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_c_73_n N_VGND_c_488_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_72_n N_VGND_c_492_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_c_73_n N_VGND_c_492_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_c_72_n N_VGND_c_499_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_73_n N_VGND_c_499_n 0.0057435f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_105 B N_C_c_158_n 0.0140819f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_106 N_B_c_115_n N_C_c_158_n 0.00122605f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B_M1010_g N_A_27_297#_c_242_n 0.0132199f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B_M1012_g N_A_27_297#_c_242_n 0.0112055f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_109 B N_A_27_297#_c_242_n 0.0417417f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_110 N_B_c_115_n N_A_27_297#_c_242_n 0.00211509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_111 B N_A_27_297#_c_243_n 0.00942636f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_112 B N_A_27_297#_c_244_n 0.0089871f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_113 N_B_M1010_g N_VPWR_c_279_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B_M1012_g N_VPWR_c_279_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B_M1010_g N_VPWR_c_276_n 0.0106871f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B_M1012_g N_VPWR_c_276_n 0.00660224f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B_M1012_g N_A_281_297#_c_323_n 0.0119904f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_118 N_B_M1012_g N_A_475_297#_c_345_n 4.91095e-19 $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B_c_112_n N_Y_c_390_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B_c_112_n N_Y_c_377_n 0.00865686f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_121 B N_Y_c_377_n 0.0174927f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B_c_112_n N_Y_c_398_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_113_n N_Y_c_398_n 0.0109565f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_113_n N_Y_c_379_n 0.0109318f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_125 B N_Y_c_379_n 0.0171084f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_c_112_n N_Y_c_382_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_113_n N_Y_c_382_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_128 B N_Y_c_382_n 0.0266272f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B_c_115_n N_Y_c_382_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_c_112_n N_VGND_c_488_n 0.00146339f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B_c_112_n N_VGND_c_497_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_c_113_n N_VGND_c_497_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_113_n N_VGND_c_498_n 0.00336547f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B_c_112_n N_VGND_c_499_n 0.0057435f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B_c_113_n N_VGND_c_499_n 0.0070399f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_136 N_C_c_157_n N_D_c_197_n 0.0194216f $X=3.15 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_137 N_C_M1003_g N_D_M1005_g 0.0194216f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_138 N_C_c_158_n N_D_c_199_n 0.01435f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_139 N_C_c_159_n N_D_c_199_n 0.00192374f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_140 N_C_c_159_n N_D_c_200_n 0.0194216f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C_M1000_g N_A_27_297#_c_244_n 4.91095e-19 $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_C_M1000_g N_VPWR_c_279_n 0.00357877f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_143 N_C_M1003_g N_VPWR_c_279_n 0.00585385f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_144 N_C_M1000_g N_VPWR_c_276_n 0.00660224f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_145 N_C_M1003_g N_VPWR_c_276_n 0.0106871f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_146 N_C_M1000_g N_A_281_297#_c_323_n 0.0119904f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_147 N_C_M1000_g N_A_475_297#_c_342_n 0.0111613f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_148 N_C_M1003_g N_A_475_297#_c_342_n 0.0146546f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_149 N_C_c_158_n N_A_475_297#_c_342_n 0.0327461f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_150 N_C_c_159_n N_A_475_297#_c_342_n 0.00211509f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_151 N_C_c_158_n N_A_475_297#_c_345_n 0.0213978f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_152 N_C_c_156_n N_Y_c_379_n 0.0109318f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_153 N_C_c_158_n N_Y_c_379_n 0.0424717f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_154 N_C_c_156_n N_Y_c_412_n 0.0109565f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C_c_157_n N_Y_c_412_n 0.00630972f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C_c_157_n N_Y_c_380_n 0.0101343f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_157 N_C_c_157_n N_Y_c_415_n 5.22228e-19 $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_158 N_C_c_156_n N_Y_c_383_n 0.00113286f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_159 N_C_c_157_n N_Y_c_383_n 0.00113286f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_160 N_C_c_158_n N_Y_c_383_n 0.0266272f $X=2.94 $Y=1.16 $X2=0 $Y2=0
cc_161 N_C_c_159_n N_Y_c_383_n 0.00230339f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_162 N_C_c_157_n N_VGND_c_489_n 0.00146339f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_163 N_C_c_156_n N_VGND_c_494_n 0.00423334f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C_c_157_n N_VGND_c_494_n 0.00423334f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C_c_156_n N_VGND_c_498_n 0.00336547f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_166 N_C_c_156_n N_VGND_c_499_n 0.0070399f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_167 N_C_c_157_n N_VGND_c_499_n 0.0057435f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_168 N_D_M1005_g N_VPWR_c_279_n 0.00357877f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_169 N_D_M1013_g N_VPWR_c_279_n 0.00357877f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_170 N_D_M1005_g N_VPWR_c_276_n 0.00525237f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_171 N_D_M1013_g N_VPWR_c_276_n 0.00628918f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_172 N_D_M1005_g N_A_475_297#_c_343_n 2.57315e-19 $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_173 N_D_c_199_n N_A_475_297#_c_343_n 0.0124257f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_174 N_D_M1005_g N_A_475_297#_c_344_n 0.0121306f $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_175 N_D_M1013_g N_A_475_297#_c_344_n 0.00984328f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_176 N_D_c_197_n N_Y_c_412_n 5.22228e-19 $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_177 N_D_c_197_n N_Y_c_380_n 0.00865686f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_178 N_D_c_199_n N_Y_c_380_n 0.0201828f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_179 N_D_c_197_n N_Y_c_415_n 0.00630972f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_180 N_D_c_198_n N_Y_c_415_n 0.0109314f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_181 N_D_M1013_g N_Y_c_387_n 0.0143208f $X=3.99 $Y=1.985 $X2=0 $Y2=0
cc_182 N_D_c_199_n N_Y_c_387_n 0.00137795f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_183 N_D_c_198_n N_Y_c_381_n 0.0119544f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_184 N_D_c_197_n N_Y_c_384_n 0.00113286f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_185 N_D_c_198_n N_Y_c_384_n 0.00133956f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_186 N_D_c_199_n N_Y_c_384_n 0.0250867f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_187 N_D_c_200_n N_Y_c_384_n 0.00230339f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_188 N_D_M1005_g N_Y_c_388_n 2.57315e-19 $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_189 N_D_c_199_n N_Y_c_388_n 0.0204292f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_190 N_D_c_200_n N_Y_c_388_n 0.00219557f $X=3.99 $Y=1.16 $X2=0 $Y2=0
cc_191 N_D_c_198_n Y 0.0201093f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_192 N_D_c_199_n Y 0.0127368f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_193 N_D_c_197_n N_VGND_c_489_n 0.00146448f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_194 N_D_c_198_n N_VGND_c_491_n 0.0032322f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_195 N_D_c_197_n N_VGND_c_496_n 0.00423334f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_196 N_D_c_198_n N_VGND_c_496_n 0.00423334f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_197 N_D_c_197_n N_VGND_c_499_n 0.0057435f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_198 N_D_c_198_n N_VGND_c_499_n 0.00678032f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_27_297#_c_241_n N_VPWR_M1001_d 0.00165831f $X=0.995 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_200 N_A_27_297#_c_241_n N_VPWR_c_277_n 0.0126919f $X=0.995 $Y=1.54 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_259_p N_VPWR_c_278_n 0.0161885f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_202 N_A_27_297#_c_260_p N_VPWR_c_279_n 0.0142343f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_203 N_A_27_297#_M1001_s N_VPWR_c_276_n 0.00315976f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_M1015_s N_VPWR_c_276_n 0.00284632f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_M1012_d N_VPWR_c_276_n 0.00226545f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_259_p N_VPWR_c_276_n 0.00974347f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_207 N_A_27_297#_c_260_p N_VPWR_c_276_n 0.00955092f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_208 N_A_27_297#_c_242_n N_A_281_297#_M1010_s 0.00165831f $X=1.835 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_209 N_A_27_297#_c_242_n N_A_281_297#_c_327_n 0.0126766f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_210 N_A_27_297#_M1012_d N_A_281_297#_c_323_n 0.00593473f $X=1.825 $Y=1.485
+ $X2=0 $Y2=0
cc_211 N_A_27_297#_c_242_n N_A_281_297#_c_323_n 0.00320918f $X=1.835 $Y=1.54
+ $X2=0 $Y2=0
cc_212 N_A_27_297#_c_244_n N_A_281_297#_c_323_n 0.0153739f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_244_n N_A_475_297#_c_345_n 0.0346205f $X=1.96 $Y=1.62 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_241_n N_Y_c_377_n 8.37688e-19 $X=0.995 $Y=1.54 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_243_n N_Y_c_377_n 0.00524452f $X=1.12 $Y=1.62 $X2=0 $Y2=0
cc_216 N_A_27_297#_c_244_n N_Y_c_379_n 0.00542522f $X=1.96 $Y=1.62 $X2=0 $Y2=0
cc_217 N_A_27_297#_c_240_n N_VGND_c_487_n 0.00206382f $X=0.277 $Y=1.625 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_276_n N_A_281_297#_M1010_s 0.00246446f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_219 N_VPWR_c_276_n N_A_281_297#_M1000_s 0.00246446f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_279_n N_A_281_297#_c_323_n 0.0830896f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_276_n N_A_281_297#_c_323_n 0.0509444f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_279_n N_A_281_297#_c_335_n 0.0142933f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_276_n N_A_281_297#_c_335_n 0.00962421f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_276_n N_A_475_297#_M1000_d 0.00226545f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_225 N_VPWR_c_276_n N_A_475_297#_M1003_d 0.00246446f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_276_n N_A_475_297#_M1013_d 0.0020932f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_279_n N_A_475_297#_c_360_n 0.0143053f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_276_n N_A_475_297#_c_360_n 0.00962794f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_279_n N_A_475_297#_c_344_n 0.0489446f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_276_n N_A_475_297#_c_344_n 0.0300869f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_276_n N_Y_M1005_s 0.00216833f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_232 N_A_281_297#_c_323_n N_A_475_297#_M1000_d 0.00593473f $X=2.815 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_233 N_A_281_297#_M1000_s N_A_475_297#_c_342_n 0.00165831f $X=2.805 $Y=1.485
+ $X2=0 $Y2=0
cc_234 N_A_281_297#_c_323_n N_A_475_297#_c_342_n 0.00320918f $X=2.815 $Y=2.38
+ $X2=0 $Y2=0
cc_235 N_A_281_297#_c_340_p N_A_475_297#_c_342_n 0.0126766f $X=2.94 $Y=1.96
+ $X2=0 $Y2=0
cc_236 N_A_281_297#_c_323_n N_A_475_297#_c_345_n 0.0153739f $X=2.815 $Y=2.38
+ $X2=0 $Y2=0
cc_237 N_A_475_297#_c_344_n N_Y_M1005_s 0.00312348f $X=4.075 $Y=2.38 $X2=0 $Y2=0
cc_238 N_A_475_297#_c_342_n N_Y_c_380_n 0.00342102f $X=3.235 $Y=1.54 $X2=0 $Y2=0
cc_239 N_A_475_297#_c_343_n N_Y_c_380_n 0.00393339f $X=3.36 $Y=1.625 $X2=0 $Y2=0
cc_240 N_A_475_297#_M1013_d N_Y_c_387_n 0.00281938f $X=4.065 $Y=1.485 $X2=0
+ $Y2=0
cc_241 N_A_475_297#_c_344_n N_Y_c_387_n 0.00320918f $X=4.075 $Y=2.38 $X2=0 $Y2=0
cc_242 N_A_475_297#_c_374_p N_Y_c_387_n 0.0176457f $X=4.2 $Y=1.96 $X2=0 $Y2=0
cc_243 N_A_475_297#_c_343_n N_Y_c_388_n 0.00271526f $X=3.36 $Y=1.625 $X2=0 $Y2=0
cc_244 N_A_475_297#_c_344_n N_Y_c_388_n 0.0118729f $X=4.075 $Y=2.38 $X2=0 $Y2=0
cc_245 N_Y_c_377_n N_VGND_M1007_d 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_246 N_Y_c_379_n N_VGND_M1006_s 0.00320259f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_247 N_Y_c_379_n N_VGND_M1008_s 0.00320259f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_248 N_Y_c_380_n N_VGND_M1014_s 0.00162089f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_249 N_Y_c_381_n N_VGND_M1011_d 5.9225e-19 $X=4.18 $Y=0.815 $X2=0 $Y2=0
cc_250 N_Y_c_386_n N_VGND_M1011_d 0.00227404f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_251 N_Y_c_378_n N_VGND_c_487_n 0.00835456f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_252 N_Y_c_377_n N_VGND_c_488_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_253 N_Y_c_380_n N_VGND_c_489_n 0.0122559f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_254 N_Y_c_386_n N_VGND_c_490_n 0.00187739f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_255 N_Y_c_381_n N_VGND_c_491_n 0.00452261f $X=4.18 $Y=0.815 $X2=0 $Y2=0
cc_256 N_Y_c_386_n N_VGND_c_491_n 0.0196389f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_257 N_Y_c_390_n N_VGND_c_492_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_258 N_Y_c_377_n N_VGND_c_492_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_259 N_Y_c_379_n N_VGND_c_494_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_260 N_Y_c_412_n N_VGND_c_494_n 0.0188551f $X=2.94 $Y=0.39 $X2=0 $Y2=0
cc_261 N_Y_c_380_n N_VGND_c_494_n 0.00198695f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_262 N_Y_c_380_n N_VGND_c_496_n 0.00198695f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_263 N_Y_c_415_n N_VGND_c_496_n 0.0188551f $X=3.78 $Y=0.39 $X2=0 $Y2=0
cc_264 N_Y_c_381_n N_VGND_c_496_n 0.00198695f $X=4.18 $Y=0.815 $X2=0 $Y2=0
cc_265 N_Y_c_377_n N_VGND_c_497_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_266 N_Y_c_398_n N_VGND_c_497_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_267 N_Y_c_379_n N_VGND_c_497_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_268 N_Y_c_379_n N_VGND_c_498_n 0.0567707f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_269 N_Y_M1004_s N_VGND_c_499_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_270 N_Y_M1002_d N_VGND_c_499_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_271 N_Y_M1008_d N_VGND_c_499_n 0.00215201f $X=2.805 $Y=0.235 $X2=0 $Y2=0
cc_272 N_Y_M1009_s N_VGND_c_499_n 0.00215201f $X=3.645 $Y=0.235 $X2=0 $Y2=0
cc_273 N_Y_c_390_n N_VGND_c_499_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_274 N_Y_c_377_n N_VGND_c_499_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_275 N_Y_c_398_n N_VGND_c_499_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_276 N_Y_c_379_n N_VGND_c_499_n 0.0104789f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_277 N_Y_c_412_n N_VGND_c_499_n 0.0122069f $X=2.94 $Y=0.39 $X2=0 $Y2=0
cc_278 N_Y_c_380_n N_VGND_c_499_n 0.00835832f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_279 N_Y_c_415_n N_VGND_c_499_n 0.0122069f $X=3.78 $Y=0.39 $X2=0 $Y2=0
cc_280 N_Y_c_381_n N_VGND_c_499_n 0.00410102f $X=4.18 $Y=0.815 $X2=0 $Y2=0
cc_281 N_Y_c_386_n N_VGND_c_499_n 0.00410715f $X=4.347 $Y=0.905 $X2=0 $Y2=0

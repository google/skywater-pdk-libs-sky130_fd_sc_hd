* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.08e+12p pd=1.016e+07u as=2.97e+12p ps=2.394e+07u
M1001 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=1.08e+12p pd=1.016e+07u as=0p ps=0u
M1002 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_297# B2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_803_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=8.645e+11p ps=9.16e+06u
M1009 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y A1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=0p ps=0u
M1011 a_803_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=9.16e+06u as=0p ps=0u
M1014 Y A1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_803_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_803_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A2 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y B2 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_803_47# A1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y B1 a_27_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_27_297# B2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_27_297# B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

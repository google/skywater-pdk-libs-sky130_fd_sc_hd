* File: sky130_fd_sc_hd__mux4_2.pex.spice
* Created: Tue Sep  1 19:15:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX4_2%S0 3 7 9 11 13 17 21 23 24 27 29 30 33 34 35
+ 36 43 45 46 52 58
c204 46 0 7.62213e-20 $X=6.21 $Y=1.53
c205 43 0 9.63205e-21 $X=1.15 $Y=1.53
c206 35 0 7.52734e-20 $X=6.065 $Y=1.53
c207 33 0 9.17818e-20 $X=1.005 $Y=1.53
c208 17 0 1.33206e-19 $X=1.91 $Y=0.415
r209 61 63 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.41
+ $X2=6.38 $Y2=1.575
r210 58 61 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.38 $Y=1.32 $X2=6.38
+ $Y2=1.41
r211 54 56 24.3813 $w=2.57e-07 $l=1.3e-07 $layer=POLY_cond $X=1.305 $Y=1.32
+ $X2=1.305 $Y2=1.45
r212 49 52 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r213 46 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.38
+ $Y=1.41 $X2=6.38 $Y2=1.41
r214 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.53
+ $X2=6.21 $Y2=1.53
r215 43 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.305
+ $Y=1.45 $X2=1.305 $Y2=1.45
r216 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.53
+ $X2=1.15 $Y2=1.53
r217 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.53
+ $X2=1.15 $Y2=1.53
r218 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.065 $Y=1.53
+ $X2=6.21 $Y2=1.53
r219 35 36 5.90345 $w=1.4e-07 $l=4.77e-06 $layer=MET1_cond $X=6.065 $Y=1.53
+ $X2=1.295 $Y2=1.53
r220 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.375 $Y=1.53
+ $X2=0.23 $Y2=1.53
r221 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.005 $Y=1.53
+ $X2=1.15 $Y2=1.53
r222 33 34 0.779701 $w=1.4e-07 $l=6.3e-07 $layer=MET1_cond $X=1.005 $Y=1.53
+ $X2=0.375 $Y2=1.53
r223 30 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=1.53
+ $X2=0.23 $Y2=1.53
r224 29 30 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.235 $Y2=1.53
r225 29 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r226 27 63 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.32 $Y=2.275
+ $X2=6.32 $Y2=1.575
r227 23 58 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.245 $Y=1.32
+ $X2=6.38 $Y2=1.32
r228 23 24 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.245 $Y=1.32
+ $X2=5.855 $Y2=1.32
r229 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.78 $Y=1.245
+ $X2=5.855 $Y2=1.32
r230 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.78 $Y=1.245
+ $X2=5.78 $Y2=0.415
r231 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.91 $Y=1.245
+ $X2=1.91 $Y2=0.415
r232 14 54 15.359 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.44 $Y=1.32
+ $X2=1.305 $Y2=1.32
r233 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.835 $Y=1.32
+ $X2=1.91 $Y2=1.245
r234 13 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.835 $Y=1.32
+ $X2=1.44 $Y2=1.32
r235 9 56 39.2307 $w=2.57e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.365 $Y=1.615
+ $X2=1.305 $Y2=1.45
r236 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=1.615
+ $X2=1.365 $Y2=2.275
r237 5 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r238 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=2.165
r239 1 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r240 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A2 5 8 10 11 12 13 18 20
c64 13 0 1.60286e-19 $X=1.15 $Y=0.85
c65 11 0 9.17818e-20 $X=0.887 $Y=1.715
r66 19 29 7.22896 $w=3.28e-07 $l=2.07e-07 $layer=LI1_cond $X=0.92 $Y=0.93
+ $X2=1.127 $Y2=0.93
r67 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=0.93
+ $X2=0.92 $Y2=1.095
r68 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=0.93
+ $X2=0.92 $Y2=0.765
r69 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.92
+ $Y=0.93 $X2=0.92 $Y2=0.93
r70 13 29 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=1.15 $Y=0.93
+ $X2=1.127 $Y2=0.93
r71 13 29 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.127 $Y=0.765
+ $X2=1.127 $Y2=0.93
r72 12 13 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.127 $Y=0.51
+ $X2=1.127 $Y2=0.765
r73 10 11 19.1365 $w=1.55e-07 $l=4e-08 $layer=POLY_cond $X=0.887 $Y=1.675
+ $X2=0.887 $Y2=1.715
r74 10 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.885 $Y=1.675
+ $X2=0.885 $Y2=1.095
r75 8 11 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.89 $Y=2.165
+ $X2=0.89 $Y2=1.715
r76 5 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A_27_47# 1 2 7 9 12 16 18 20 23 27 30 31 32
+ 37 43 45 51 54 55 61 69 70 74 75 80 85
c242 69 0 9.63205e-21 $X=1.815 $Y=1.74
c243 51 0 3.21039e-20 $X=6.2 $Y=0.87
r244 74 77 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.87 $Y=1.74
+ $X2=5.87 $Y2=1.875
r245 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.74 $X2=5.87 $Y2=1.74
r246 70 85 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=1.74
+ $X2=1.73 $Y2=1.575
r247 69 72 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.815 $Y=1.74
+ $X2=1.815 $Y2=1.875
r248 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.74 $X2=1.815 $Y2=1.74
r249 61 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.87
+ $X2=5.75 $Y2=1.87
r250 58 70 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.73 $Y=1.87
+ $X2=1.73 $Y2=1.74
r251 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.87
+ $X2=1.61 $Y2=1.87
r252 55 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.87
+ $X2=1.61 $Y2=1.87
r253 54 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.605 $Y=1.87
+ $X2=5.75 $Y2=1.87
r254 54 55 4.76484 $w=1.4e-07 $l=3.85e-06 $layer=MET1_cond $X=5.605 $Y=1.87
+ $X2=1.755 $Y2=1.87
r255 52 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=6.2 $Y=0.87 $X2=6.33
+ $Y2=0.87
r256 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.2
+ $Y=0.87 $X2=6.2 $Y2=0.87
r257 48 75 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.81 $Y=1.035
+ $X2=5.81 $Y2=1.74
r258 47 51 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.81 $Y=0.87
+ $X2=6.2 $Y2=0.87
r259 47 48 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=0.87
+ $X2=5.81 $Y2=1.035
r260 43 64 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.49 $Y=0.87
+ $X2=1.365 $Y2=0.87
r261 42 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.49 $Y=0.87
+ $X2=1.645 $Y2=0.87
r262 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=0.87 $X2=1.49 $Y2=0.87
r263 39 40 18.1581 $w=2.15e-07 $l=3.2e-07 $layer=LI1_cond $X=0.26 $Y=1.935
+ $X2=0.58 $Y2=1.935
r264 35 37 21.0727 $w=1.68e-07 $l=3.23e-07 $layer=LI1_cond $X=0.257 $Y=0.72
+ $X2=0.58 $Y2=0.72
r265 33 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=1.035
+ $X2=1.645 $Y2=0.87
r266 33 85 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.645 $Y=1.035
+ $X2=1.645 $Y2=1.575
r267 32 40 5.39194 $w=2.15e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.665 $Y=1.87
+ $X2=0.58 $Y2=1.935
r268 31 58 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.56 $Y=1.87
+ $X2=1.73 $Y2=1.87
r269 31 32 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.56 $Y=1.87
+ $X2=0.665 $Y2=1.87
r270 30 40 2.11506 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.58 $Y=1.785
+ $X2=0.58 $Y2=1.935
r271 29 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.58 $Y=0.805
+ $X2=0.58 $Y2=0.72
r272 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.58 $Y=0.805
+ $X2=0.58 $Y2=1.785
r273 25 39 2.11506 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=1.935
r274 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=2.085
+ $X2=0.26 $Y2=2.21
r275 21 35 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.72
r276 21 23 7.92208 $w=1.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.257 $Y=0.635
+ $X2=0.257 $Y2=0.51
r277 18 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.33 $Y=0.705
+ $X2=6.33 $Y2=0.87
r278 18 20 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.33 $Y=0.705
+ $X2=6.33 $Y2=0.415
r279 16 77 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.9 $Y=2.275 $X2=5.9
+ $Y2=1.875
r280 12 72 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.785 $Y=2.275
+ $X2=1.785 $Y2=1.875
r281 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.705
+ $X2=1.365 $Y2=0.87
r282 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.365 $Y=0.705
+ $X2=1.365 $Y2=0.415
r283 2 27 600 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.21
r284 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A3 3 5 6 8 11 13 14 18 20
c59 20 0 1.3041e-19 $X=2.405 $Y=0.765
c60 18 0 1.47056e-19 $X=2.405 $Y=0.93
c61 13 0 4.84598e-20 $X=2.53 $Y=0.85
r62 19 30 4.96365 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=2.427 $Y=0.93
+ $X2=2.427 $Y2=1.015
r63 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=0.93
+ $X2=2.405 $Y2=1.095
r64 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=0.93
+ $X2=2.405 $Y2=0.765
r65 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=0.93 $X2=2.405 $Y2=0.93
r66 14 30 9.46785 $w=2.03e-07 $l=1.75e-07 $layer=LI1_cond $X=2.512 $Y=1.19
+ $X2=2.512 $Y2=1.015
r67 13 19 2.45854 $w=3.73e-07 $l=8e-08 $layer=LI1_cond $X=2.427 $Y=0.85
+ $X2=2.427 $Y2=0.93
r68 9 11 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=2.39 $Y=1.575
+ $X2=2.505 $Y2=1.575
r69 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.65
+ $X2=2.505 $Y2=1.575
r70 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.505 $Y=1.65
+ $X2=2.505 $Y2=2.045
r71 5 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.39 $Y=1.5 $X2=2.39
+ $Y2=1.575
r72 5 21 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.39 $Y=1.5 $X2=2.39
+ $Y2=1.095
r73 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.39 $Y=0.445
+ $X2=2.39 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%S1 1 4 5 7 8 9 10 12 14 17 19 20
c86 19 0 1.3041e-19 $X=2.99 $Y=0.85
c87 5 0 4.84598e-20 $X=2.93 $Y=0.73
c88 1 0 3.58022e-19 $X=2.925 $Y=1.095
r89 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.885
+ $Y=0.93 $X2=2.885 $Y2=0.93
r90 23 25 23.1731 $w=2.6e-07 $l=1.25e-07 $layer=POLY_cond $X=2.885 $Y=0.805
+ $X2=2.885 $Y2=0.93
r91 20 26 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=2.93 $Y=1.19
+ $X2=2.93 $Y2=0.93
r92 19 26 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=2.93 $Y=0.85 $X2=2.93
+ $Y2=0.93
r93 15 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.285 $Y=2.465
+ $X2=4.285 $Y2=1.85
r94 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.445
r95 11 23 15.628 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.02 $Y=0.805
+ $X2=2.885 $Y2=0.805
r96 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.805 $Y=0.805
+ $X2=3.88 $Y2=0.73
r97 10 11 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.805 $Y=0.805
+ $X2=3.02 $Y2=0.805
r98 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.21 $Y=2.54
+ $X2=4.285 $Y2=2.465
r99 8 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=4.21 $Y=2.54 $X2=3
+ $Y2=2.54
r100 5 23 22.4589 $w=2.6e-07 $l=9.48683e-08 $layer=POLY_cond $X=2.93 $Y=0.73
+ $X2=2.885 $Y2=0.805
r101 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.93 $Y=0.73 $X2=2.93
+ $Y2=0.445
r102 2 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.925 $Y=2.465
+ $X2=3 $Y2=2.54
r103 2 4 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.925 $Y=2.465
+ $X2=2.925 $Y2=2.045
r104 1 25 39.1435 $w=2.6e-07 $l=1.83916e-07 $layer=POLY_cond $X=2.925 $Y=1.095
+ $X2=2.885 $Y2=0.93
r105 1 4 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.925 $Y=1.095
+ $X2=2.925 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A_600_345# 1 2 9 11 15 17 18 20 22 29
c69 22 0 2.63684e-19 $X=3.395 $Y=1.225
r70 27 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.15 $Y=0.38
+ $X2=3.33 $Y2=0.38
r71 22 25 31.9878 $w=2.46e-07 $l=7.25034e-07 $layer=LI1_cond $X=3.395 $Y=1.225
+ $X2=3.225 $Y2=1.87
r72 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.395
+ $Y=1.225 $X2=3.395 $Y2=1.225
r73 20 22 9.35836 $w=2.46e-07 $l=1.94808e-07 $layer=LI1_cond $X=3.33 $Y=1.06
+ $X2=3.395 $Y2=1.225
r74 19 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.465
+ $X2=3.33 $Y2=0.38
r75 19 20 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.33 $Y=0.465
+ $X2=3.33 $Y2=1.06
r76 17 23 87.7586 $w=2.7e-07 $l=3.95e-07 $layer=POLY_cond $X=3.79 $Y=1.225
+ $X2=3.395 $Y2=1.225
r77 17 18 15.2969 $w=2.1e-07 $l=7.5e-08 $layer=POLY_cond $X=3.79 $Y=1.225
+ $X2=3.865 $Y2=1.225
r78 13 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.305 $Y=1.09
+ $X2=4.305 $Y2=0.445
r79 12 18 15.2969 $w=2.1e-07 $l=1.00623e-07 $layer=POLY_cond $X=3.94 $Y=1.165
+ $X2=3.865 $Y2=1.225
r80 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.23 $Y=1.165
+ $X2=4.305 $Y2=1.09
r81 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.23 $Y=1.165
+ $X2=3.94 $Y2=1.165
r82 7 18 10.1846 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.865 $Y=1.36
+ $X2=3.865 $Y2=1.225
r83 7 9 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.865 $Y=1.36
+ $X2=3.865 $Y2=1.85
r84 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3
+ $Y=1.725 $X2=3.135 $Y2=1.87
r85 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.15 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A1 3 7 9 10 18
r40 17 18 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.225 $Y=1.23
+ $X2=5.245 $Y2=1.23
r41 14 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.03 $Y=1.23
+ $X2=5.225 $Y2=1.23
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.03
+ $Y=1.23 $X2=5.03 $Y2=1.23
r43 10 15 1.24588 $w=3.68e-07 $l=4e-08 $layer=LI1_cond $X=4.93 $Y=1.19 $X2=4.93
+ $Y2=1.23
r44 9 10 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.93 $Y=0.85 $X2=4.93
+ $Y2=1.19
r45 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.245 $Y=1.065
+ $X2=5.245 $Y2=1.23
r46 5 7 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.245 $Y=1.065
+ $X2=5.245 $Y2=0.445
r47 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.225 $Y=1.395
+ $X2=5.225 $Y2=1.23
r48 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.225 $Y=1.395
+ $X2=5.225 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A0 3 7 9 12 13 14
c49 12 0 3.6404e-19 $X=6.86 $Y=1.16
c50 9 0 4.70922e-20 $X=6.69 $Y=0.995
r51 13 14 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=6.69 $Y=0.51
+ $X2=6.69 $Y2=0.85
r52 12 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.86 $Y=1.16
+ $X2=6.86 $Y2=1.325
r53 12 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.86 $Y=1.16
+ $X2=6.86 $Y2=0.995
r54 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.16 $X2=6.86 $Y2=1.16
r55 9 14 5.39046 $w=3.08e-07 $l=1.45e-07 $layer=LI1_cond $X=6.69 $Y=0.995
+ $X2=6.69 $Y2=0.85
r56 9 11 6.10881 $w=3.34e-07 $l=1.88348e-07 $layer=LI1_cond $X=6.69 $Y=0.995
+ $X2=6.74 $Y2=1.16
r57 7 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.825 $Y=2.165
+ $X2=6.825 $Y2=1.325
r58 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.805 $Y=0.445
+ $X2=6.805 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A_788_316# 1 2 7 9 12 14 16 19 23 28 29 30 32
+ 33 37 40 41 44 47 53 59
c148 32 0 1.33968e-19 $X=7.2 $Y=1.495
c149 30 0 1.93706e-19 $X=6.845 $Y=1.58
c150 23 0 1.35566e-19 $X=4.095 $Y=0.51
r151 48 59 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.67 $Y=2.21 $X2=6.76
+ $Y2=2.21
r152 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.21
+ $X2=6.67 $Y2=2.21
r153 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.21
+ $X2=4.37 $Y2=2.21
r154 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.515 $Y=2.21
+ $X2=4.37 $Y2=2.21
r155 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.525 $Y=2.21
+ $X2=6.67 $Y2=2.21
r156 40 41 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=6.525 $Y=2.21
+ $X2=4.515 $Y2=2.21
r157 38 53 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.34 $Y=1.16
+ $X2=7.73 $Y2=1.16
r158 38 50 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.34 $Y=1.16 $X2=7.31
+ $Y2=1.16
r159 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.16 $X2=7.34 $Y2=1.16
r160 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.2 $Y=1.16
+ $X2=7.34 $Y2=1.16
r161 33 44 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.18 $Y=2.21
+ $X2=4.37 $Y2=2.21
r162 31 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.2 $Y=1.325
+ $X2=7.2 $Y2=1.16
r163 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.2 $Y=1.325
+ $X2=7.2 $Y2=1.495
r164 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.115 $Y=1.58
+ $X2=7.2 $Y2=1.495
r165 29 30 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.115 $Y=1.58
+ $X2=6.845 $Y2=1.58
r166 28 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.125
+ $X2=6.76 $Y2=2.21
r167 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.76 $Y=1.665
+ $X2=6.845 $Y2=1.58
r168 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.76 $Y=1.665
+ $X2=6.76 $Y2=2.125
r169 23 26 70.9234 $w=1.88e-07 $l=1.215e-06 $layer=LI1_cond $X=4.085 $Y=0.51
+ $X2=4.085 $Y2=1.725
r170 21 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.085 $Y=2.125
+ $X2=4.18 $Y2=2.21
r171 21 26 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=4.085 $Y=2.125
+ $X2=4.085 $Y2=1.725
r172 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.73 $Y=1.325
+ $X2=7.73 $Y2=1.16
r173 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.73 $Y=1.325
+ $X2=7.73 $Y2=1.985
r174 14 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.73 $Y=0.995
+ $X2=7.73 $Y2=1.16
r175 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.73 $Y=0.995
+ $X2=7.73 $Y2=0.56
r176 10 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=1.325
+ $X2=7.31 $Y2=1.16
r177 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.31 $Y=1.325
+ $X2=7.31 $Y2=1.985
r178 7 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.31 $Y=0.995
+ $X2=7.31 $Y2=1.16
r179 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.31 $Y=0.995
+ $X2=7.31 $Y2=0.56
r180 2 26 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.58 $X2=4.075 $Y2=1.725
r181 1 23 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.095 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42 43
+ 44 46 58 69 74 77 81
c130 4 0 1.33968e-19 $X=6.9 $Y=1.845
r131 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r132 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r133 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 72 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r135 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r136 69 80 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=8.107 $Y2=2.72
r137 69 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=2.72
+ $X2=7.59 $Y2=2.72
r138 68 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r139 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r140 65 68 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 65 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r142 64 67 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=6.67 $Y2=2.72
r143 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r144 62 77 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.1 $Y=2.72
+ $X2=4.927 $Y2=2.72
r145 62 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=2.72
+ $X2=5.29 $Y2=2.72
r146 61 78 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.83 $Y2=2.72
r147 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r148 58 77 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.755 $Y=2.72
+ $X2=4.927 $Y2=2.72
r149 58 60 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=4.755 $Y=2.72
+ $X2=2.99 $Y2=2.72
r150 57 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r151 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r152 54 57 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r153 54 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 53 56 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r155 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r156 51 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r157 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r158 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r159 46 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r160 44 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r161 44 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r162 42 67 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=6.67 $Y2=2.72
r163 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=7.1 $Y2=2.72
r164 41 71 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.185 $Y=2.72
+ $X2=7.59 $Y2=2.72
r165 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.185 $Y=2.72
+ $X2=7.1 $Y2=2.72
r166 39 56 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.595 $Y=2.72
+ $X2=2.53 $Y2=2.72
r167 39 40 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.595 $Y=2.72
+ $X2=2.71 $Y2=2.72
r168 38 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.99 $Y2=2.72
r169 38 40 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.825 $Y=2.72
+ $X2=2.71 $Y2=2.72
r170 34 37 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=8.06 $Y=1.66
+ $X2=8.06 $Y2=2.34
r171 32 80 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=8.06 $Y=2.635
+ $X2=8.107 $Y2=2.72
r172 32 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.06 $Y=2.635
+ $X2=8.06 $Y2=2.34
r173 28 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.1 $Y=2.635 $X2=7.1
+ $Y2=2.72
r174 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.1 $Y=2.635
+ $X2=7.1 $Y2=2
r175 24 77 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.927 $Y=2.635
+ $X2=4.927 $Y2=2.72
r176 24 26 13.1946 $w=3.43e-07 $l=3.95e-07 $layer=LI1_cond $X=4.927 $Y=2.635
+ $X2=4.927 $Y2=2.24
r177 20 40 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.72
r178 20 22 20.7941 $w=2.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.22
r179 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r180 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r181 5 37 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=7.805
+ $Y=1.485 $X2=8.02 $Y2=2.34
r182 5 34 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=7.805
+ $Y=1.485 $X2=8.02 $Y2=1.66
r183 4 30 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=6.9
+ $Y=1.845 $X2=7.1 $Y2=2
r184 3 26 600 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=1.845 $X2=5.015 $Y2=2.24
r185 2 22 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.725 $X2=2.715 $Y2=2.22
r186 1 18 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.845 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A_288_47# 1 2 3 4 13 17 22 24 25 26 28 33 35
+ 37 40 41 47
c132 47 0 2.0604e-19 $X=3.45 $Y=2.21
c133 22 0 2.70803e-20 $X=1.985 $Y=1.235
c134 13 0 7.52734e-20 $X=2.07 $Y=2.21
r135 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.21
+ $X2=3.45 $Y2=2.21
r136 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.21
+ $X2=2.07 $Y2=2.21
r137 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.215 $Y=2.21
+ $X2=2.07 $Y2=2.21
r138 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.305 $Y=2.21
+ $X2=3.45 $Y2=2.21
r139 40 41 1.34901 $w=1.4e-07 $l=1.09e-06 $layer=MET1_cond $X=3.305 $Y=2.21
+ $X2=2.215 $Y2=2.21
r140 37 39 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.702 $Y=0.51
+ $X2=3.702 $Y2=0.675
r141 35 39 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=3.735 $Y=1.81
+ $X2=3.735 $Y2=0.675
r142 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.985 $Y=1.32
+ $X2=2.155 $Y2=1.32
r143 26 48 15.7882 $w=1.68e-07 $l=2.42e-07 $layer=LI1_cond $X=3.692 $Y=2.21
+ $X2=3.45 $Y2=2.21
r144 26 28 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=3.692 $Y=2.125
+ $X2=3.692 $Y2=1.975
r145 25 35 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=3.692 $Y=1.937
+ $X2=3.692 $Y2=1.81
r146 25 28 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=3.692 $Y=1.937
+ $X2=3.692 $Y2=1.975
r147 24 44 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.125
+ $X2=2.155 $Y2=2.21
r148 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.405
+ $X2=2.155 $Y2=1.32
r149 23 24 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.155 $Y=1.405
+ $X2=2.155 $Y2=2.125
r150 22 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=1.235
+ $X2=1.985 $Y2=1.32
r151 21 22 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.985 $Y=0.535
+ $X2=1.985 $Y2=1.235
r152 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.9 $Y=0.45
+ $X2=1.985 $Y2=0.535
r153 17 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.9 $Y=0.45
+ $X2=1.635 $Y2=0.45
r154 13 44 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.21
+ $X2=2.155 $Y2=2.21
r155 13 15 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.07 $Y=2.21
+ $X2=1.575 $Y2=2.21
r156 4 28 600 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.58 $X2=3.655 $Y2=1.975
r157 3 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=2.065 $X2=1.575 $Y2=2.21
r158 2 37 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.235 $X2=3.67 $Y2=0.51
r159 1 19 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.635 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%A_872_316# 1 2 3 4 14 15 18 20 21 23 25 27 30
+ 35
r87 30 32 9.2829 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=4.497 $Y=0.42
+ $X2=4.497 $Y2=0.585
r88 25 27 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.495 $Y=2.24
+ $X2=6.11 $Y2=2.24
r89 21 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.495 $Y=0.38
+ $X2=6.055 $Y2=0.38
r90 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.41 $Y=2.155
+ $X2=5.495 $Y2=2.24
r91 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=1.735
+ $X2=5.41 $Y2=1.65
r92 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.41 $Y=1.735
+ $X2=5.41 $Y2=2.155
r93 18 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=1.565
+ $X2=5.41 $Y2=1.65
r94 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.41 $Y=0.465
+ $X2=5.495 $Y2=0.38
r95 17 18 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=5.41 $Y=0.465
+ $X2=5.41 $Y2=1.565
r96 16 34 3.40825 $w=1.7e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.585 $Y=1.65
+ $X2=4.49 $Y2=1.73
r97 15 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=1.65
+ $X2=5.41 $Y2=1.65
r98 15 16 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.325 $Y=1.65
+ $X2=4.585 $Y2=1.65
r99 14 34 3.40825 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.48 $Y=1.565
+ $X2=4.49 $Y2=1.73
r100 14 32 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=4.48 $Y=1.565
+ $X2=4.48 $Y2=0.585
r101 4 27 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=2.065 $X2=6.11 $Y2=2.24
r102 3 34 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.58 $X2=4.495 $Y2=1.73
r103 2 23 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=5.855
+ $Y=0.235 $X2=6.055 $Y2=0.38
r104 1 30 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.235 $X2=4.515 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%X 1 2 9 10 11 12 13 30
c31 10 0 1.09101e-19 $X=7.61 $Y=1.495
r32 30 31 1.69646 $w=4.08e-07 $l=3.5e-08 $layer=LI1_cond $X=7.56 $Y=1.87
+ $X2=7.56 $Y2=1.835
r33 13 20 4.77842 $w=4.08e-07 $l=1.7e-07 $layer=LI1_cond $X=7.56 $Y=2.21
+ $X2=7.56 $Y2=2.04
r34 12 20 4.07571 $w=4.08e-07 $l=1.45e-07 $layer=LI1_cond $X=7.56 $Y=1.895
+ $X2=7.56 $Y2=2.04
r35 12 30 0.702709 $w=4.08e-07 $l=2.5e-08 $layer=LI1_cond $X=7.56 $Y=1.895
+ $X2=7.56 $Y2=1.87
r36 12 31 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=7.61 $Y=1.81
+ $X2=7.61 $Y2=1.835
r37 11 28 13.0021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.6 $Y=0.43 $X2=7.6
+ $Y2=0.725
r38 10 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.68 $Y=1.495
+ $X2=7.68 $Y2=0.725
r39 9 12 5.94809 $w=3.08e-07 $l=1.6e-07 $layer=LI1_cond $X=7.61 $Y=1.65 $X2=7.61
+ $Y2=1.81
r40 9 10 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=7.61 $Y=1.65
+ $X2=7.61 $Y2=1.495
r41 2 12 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=7.385
+ $Y=1.485 $X2=7.52 $Y2=1.92
r42 1 11 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.235 $X2=7.52 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__MUX4_2%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 61 67 70 73 76 80
c130 80 0 1.64811e-19 $X=8.05 $Y=0
c131 43 0 1.47056e-19 $X=2.45 $Y=0
r132 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r133 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r134 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r135 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r136 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r137 65 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r138 65 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r139 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r140 62 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=0 $X2=7.14
+ $Y2=0
r141 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=7.59 $Y2=0
r142 61 79 4.08769 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=7.935 $Y=0
+ $X2=8.107 $Y2=0
r143 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r144 60 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r145 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r146 57 60 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r147 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r148 56 59 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=6.67
+ $Y2=0
r149 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r150 54 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r151 54 56 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0
+ $X2=5.29 $Y2=0
r152 53 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.015 $Y=0 $X2=7.14
+ $Y2=0
r153 53 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.015 $Y=0 $X2=6.67
+ $Y2=0
r154 52 74 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.83 $Y2=0
r155 52 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r156 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r157 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.615
+ $Y2=0
r158 49 51 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.99
+ $Y2=0
r159 48 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r160 48 51 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=2.99 $Y2=0
r161 47 71 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.53 $Y2=0
r162 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r163 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r164 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r165 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r166 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.615
+ $Y2=0
r167 43 46 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=2.45 $Y=0 $X2=1.15
+ $Y2=0
r168 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r169 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r170 36 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r171 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r172 32 79 3.08953 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.062 $Y=0.085
+ $X2=8.107 $Y2=0
r173 32 34 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=8.062 $Y=0.085
+ $X2=8.062 $Y2=0.38
r174 28 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0
r175 28 30 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0.51
r176 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r177 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.38
r178 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r179 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.38
r180 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r181 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r182 5 34 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=7.805
+ $Y=0.235 $X2=8.02 $Y2=0.38
r183 4 30 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=6.88
+ $Y=0.235 $X2=7.1 $Y2=0.51
r184 3 26 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.235 $X2=5.035 $Y2=0.38
r185 2 22 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.655 $Y2=0.38
r186 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__or3b_1.spice.SKY130_FD_SC_HD__OR3B_1.pxi
* Created: Thu Aug 27 14:43:38 2020
* 
x_PM_SKY130_FD_SC_HD__OR3B_1%C_N N_C_N_c_71_n N_C_N_M1009_g N_C_N_M1007_g C_N
+ N_C_N_c_73_n C_N PM_SKY130_FD_SC_HD__OR3B_1%C_N
x_PM_SKY130_FD_SC_HD__OR3B_1%A_109_93# N_A_109_93#_M1009_d N_A_109_93#_M1007_d
+ N_A_109_93#_M1005_g N_A_109_93#_M1000_g N_A_109_93#_c_94_n N_A_109_93#_c_95_n
+ N_A_109_93#_c_96_n N_A_109_93#_c_102_n N_A_109_93#_c_97_n
+ PM_SKY130_FD_SC_HD__OR3B_1%A_109_93#
x_PM_SKY130_FD_SC_HD__OR3B_1%B N_B_c_139_n N_B_M1002_g N_B_M1004_g N_B_c_137_n
+ N_B_c_138_n B B B N_B_c_141_n PM_SKY130_FD_SC_HD__OR3B_1%B
x_PM_SKY130_FD_SC_HD__OR3B_1%A N_A_c_178_n N_A_M1008_g N_A_M1006_g A A A
+ N_A_c_180_n N_A_c_181_n PM_SKY130_FD_SC_HD__OR3B_1%A
x_PM_SKY130_FD_SC_HD__OR3B_1%A_215_53# N_A_215_53#_M1005_s N_A_215_53#_M1004_d
+ N_A_215_53#_M1000_s N_A_215_53#_M1001_g N_A_215_53#_M1003_g
+ N_A_215_53#_c_230_n N_A_215_53#_c_231_n N_A_215_53#_c_232_n
+ N_A_215_53#_c_240_n N_A_215_53#_c_321_p N_A_215_53#_c_233_n
+ N_A_215_53#_c_278_n N_A_215_53#_c_241_n N_A_215_53#_c_242_n
+ N_A_215_53#_c_234_n N_A_215_53#_c_243_n N_A_215_53#_c_235_n
+ N_A_215_53#_c_236_n N_A_215_53#_c_237_n N_A_215_53#_c_238_n
+ PM_SKY130_FD_SC_HD__OR3B_1%A_215_53#
x_PM_SKY130_FD_SC_HD__OR3B_1%VPWR N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_c_331_n
+ N_VPWR_c_332_n N_VPWR_c_333_n VPWR N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_330_n N_VPWR_c_337_n PM_SKY130_FD_SC_HD__OR3B_1%VPWR
x_PM_SKY130_FD_SC_HD__OR3B_1%X N_X_M1001_d N_X_M1003_d N_X_c_367_n N_X_c_369_n
+ N_X_c_368_n X PM_SKY130_FD_SC_HD__OR3B_1%X
x_PM_SKY130_FD_SC_HD__OR3B_1%VGND N_VGND_M1009_s N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n VGND
+ N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n
+ N_VGND_c_394_n PM_SKY130_FD_SC_HD__OR3B_1%VGND
cc_1 VNB N_C_N_c_71_n 0.0213675f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB C_N 0.00874107f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_73_n 0.0409146f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_109_93#_M1005_g 0.0311233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_109_93#_c_94_n 0.0256218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_109_93#_c_95_n 0.010112f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_7 VNB N_A_109_93#_c_96_n 0.0131817f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_8 VNB N_A_109_93#_c_97_n 0.00573936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_M1002_g 0.016298f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_10 VNB N_B_c_137_n 0.013575f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_B_c_138_n 0.0110772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_c_178_n 0.0206627f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_13 VNB N_A_M1006_g 0.0265612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_c_180_n 0.00220933f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_15 VNB N_A_c_181_n 0.00354585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_215_53#_c_230_n 0.0088368f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_17 VNB N_A_215_53#_c_231_n 0.00375101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_215_53#_c_232_n 0.00351712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_215_53#_c_233_n 0.00111114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_215_53#_c_234_n 0.00147682f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_215_53#_c_235_n 0.00185649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_215_53#_c_236_n 0.0234012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_215_53#_c_237_n 0.00106484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_215_53#_c_238_n 0.019683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_330_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_367_n 0.0137601f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_27 VNB N_X_c_368_n 0.0241563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_385_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_29 VNB N_VGND_c_386_n 0.0388179f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_30 VNB N_VGND_c_387_n 0.00101984f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_31 VNB N_VGND_c_388_n 6.33915e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.0292709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_390_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_391_n 0.0166241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_392_n 0.199288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_393_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_394_n 0.00516646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VPB N_C_N_M1007_g 0.0287031f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_39 VPB C_N 8.94523e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_40 VPB N_C_N_c_73_n 0.0102214f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_41 VPB N_A_109_93#_M1000_g 0.0226299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_109_93#_c_94_n 0.00983741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_109_93#_c_95_n 6.52385e-19 $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_44 VPB N_A_109_93#_c_96_n 0.00352947f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_45 VPB N_A_109_93#_c_102_n 0.00453781f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_46 VPB N_A_109_93#_c_97_n 0.00573936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_B_c_139_n 0.0380443f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_48 VPB N_B_M1002_g 0.0241666f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_49 VPB N_B_c_141_n 0.0495672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_c_178_n 0.00403991f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_51 VPB N_A_M1008_g 0.021348f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.675
cc_52 VPB A 0.00149589f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_53 VPB N_A_c_180_n 0.00320355f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_54 VPB N_A_215_53#_M1003_g 0.0244726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_215_53#_c_240_n 0.00296402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_215_53#_c_241_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_215_53#_c_242_n 0.00814787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_215_53#_c_243_n 0.00130886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_215_53#_c_236_n 0.00544454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_331_n 0.00983572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_332_n 0.056538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_333_n 0.0114582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_334_n 0.0495055f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_64 VPB N_VPWR_c_335_n 0.0177135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_330_n 0.0670701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_337_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_X_c_369_n 0.00524127f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_68 VPB N_X_c_368_n 0.00880472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB X 0.032187f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_70 N_C_N_c_73_n N_A_109_93#_c_94_n 0.00702512f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C_N_c_71_n N_A_109_93#_c_96_n 0.0177192f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_72 C_N N_A_109_93#_c_96_n 0.0211231f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_73 N_C_N_M1007_g N_A_109_93#_c_102_n 0.00734101f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_74 N_C_N_c_71_n N_A_215_53#_c_230_n 0.00428704f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_75 N_C_N_M1007_g N_A_215_53#_c_242_n 0.00270689f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_76 N_C_N_M1007_g N_VPWR_c_332_n 0.00627879f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_77 C_N N_VPWR_c_332_n 0.0204657f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_78 N_C_N_c_73_n N_VPWR_c_332_n 0.0054329f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C_N_M1007_g N_VPWR_c_334_n 0.00327927f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_80 N_C_N_M1007_g N_VPWR_c_330_n 0.00417489f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_81 N_C_N_c_71_n N_VGND_c_386_n 0.00710775f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_82 C_N N_VGND_c_386_n 0.0210991f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_83 N_C_N_c_73_n N_VGND_c_386_n 0.00600816f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_84 N_C_N_c_71_n N_VGND_c_389_n 0.00483902f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_85 N_C_N_c_71_n N_VGND_c_392_n 0.00512902f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_109_93#_c_95_n N_B_M1002_g 0.0396727f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_109_93#_c_97_n N_B_M1002_g 2.39755e-19 $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_109_93#_M1005_g N_B_c_137_n 0.0136742f $X=1.41 $Y=0.475 $X2=0 $Y2=0
cc_89 N_A_109_93#_M1005_g N_B_c_138_n 0.0396727f $X=1.41 $Y=0.475 $X2=0 $Y2=0
cc_90 N_A_109_93#_M1000_g N_B_c_141_n 0.00442437f $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_91 N_A_109_93#_c_102_n N_B_c_141_n 0.0104825f $X=0.68 $Y=1.63 $X2=0 $Y2=0
cc_92 N_A_109_93#_M1000_g A 0.00440502f $X=1.41 $Y=1.695 $X2=0 $Y2=0
cc_93 N_A_109_93#_c_95_n N_A_c_181_n 0.0031188f $X=1.41 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_109_93#_c_97_n N_A_c_181_n 0.0245668f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_109_93#_M1005_g N_A_215_53#_c_230_n 9.90912e-19 $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_96 N_A_109_93#_c_96_n N_A_215_53#_c_230_n 0.0133756f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_97 N_A_109_93#_M1005_g N_A_215_53#_c_231_n 0.0170416f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_98 N_A_109_93#_c_94_n N_A_215_53#_c_231_n 0.00122152f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_99 N_A_109_93#_c_97_n N_A_215_53#_c_231_n 0.00184128f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_109_93#_c_94_n N_A_215_53#_c_232_n 0.00601607f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_109_93#_c_96_n N_A_215_53#_c_232_n 0.014504f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_102 N_A_109_93#_c_97_n N_A_215_53#_c_232_n 0.0216117f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_109_93#_M1000_g N_A_215_53#_c_240_n 0.0107819f $X=1.41 $Y=1.695 $X2=0
+ $Y2=0
cc_104 N_A_109_93#_M1000_g N_A_215_53#_c_242_n 0.00733409f $X=1.41 $Y=1.695
+ $X2=0 $Y2=0
cc_105 N_A_109_93#_c_94_n N_A_215_53#_c_242_n 0.00692982f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_A_109_93#_c_102_n N_A_215_53#_c_242_n 0.0224383f $X=0.68 $Y=1.63 $X2=0
+ $Y2=0
cc_107 N_A_109_93#_c_97_n N_A_215_53#_c_242_n 0.0214591f $X=1.135 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_109_93#_c_96_n N_VGND_c_386_n 0.0166146f $X=0.68 $Y=1.325 $X2=0 $Y2=0
cc_109 N_A_109_93#_M1005_g N_VGND_c_387_n 0.00789578f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_110 N_A_109_93#_M1005_g N_VGND_c_389_n 0.00322006f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_111 N_A_109_93#_c_96_n N_VGND_c_389_n 0.00840435f $X=0.68 $Y=1.325 $X2=0
+ $Y2=0
cc_112 N_A_109_93#_M1005_g N_VGND_c_392_n 0.00494938f $X=1.41 $Y=0.475 $X2=0
+ $Y2=0
cc_113 N_A_109_93#_c_96_n N_VGND_c_392_n 0.0109761f $X=0.68 $Y=1.325 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_c_178_n 0.0171538f $X=1.77 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_115 N_B_M1002_g N_A_M1008_g 0.025099f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_116 N_B_c_141_n N_A_M1008_g 8.99686e-19 $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_117 N_B_M1002_g N_A_M1006_g 0.00338246f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_118 N_B_c_137_n N_A_M1006_g 0.0187914f $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_119 N_B_M1002_g A 0.00846003f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_120 N_B_M1002_g N_A_c_180_n 0.00860145f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_121 N_B_c_138_n N_A_c_180_n 0.00177283f $X=1.8 $Y=0.91 $X2=0 $Y2=0
cc_122 N_B_M1002_g N_A_c_181_n 0.00540928f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_123 N_B_c_137_n N_A_215_53#_c_231_n 0.00683722f $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_124 N_B_c_138_n N_A_215_53#_c_231_n 0.00604464f $X=1.8 $Y=0.91 $X2=0 $Y2=0
cc_125 N_B_c_139_n N_A_215_53#_c_240_n 0.00120224f $X=1.77 $Y=2.145 $X2=0 $Y2=0
cc_126 N_B_M1002_g N_A_215_53#_c_240_n 0.0102586f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_127 N_B_c_141_n N_A_215_53#_c_240_n 0.050268f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_128 N_B_M1002_g N_A_215_53#_c_242_n 6.74356e-19 $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_129 N_B_c_141_n N_A_215_53#_c_242_n 0.0271442f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_130 N_B_M1002_g N_A_215_53#_c_243_n 0.00282377f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_131 N_B_c_141_n N_A_215_53#_c_243_n 0.0138251f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_132 N_B_c_141_n N_VPWR_c_332_n 0.0224011f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_133 N_B_c_139_n N_VPWR_c_333_n 7.16675e-19 $X=1.77 $Y=2.145 $X2=0 $Y2=0
cc_134 N_B_M1002_g N_VPWR_c_333_n 0.0025092f $X=1.77 $Y=1.695 $X2=0 $Y2=0
cc_135 N_B_c_141_n N_VPWR_c_333_n 0.0286775f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_136 N_B_c_139_n N_VPWR_c_334_n 0.00189221f $X=1.77 $Y=2.145 $X2=0 $Y2=0
cc_137 N_B_c_141_n N_VPWR_c_334_n 0.102616f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_138 N_B_c_141_n N_VPWR_c_330_n 0.0607178f $X=1.825 $Y=2.28 $X2=0 $Y2=0
cc_139 N_B_c_137_n N_VGND_c_387_n 0.00679416f $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_140 N_B_c_138_n N_VGND_c_387_n 2.19529e-19 $X=1.8 $Y=0.91 $X2=0 $Y2=0
cc_141 N_B_c_137_n N_VGND_c_388_n 5.25443e-19 $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_142 N_B_c_137_n N_VGND_c_390_n 0.00322006f $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_143 N_B_c_137_n N_VGND_c_392_n 0.00390029f $X=1.8 $Y=0.76 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_A_215_53#_M1003_g 0.0189405f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_145 N_A_c_180_n N_A_215_53#_c_231_n 0.0137749f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_181_n N_A_215_53#_c_231_n 0.0199192f $X=1.647 $Y=1.325 $X2=0 $Y2=0
cc_147 N_A_M1008_g N_A_215_53#_c_240_n 2.20055e-19 $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_148 A N_A_215_53#_c_240_n 0.0133453f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_149 N_A_c_180_n N_A_215_53#_c_240_n 0.00847219f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_178_n N_A_215_53#_c_233_n 0.00210922f $X=2.245 $Y=1.325 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_A_215_53#_c_233_n 0.0116153f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_152 N_A_c_180_n N_A_215_53#_c_233_n 0.016311f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_M1008_g N_A_215_53#_c_278_n 0.0112175f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_154 N_A_c_180_n N_A_215_53#_c_278_n 0.00969518f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_M1008_g N_A_215_53#_c_241_n 0.0034529f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_156 N_A_c_178_n N_A_215_53#_c_234_n 5.36764e-19 $X=2.245 $Y=1.325 $X2=0 $Y2=0
cc_157 N_A_c_180_n N_A_215_53#_c_234_n 0.0146459f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_c_178_n N_A_215_53#_c_243_n 0.00156674f $X=2.245 $Y=1.325 $X2=0 $Y2=0
cc_159 N_A_M1008_g N_A_215_53#_c_243_n 0.0100503f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_160 A N_A_215_53#_c_243_n 0.00624989f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_161 N_A_c_180_n N_A_215_53#_c_243_n 0.0112207f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_c_178_n N_A_215_53#_c_235_n 0.00186306f $X=2.245 $Y=1.325 $X2=0 $Y2=0
cc_163 N_A_c_180_n N_A_215_53#_c_235_n 0.0271506f $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_178_n N_A_215_53#_c_236_n 0.0202654f $X=2.245 $Y=1.325 $X2=0 $Y2=0
cc_165 N_A_c_180_n N_A_215_53#_c_236_n 3.55971e-19 $X=2.23 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_M1006_g N_A_215_53#_c_237_n 0.00346594f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_167 N_A_M1006_g N_A_215_53#_c_238_n 0.0175873f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_168 N_A_M1008_g N_VPWR_c_333_n 0.00293484f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_169 N_A_M1008_g N_VPWR_c_334_n 0.00264181f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_170 N_A_M1008_g N_VPWR_c_330_n 0.00333991f $X=2.245 $Y=1.695 $X2=0 $Y2=0
cc_171 A A_297_297# 0.00106198f $X=1.525 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_172 N_A_M1006_g N_VGND_c_387_n 5.2354e-19 $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_173 N_A_M1006_g N_VGND_c_388_n 0.00707341f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_174 N_A_M1006_g N_VGND_c_390_n 0.00322006f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_175 N_A_M1006_g N_VGND_c_392_n 0.00390029f $X=2.25 $Y=0.475 $X2=0 $Y2=0
cc_176 N_A_215_53#_c_278_n N_VPWR_M1008_d 0.00526233f $X=2.52 $Y=1.58 $X2=0
+ $Y2=0
cc_177 N_A_215_53#_M1003_g N_VPWR_c_333_n 0.00485906f $X=2.735 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_215_53#_c_278_n N_VPWR_c_333_n 0.0190361f $X=2.52 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A_215_53#_c_243_n N_VPWR_c_333_n 0.00605542f $X=2.115 $Y=1.58 $X2=0
+ $Y2=0
cc_180 N_A_215_53#_c_236_n N_VPWR_c_333_n 2.11345e-19 $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_215_53#_M1003_g N_VPWR_c_335_n 0.00585385f $X=2.735 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_215_53#_M1003_g N_VPWR_c_330_n 0.0128443f $X=2.735 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_215_53#_c_240_n A_297_297# 0.0010205f $X=2.03 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A_215_53#_c_240_n A_369_297# 0.0024965f $X=2.03 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_185 N_A_215_53#_c_243_n A_369_297# 0.00476392f $X=2.115 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_186 N_A_215_53#_M1003_g N_X_c_368_n 0.00349311f $X=2.735 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_215_53#_c_233_n N_X_c_368_n 0.0035218f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_215_53#_c_241_n N_X_c_368_n 0.00841221f $X=2.605 $Y=1.495 $X2=0 $Y2=0
cc_189 N_A_215_53#_c_235_n N_X_c_368_n 0.024459f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_215_53#_c_236_n N_X_c_368_n 0.00753248f $X=2.71 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_215_53#_c_237_n N_X_c_368_n 0.00836618f $X=2.657 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_215_53#_c_238_n N_X_c_368_n 0.00441003f $X=2.71 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_215_53#_c_231_n N_VGND_M1005_d 0.00160115f $X=1.955 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_215_53#_c_233_n N_VGND_M1006_d 0.00467744f $X=2.52 $Y=0.74 $X2=0
+ $Y2=0
cc_195 N_A_215_53#_c_237_n N_VGND_M1006_d 6.96297e-19 $X=2.657 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A_215_53#_c_230_n N_VGND_c_387_n 0.00899132f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_197 N_A_215_53#_c_231_n N_VGND_c_387_n 0.0160613f $X=1.955 $Y=0.74 $X2=0
+ $Y2=0
cc_198 N_A_215_53#_c_233_n N_VGND_c_388_n 0.0203172f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_215_53#_c_236_n N_VGND_c_388_n 2.33671e-19 $X=2.71 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_215_53#_c_238_n N_VGND_c_388_n 0.0132163f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_215_53#_c_230_n N_VGND_c_389_n 0.0182527f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_202 N_A_215_53#_c_231_n N_VGND_c_389_n 0.0023303f $X=1.955 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_A_215_53#_c_231_n N_VGND_c_390_n 0.00232396f $X=1.955 $Y=0.74 $X2=0
+ $Y2=0
cc_204 N_A_215_53#_c_321_p N_VGND_c_390_n 0.00846569f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_205 N_A_215_53#_c_233_n N_VGND_c_390_n 0.00232396f $X=2.52 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_215_53#_c_233_n N_VGND_c_391_n 3.34073e-19 $X=2.52 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_215_53#_c_238_n N_VGND_c_391_n 0.00524631f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_215_53#_c_230_n N_VGND_c_392_n 0.00989054f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_209 N_A_215_53#_c_231_n N_VGND_c_392_n 0.00971545f $X=1.955 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_215_53#_c_321_p N_VGND_c_392_n 0.00625722f $X=2.04 $Y=0.47 $X2=0
+ $Y2=0
cc_211 N_A_215_53#_c_233_n N_VGND_c_392_n 0.00635763f $X=2.52 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_215_53#_c_238_n N_VGND_c_392_n 0.00951738f $X=2.71 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_330_n N_X_M1003_d 0.00399469f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_335_n X 0.0190559f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_c_330_n X 0.0105137f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_216 N_X_c_367_n N_VGND_c_391_n 0.00892672f $X=3.05 $Y=0.587 $X2=0 $Y2=0
cc_217 N_X_M1001_d N_VGND_c_392_n 0.00416042f $X=2.81 $Y=0.235 $X2=0 $Y2=0
cc_218 N_X_c_367_n N_VGND_c_392_n 0.00941771f $X=3.05 $Y=0.587 $X2=0 $Y2=0

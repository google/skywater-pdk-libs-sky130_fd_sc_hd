* File: sky130_fd_sc_hd__ebufn_1.spice.SKY130_FD_SC_HD__EBUFN_1.pxi
* Created: Thu Aug 27 14:19:19 2020
* 
x_PM_SKY130_FD_SC_HD__EBUFN_1%A N_A_M1005_g N_A_M1003_g A A N_A_c_63_n
+ PM_SKY130_FD_SC_HD__EBUFN_1%A
x_PM_SKY130_FD_SC_HD__EBUFN_1%TE_B N_TE_B_M1001_g N_TE_B_c_88_n N_TE_B_M1007_g
+ N_TE_B_M1004_g N_TE_B_c_89_n N_TE_B_c_90_n TE_B TE_B
+ PM_SKY130_FD_SC_HD__EBUFN_1%TE_B
x_PM_SKY130_FD_SC_HD__EBUFN_1%A_193_369# N_A_193_369#_M1007_d
+ N_A_193_369#_M1001_d N_A_193_369#_c_137_n N_A_193_369#_M1002_g
+ N_A_193_369#_c_142_n N_A_193_369#_c_138_n N_A_193_369#_c_143_n
+ N_A_193_369#_c_139_n N_A_193_369#_c_140_n N_A_193_369#_c_156_n
+ N_A_193_369#_c_141_n PM_SKY130_FD_SC_HD__EBUFN_1%A_193_369#
x_PM_SKY130_FD_SC_HD__EBUFN_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1003_s
+ N_A_27_47#_M1006_g N_A_27_47#_M1000_g N_A_27_47#_c_193_n N_A_27_47#_c_205_n
+ N_A_27_47#_c_194_n N_A_27_47#_c_224_n N_A_27_47#_c_195_n N_A_27_47#_c_217_n
+ N_A_27_47#_c_196_n N_A_27_47#_c_197_n N_A_27_47#_c_198_n N_A_27_47#_c_199_n
+ N_A_27_47#_c_200_n N_A_27_47#_c_207_n N_A_27_47#_c_201_n N_A_27_47#_c_202_n
+ N_A_27_47#_c_203_n PM_SKY130_FD_SC_HD__EBUFN_1%A_27_47#
x_PM_SKY130_FD_SC_HD__EBUFN_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_s N_VPWR_c_305_n
+ N_VPWR_c_306_n VPWR N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_304_n N_VPWR_c_311_n N_VPWR_c_312_n PM_SKY130_FD_SC_HD__EBUFN_1%VPWR
x_PM_SKY130_FD_SC_HD__EBUFN_1%Z N_Z_M1006_d N_Z_M1000_d Z Z Z Z Z Z Z
+ N_Z_c_353_n N_Z_c_351_n Z N_Z_c_350_n PM_SKY130_FD_SC_HD__EBUFN_1%Z
x_PM_SKY130_FD_SC_HD__EBUFN_1%VGND N_VGND_M1005_d N_VGND_M1002_s N_VGND_c_379_n
+ VGND N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n
+ N_VGND_c_384_n N_VGND_c_385_n PM_SKY130_FD_SC_HD__EBUFN_1%VGND
cc_1 VNB N_A_M1005_g 0.0382186f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.0137853f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_c_63_n 0.0336001f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_TE_B_c_88_n 0.030021f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_5 VNB N_TE_B_c_89_n 0.0159446f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_6 VNB N_TE_B_c_90_n 0.0583658f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_A_193_369#_c_137_n 0.0194389f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.165
cc_8 VNB N_A_193_369#_c_138_n 0.00467887f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_9 VNB N_A_193_369#_c_139_n 0.00295737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_193_369#_c_140_n 0.0031322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_193_369#_c_141_n 0.0303691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_193_n 0.0132408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_194_n 0.00347289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_195_n 0.0118279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_196_n 0.02026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_197_n 9.80023e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_198_n 0.00797971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_199_n 0.0069638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_200_n 0.00396693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_201_n 0.00561681f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_202_n 0.0235061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_203_n 0.0177457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_304_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB Z 0.0260135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Z_c_350_n 0.026125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_379_n 0.0043076f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_VGND_c_380_n 0.0143746f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_28 VNB N_VGND_c_381_n 0.0197588f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_382_n 0.210732f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_383_n 0.00506674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_384_n 0.0318824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_385_n 0.0137805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_M1003_g 0.04382f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.165
cc_34 VPB A 0.0164877f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_35 VPB N_A_c_63_n 0.00918023f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_36 VPB N_TE_B_M1001_g 0.0451227f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_37 VPB N_TE_B_M1004_g 0.0295458f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_38 VPB N_TE_B_c_89_n 8.85159e-19 $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_39 VPB N_TE_B_c_90_n 0.020063f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_40 VPB TE_B 0.00674563f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_41 VPB N_A_193_369#_c_142_n 0.00550333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_193_369#_c_143_n 0.0150089f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_43 VPB N_A_193_369#_c_139_n 0.00456577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_193_369#_c_141_n 0.0119577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_M1000_g 0.0296819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_205_n 0.0179778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_194_n 0.0040448f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_207_n 0.0130872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_201_n 0.00225912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_202_n 0.00443776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_305_n 4.10133e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_52 VPB N_VPWR_c_306_n 0.00575184f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_53 VPB N_VPWR_c_307_n 0.0144009f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_54 VPB N_VPWR_c_308_n 0.0148099f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.53
cc_55 VPB N_VPWR_c_309_n 0.0453881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_304_n 0.0486892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.00436611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_312_n 0.00569002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_Z_c_351_n 0.0509353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB Z 0.01123f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 N_A_M1003_g N_TE_B_M1001_g 0.0286267f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_TE_B_c_88_n 0.0195145f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_c_63_n N_TE_B_c_89_n 0.0286267f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_c_63_n TE_B 4.43686e-19 $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1005_g N_A_27_47#_c_194_n 0.00869167f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_A_27_47#_c_194_n 0.0138015f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_67 A N_A_27_47#_c_194_n 0.0454615f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_c_63_n N_A_27_47#_c_194_n 0.00785916f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_A_27_47#_c_195_n 0.0186376f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_70 A N_A_27_47#_c_195_n 0.0218104f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_c_63_n N_A_27_47#_c_195_n 0.0031434f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_A_27_47#_c_217_n 2.64984e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_A_27_47#_c_207_n 0.0187297f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_207_n 0.0228675f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_63_n N_A_27_47#_c_207_n 0.0019986f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_VPWR_c_305_n 0.00919555f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_77 N_A_M1003_g N_VPWR_c_307_n 0.00348405f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_78 N_A_M1003_g N_VPWR_c_304_n 0.00513647f $X=0.47 $Y=2.165 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_VGND_c_379_n 0.00973188f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_80 N_A_M1005_g N_VGND_c_380_n 0.00337001f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_VGND_c_382_n 0.00493924f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_82 N_TE_B_M1004_g N_A_193_369#_c_142_n 0.00341043f $X=1.84 $Y=1.985 $X2=0
+ $Y2=0
cc_83 N_TE_B_c_88_n N_A_193_369#_c_138_n 0.0021256f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_84 N_TE_B_c_90_n N_A_193_369#_c_138_n 0.0113232f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_85 N_TE_B_M1001_g N_A_193_369#_c_143_n 0.00850888f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_86 N_TE_B_M1004_g N_A_193_369#_c_143_n 0.029281f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_87 N_TE_B_c_90_n N_A_193_369#_c_143_n 0.00606406f $X=1.765 $Y=1.16 $X2=0
+ $Y2=0
cc_88 TE_B N_A_193_369#_c_143_n 0.044553f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_89 N_TE_B_c_90_n N_A_193_369#_c_139_n 0.0122035f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_90 N_TE_B_c_88_n N_A_193_369#_c_140_n 0.00226565f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_91 N_TE_B_c_90_n N_A_193_369#_c_140_n 0.00226247f $X=1.765 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_TE_B_c_90_n N_A_193_369#_c_156_n 0.0209048f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_93 TE_B N_A_193_369#_c_156_n 0.0199562f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_94 N_TE_B_c_90_n N_A_193_369#_c_141_n 0.0136095f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_95 N_TE_B_c_88_n N_A_27_47#_c_194_n 0.00198111f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_96 N_TE_B_c_89_n N_A_27_47#_c_194_n 0.00730791f $X=0.932 $Y=1.16 $X2=0 $Y2=0
cc_97 TE_B N_A_27_47#_c_194_n 0.0424281f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 N_TE_B_c_88_n N_A_27_47#_c_224_n 0.0147309f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_99 N_TE_B_c_89_n N_A_27_47#_c_224_n 0.00256391f $X=0.932 $Y=1.16 $X2=0 $Y2=0
cc_100 N_TE_B_c_90_n N_A_27_47#_c_224_n 0.00304871f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_101 TE_B N_A_27_47#_c_224_n 0.0144816f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_102 N_TE_B_c_88_n N_A_27_47#_c_217_n 0.00559256f $X=0.975 $Y=0.995 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_90_n N_A_27_47#_c_196_n 0.0084907f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_104 TE_B N_A_27_47#_c_196_n 0.00160979f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_105 N_TE_B_c_88_n N_A_27_47#_c_197_n 0.0077697f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_106 N_TE_B_c_90_n N_A_27_47#_c_200_n 0.00179376f $X=1.765 $Y=1.16 $X2=0 $Y2=0
cc_107 N_TE_B_M1001_g N_A_27_47#_c_207_n 0.00217457f $X=0.89 $Y=2.165 $X2=0
+ $Y2=0
cc_108 N_TE_B_M1001_g N_VPWR_c_305_n 0.00893175f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_109 N_TE_B_M1001_g N_VPWR_c_306_n 0.00217989f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_110 N_TE_B_M1004_g N_VPWR_c_306_n 0.0116894f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_111 N_TE_B_M1001_g N_VPWR_c_308_n 0.0046653f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_112 N_TE_B_M1004_g N_VPWR_c_309_n 0.00427505f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_113 N_TE_B_M1001_g N_VPWR_c_304_n 0.00934473f $X=0.89 $Y=2.165 $X2=0 $Y2=0
cc_114 N_TE_B_M1004_g N_VPWR_c_304_n 0.00873046f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_115 N_TE_B_M1004_g N_Z_c_353_n 0.026188f $X=1.84 $Y=1.985 $X2=0 $Y2=0
cc_116 N_TE_B_c_88_n N_VGND_c_379_n 0.0030314f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_117 N_TE_B_c_88_n N_VGND_c_382_n 0.00510711f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_118 N_TE_B_c_88_n N_VGND_c_384_n 0.00341702f $X=0.975 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_193_369#_c_138_n N_A_27_47#_c_194_n 0.00538875f $X=1.547 $Y=1.075
+ $X2=0 $Y2=0
cc_120 N_A_193_369#_c_143_n N_A_27_47#_c_194_n 0.00480517f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_121 N_A_193_369#_c_140_n N_A_27_47#_c_194_n 0.0017713f $X=1.52 $Y=0.76 $X2=0
+ $Y2=0
cc_122 N_A_193_369#_M1007_d N_A_27_47#_c_224_n 0.00329588f $X=1.05 $Y=0.465
+ $X2=0 $Y2=0
cc_123 N_A_193_369#_c_140_n N_A_27_47#_c_224_n 0.016181f $X=1.52 $Y=0.76 $X2=0
+ $Y2=0
cc_124 N_A_193_369#_M1007_d N_A_27_47#_c_217_n 0.00296563f $X=1.05 $Y=0.465
+ $X2=0 $Y2=0
cc_125 N_A_193_369#_c_137_n N_A_27_47#_c_196_n 8.64558e-19 $X=2.58 $Y=0.995
+ $X2=0 $Y2=0
cc_126 N_A_193_369#_c_139_n N_A_27_47#_c_196_n 0.00139349f $X=2.37 $Y=1.16 $X2=0
+ $Y2=0
cc_127 N_A_193_369#_c_140_n N_A_27_47#_c_196_n 0.0257699f $X=1.52 $Y=0.76 $X2=0
+ $Y2=0
cc_128 N_A_193_369#_c_156_n N_A_27_47#_c_196_n 0.00365147f $X=1.607 $Y=1.2 $X2=0
+ $Y2=0
cc_129 N_A_193_369#_c_137_n N_A_27_47#_c_198_n 0.0045733f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_130 N_A_193_369#_c_140_n N_A_27_47#_c_198_n 0.0078909f $X=1.52 $Y=0.76 $X2=0
+ $Y2=0
cc_131 N_A_193_369#_c_137_n N_A_27_47#_c_199_n 0.0131208f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_A_193_369#_c_139_n N_A_27_47#_c_199_n 0.0382161f $X=2.37 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_193_369#_c_141_n N_A_27_47#_c_199_n 0.00665475f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_193_369#_c_139_n N_A_27_47#_c_200_n 0.0144531f $X=2.37 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_193_369#_c_140_n N_A_27_47#_c_200_n 0.014975f $X=1.52 $Y=0.76 $X2=0
+ $Y2=0
cc_136 N_A_193_369#_c_143_n N_A_27_47#_c_207_n 0.00834979f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_137 N_A_193_369#_c_137_n N_A_27_47#_c_201_n 0.00640393f $X=2.58 $Y=0.995
+ $X2=0 $Y2=0
cc_138 N_A_193_369#_c_139_n N_A_27_47#_c_201_n 0.0211345f $X=2.37 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_193_369#_c_141_n N_A_27_47#_c_202_n 0.0385312f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_193_369#_c_137_n N_A_27_47#_c_203_n 0.0385312f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_141 N_A_193_369#_c_143_n N_VPWR_M1004_s 0.00590922f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_142 N_A_193_369#_c_142_n N_VPWR_c_306_n 0.0234595f $X=1.1 $Y=2.265 $X2=0
+ $Y2=0
cc_143 N_A_193_369#_c_143_n N_VPWR_c_306_n 0.0241089f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_144 N_A_193_369#_c_142_n N_VPWR_c_308_n 0.0166106f $X=1.1 $Y=2.265 $X2=0
+ $Y2=0
cc_145 N_A_193_369#_c_143_n N_VPWR_c_308_n 0.00269444f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_146 N_A_193_369#_M1001_d N_VPWR_c_304_n 0.00383011f $X=0.965 $Y=1.845 $X2=0
+ $Y2=0
cc_147 N_A_193_369#_c_142_n N_VPWR_c_304_n 0.00961964f $X=1.1 $Y=2.265 $X2=0
+ $Y2=0
cc_148 N_A_193_369#_c_143_n N_VPWR_c_304_n 0.00607035f $X=1.607 $Y=1.8 $X2=0
+ $Y2=0
cc_149 N_A_193_369#_c_143_n N_Z_c_353_n 0.0431665f $X=1.607 $Y=1.8 $X2=0 $Y2=0
cc_150 N_A_193_369#_c_139_n N_Z_c_353_n 0.0461904f $X=2.37 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_193_369#_c_141_n N_Z_c_353_n 0.011083f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_193_369#_c_137_n N_VGND_c_385_n 0.0248045f $X=2.58 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_207_n N_VPWR_M1003_d 0.0032019f $X=0.632 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_27_47#_c_207_n N_VPWR_c_305_n 0.0130719f $X=0.632 $Y=1.895 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_205_n N_VPWR_c_307_n 0.0175014f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_207_n N_VPWR_c_307_n 0.00207512f $X=0.632 $Y=1.895 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_M1000_g N_VPWR_c_309_n 0.00357877f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_M1003_s N_VPWR_c_304_n 0.00234717f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_M1000_g N_VPWR_c_304_n 0.00781618f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_205_n N_VPWR_c_304_n 0.00983733f $X=0.26 $Y=2.22 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_207_n N_VPWR_c_304_n 0.00493223f $X=0.632 $Y=1.895 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_M1000_g N_Z_c_353_n 0.0458967f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_199_n N_Z_c_353_n 0.00521932f $X=2.705 $Y=0.82 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_201_n N_Z_c_353_n 0.0274474f $X=2.895 $Y=0.82 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_202_n N_Z_c_353_n 0.00247161f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1000_g Z 0.00583687f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_201_n Z 0.0354253f $X=2.895 $Y=0.82 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_202_n Z 0.00766586f $X=3 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_203_n Z 0.00328239f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_201_n N_Z_c_350_n 0.00761256f $X=2.895 $Y=0.82 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_202_n N_Z_c_350_n 2.66949e-19 $X=3 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_203_n N_Z_c_350_n 0.0155195f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_194_n N_VGND_M1005_d 0.00121069f $X=0.632 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_27_47#_c_224_n N_VGND_M1005_d 0.0042757f $X=1.015 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_27_47#_c_195_n N_VGND_M1005_d 0.00176688f $X=0.74 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_27_47#_c_199_n N_VGND_M1002_s 0.00481109f $X=2.705 $Y=0.82 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_195_n N_VGND_c_379_n 0.0206099f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_197_n N_VGND_c_379_n 0.0159418f $X=1.185 $Y=0.36 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_193_n N_VGND_c_380_n 0.0147634f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_195_n N_VGND_c_380_n 0.00261327f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_203_n N_VGND_c_381_n 0.00232377f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1005_s N_VGND_c_382_n 0.0022816f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_193_n N_VGND_c_382_n 0.00962926f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_224_n N_VGND_c_382_n 0.00439315f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_195_n N_VGND_c_382_n 0.00594195f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_196_n N_VGND_c_382_n 0.0315989f $X=1.855 $Y=0.36 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_197_n N_VGND_c_382_n 0.00635703f $X=1.185 $Y=0.36 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_199_n N_VGND_c_382_n 0.00631289f $X=2.705 $Y=0.82 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_201_n N_VGND_c_382_n 0.00101658f $X=2.895 $Y=0.82 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_203_n N_VGND_c_382_n 0.00550891f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_224_n N_VGND_c_384_n 0.00254828f $X=1.015 $Y=0.72 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_196_n N_VGND_c_384_n 0.055889f $X=1.855 $Y=0.36 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_197_n N_VGND_c_384_n 0.0119068f $X=1.185 $Y=0.36 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_199_n N_VGND_c_384_n 0.00249653f $X=2.705 $Y=0.82 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_196_n N_VGND_c_385_n 0.019305f $X=1.855 $Y=0.36 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_198_n N_VGND_c_385_n 0.0081484f $X=1.94 $Y=0.735 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_199_n N_VGND_c_385_n 0.0307107f $X=2.705 $Y=0.82 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_201_n N_VGND_c_385_n 0.0154057f $X=2.895 $Y=0.82 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_203_n N_VGND_c_385_n 0.0160782f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_201_n A_531_47# 0.00103579f $X=2.895 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_201 N_VPWR_c_304_n A_383_297# 0.00981138f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_202 N_VPWR_c_304_n N_Z_M1000_d 0.00255234f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_306_n N_Z_c_353_n 0.0240347f $X=1.62 $Y=2.26 $X2=0 $Y2=0
cc_204 N_VPWR_c_309_n N_Z_c_353_n 0.0851375f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_205 N_VPWR_c_304_n N_Z_c_353_n 0.0485804f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_206 N_VPWR_c_309_n N_Z_c_351_n 0.0242022f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_207 N_VPWR_c_304_n N_Z_c_351_n 0.0130835f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_208 A_383_297# N_Z_c_353_n 0.0638111f $X=1.915 $Y=1.485 $X2=3.45 $Y2=2.72
cc_209 N_Z_c_350_n N_VGND_c_381_n 0.032985f $X=3.29 $Y=0.36 $X2=0 $Y2=0
cc_210 N_Z_M1006_d N_VGND_c_382_n 0.00745383f $X=3.015 $Y=0.235 $X2=0 $Y2=0
cc_211 N_Z_c_350_n N_VGND_c_382_n 0.0180008f $X=3.29 $Y=0.36 $X2=0 $Y2=0
cc_212 N_Z_c_350_n N_VGND_c_385_n 0.0261365f $X=3.29 $Y=0.36 $X2=0 $Y2=0
cc_213 N_VGND_c_385_n A_531_47# 0.00106341f $X=2.955 $Y=0.24 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__and2b_1.pex.spice
* Created: Thu Aug 27 14:07:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND2B_1%A_N 3 7 9 10 11 16
c30 16 0 1.89169e-19 $X=0.36 $Y=1.16
r31 16 19 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.37 $Y=1.16
+ $X2=0.37 $Y2=1.325
r32 16 18 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.37 $Y=1.16
+ $X2=0.37 $Y2=0.995
r33 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r34 10 11 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.53
r35 10 17 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.16
r36 9 17 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.295 $Y=0.85
+ $X2=0.295 $Y2=1.16
r37 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r38 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%A_27_413# 1 2 9 13 17 19 20 22 24 26 33 34
c64 34 0 1.56867e-21 $X=1.065 $Y=0.97
c65 33 0 1.26328e-19 $X=1.065 $Y=0.97
c66 19 0 2.5987e-19 $X=0.615 $Y=1.9
c67 9 0 1.69139e-19 $X=0.96 $Y=2.275
r68 34 36 20.004 $w=2.53e-07 $l=1.05e-07 $layer=POLY_cond $X=1.065 $Y=0.97
+ $X2=0.96 $Y2=0.97
r69 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.065
+ $Y=0.97 $X2=1.065 $Y2=0.97
r70 31 33 11.6292 $w=3.28e-07 $l=3.33e-07 $layer=LI1_cond $X=0.732 $Y=0.97
+ $X2=1.065 $Y2=0.97
r71 29 31 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=0.725 $Y=0.97
+ $X2=0.732 $Y2=0.97
r72 26 28 10.1849 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.715 $Y=0.445
+ $X2=0.715 $Y2=0.655
r73 23 31 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.732 $Y=1.135
+ $X2=0.732 $Y2=0.97
r74 23 24 31.8761 $w=2.33e-07 $l=6.5e-07 $layer=LI1_cond $X=0.732 $Y=1.135
+ $X2=0.732 $Y2=1.785
r75 22 29 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.97
r76 22 28 7.85757 $w=2.18e-07 $l=1.5e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=0.655
r77 19 24 6.81752 $w=2.3e-07 $l=1.64754e-07 $layer=LI1_cond $X=0.615 $Y=1.9
+ $X2=0.732 $Y2=1.785
r78 19 20 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.615 $Y=1.9
+ $X2=0.345 $Y2=1.9
r79 15 20 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.345 $Y2=1.9
r80 15 17 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=2.225
r81 11 34 65.7273 $w=2.53e-07 $l=4.19464e-07 $layer=POLY_cond $X=1.41 $Y=0.805
+ $X2=1.065 $Y2=0.97
r82 11 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.41 $Y=0.805
+ $X2=1.41 $Y2=0.445
r83 7 36 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.135
+ $X2=0.96 $Y2=0.97
r84 7 9 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=0.96 $Y=1.135
+ $X2=0.96 $Y2=2.275
r85 2 17 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.225
r86 1 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%B 1 3 7 9 10
c32 10 0 1.70708e-19 $X=2.07 $Y=1.87
c33 7 0 1.26328e-19 $X=1.8 $Y=0.445
c34 1 0 1.16262e-19 $X=1.4 $Y=1.895
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.73 $X2=1.645 $Y2=1.73
r36 10 15 15.7996 $w=3.08e-07 $l=4.25e-07 $layer=LI1_cond $X=2.07 $Y=1.8
+ $X2=1.645 $Y2=1.8
r37 9 15 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=1.61 $Y=1.8 $X2=1.645
+ $Y2=1.8
r38 5 14 83.5248 $w=4.5e-07 $l=6.57438e-07 $layer=POLY_cond $X=1.8 $Y=1.165
+ $X2=1.6 $Y2=1.73
r39 5 7 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.8 $Y=1.165 $X2=1.8
+ $Y2=0.445
r40 1 14 40.6804 $w=4.5e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.4 $Y=1.895
+ $X2=1.6 $Y2=1.73
r41 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.4 $Y=1.895 $X2=1.4
+ $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%A_207_413# 1 2 9 12 16 19 20 22 23 28 31
r58 28 29 9.61923 $w=2.6e-07 $l=2.05e-07 $layer=LI1_cond $X=1.2 $Y=0.44
+ $X2=1.405 $Y2=0.44
r59 23 32 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.225 $Y2=1.325
r60 23 31 50.3433 $w=2.8e-07 $l=1.75e-07 $layer=POLY_cond $X=2.225 $Y=1.16
+ $X2=2.225 $Y2=0.985
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.16 $X2=2.22 $Y2=1.16
r62 20 26 14.4021 $w=4.04e-07 $l=5.11126e-07 $layer=LI1_cond $X=1.88 $Y=1.135
+ $X2=1.405 $Y2=1.21
r63 20 22 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.88 $Y=1.135
+ $X2=2.22 $Y2=1.135
r64 19 26 5.83894 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.405 $Y=0.945
+ $X2=1.405 $Y2=1.21
r65 18 29 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.405 $Y=0.61
+ $X2=1.405 $Y2=0.44
r66 18 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.405 $Y=0.61
+ $X2=1.405 $Y2=0.945
r67 14 26 7.33812 $w=4.04e-07 $l=3.66906e-07 $layer=LI1_cond $X=1.162 $Y=1.475
+ $X2=1.405 $Y2=1.21
r68 14 16 30.3274 $w=2.83e-07 $l=7.5e-07 $layer=LI1_cond $X=1.162 $Y=1.475
+ $X2=1.162 $Y2=2.225
r69 12 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.29 $Y=1.985
+ $X2=2.29 $Y2=1.325
r70 9 31 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.29 $Y=0.56
+ $X2=2.29 $Y2=0.985
r71 2 16 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=2.065 $X2=1.18 $Y2=2.225
r72 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%VPWR 1 2 9 11 13 25 26 29 33 37
c36 33 0 7.07005e-20 $X=1.485 $Y=2.485
c37 26 0 1.16262e-19 $X=2.53 $Y=2.72
r38 35 37 9.20209 $w=6.38e-07 $l=1e-07 $layer=LI1_cond $X=2.07 $Y=2.485 $X2=2.17
+ $Y2=2.485
r39 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 32 35 1.30821 $w=6.38e-07 $l=7e-08 $layer=LI1_cond $X=2 $Y=2.485 $X2=2.07
+ $Y2=2.485
r41 32 33 16.9579 $w=6.38e-07 $l=5.15e-07 $layer=LI1_cond $X=2 $Y=2.485
+ $X2=1.485 $Y2=2.485
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 26 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 25 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.17 $Y2=2.72
r45 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 22 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 22 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 21 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.485 $Y2=2.72
r49 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 19 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r51 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r52 13 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r53 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 11 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 7 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r57 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.27
r58 2 32 300 $w=1.7e-07 $l=6.44011e-07 $layer=licon1_PDIFF $count=2 $X=1.475
+ $Y=2.065 $X2=2 $Y2=2.33
r59 1 9 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%X 1 2 9 10 12 13 14 15
r18 14 15 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=2.502 $Y=1.835
+ $X2=2.502 $Y2=2.21
r19 11 13 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=2.535 $Y=0.655
+ $X2=2.535 $Y2=0.51
r20 11 12 6.62856 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.535 $Y=0.655
+ $X2=2.535 $Y2=0.775
r21 10 12 51.0182 $w=1.73e-07 $l=8.05e-07 $layer=LI1_cond $X=2.567 $Y=1.58
+ $X2=2.567 $Y2=0.775
r22 9 14 3.89186 $w=3.03e-07 $l=1.03e-07 $layer=LI1_cond $X=2.502 $Y=1.732
+ $X2=2.502 $Y2=1.835
r23 9 10 7.81944 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=2.502 $Y=1.732
+ $X2=2.502 $Y2=1.58
r24 2 14 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.485 $X2=2.5 $Y2=1.835
r25 1 13 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=2.5 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__AND2B_1%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r38 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r39 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r40 25 34 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.047
+ $Y2=0
r41 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.53
+ $Y2=0
r42 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r43 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r44 21 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r45 20 23 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r46 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 18 31 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r48 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r49 17 34 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.047
+ $Y2=0
r50 17 23 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.61
+ $Y2=0
r51 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r52 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r53 11 34 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=0.085
+ $X2=2.047 $Y2=0
r54 11 13 11.2327 $w=3.93e-07 $l=3.85e-07 $layer=LI1_cond $X=2.047 $Y=0.085
+ $X2=2.047 $Y2=0.47
r55 7 31 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r56 7 9 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.445
r57 2 13 182 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_NDIFF $count=1 $X=1.875
+ $Y=0.235 $X2=2.08 $Y2=0.47
r58 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends


* File: sky130_fd_sc_hd__a211oi_2.spice.pex
* Created: Thu Aug 27 13:59:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211OI_2%C1 1 3 6 8 10 13 15 16 21 24
c42 13 0 1.66419e-19 $X=0.955 $Y=1.985
r43 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.525 $Y=1.16
+ $X2=0.955 $Y2=1.16
r44 20 23 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.315 $Y=1.16
+ $X2=0.525 $Y2=1.16
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.16 $X2=0.315 $Y2=1.16
r46 15 16 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.252 $Y=1.19
+ $X2=0.252 $Y2=1.53
r47 15 21 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=0.252 $Y=1.19
+ $X2=0.252 $Y2=1.16
r48 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r50 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r52 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.985
r54 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%B1 1 3 6 8 10 13 15 16 17 26 28
r53 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.6 $Y=1.16
+ $X2=1.815 $Y2=1.16
r54 21 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.6 $Y2=1.16
r55 17 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.59 $Y=1.16
+ $X2=1.255 $Y2=1.16
r56 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r57 16 28 12.834 $w=2.18e-07 $l=2.45e-07 $layer=LI1_cond $X=1.145 $Y=1.53
+ $X2=1.145 $Y2=1.285
r58 15 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.145 $Y=1.16
+ $X2=1.145 $Y2=1.285
r59 15 32 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.145 $Y=1.16
+ $X2=1.255 $Y2=1.16
r60 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.16
r61 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.815 $Y=1.325
+ $X2=1.815 $Y2=1.985
r62 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=1.16
r63 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.815 $Y=0.995
+ $X2=1.815 $Y2=0.56
r64 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.16
r65 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.985
r66 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=0.995
+ $X2=1.385 $Y2=1.16
r67 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.385 $Y=0.995
+ $X2=1.385 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%A1 1 3 6 8 10 13 15 16 24
r41 22 24 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.895 $Y=1.16
+ $X2=3.195 $Y2=1.16
r42 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.895
+ $Y=1.16 $X2=2.895 $Y2=1.16
r43 19 22 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.765 $Y=1.16
+ $X2=2.895 $Y2=1.16
r44 16 23 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.99 $Y=1.16
+ $X2=2.895 $Y2=1.16
r45 15 23 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.895 $Y2=1.16
r46 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.16
r47 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.985
r48 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=0.995
+ $X2=3.195 $Y2=1.16
r49 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.195 $Y=0.995
+ $X2=3.195 $Y2=0.56
r50 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.325
+ $X2=2.765 $Y2=1.16
r51 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.765 $Y=1.325
+ $X2=2.765 $Y2=1.985
r52 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=0.995
+ $X2=2.765 $Y2=1.16
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.765 $Y=0.995
+ $X2=2.765 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%A2 1 3 6 8 10 13 15 16 17 28 31 35
c40 1 0 1.13948e-19 $X=3.625 $Y=0.995
r41 26 28 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.055 $Y=1.16
+ $X2=4.265 $Y2=1.16
r42 24 26 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=3.925 $Y=1.16
+ $X2=4.055 $Y2=1.16
r43 21 24 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=3.625 $Y=1.16
+ $X2=3.925 $Y2=1.16
r44 17 35 8.68765 $w=3.23e-07 $l=2.45e-07 $layer=LI1_cond $X=4.337 $Y=1.53
+ $X2=4.337 $Y2=1.285
r45 16 35 3.03503 $w=3.25e-07 $l=1.25e-07 $layer=LI1_cond $X=4.337 $Y=1.16
+ $X2=4.337 $Y2=1.285
r46 16 31 3.93339 $w=2.5e-07 $l=1.62e-07 $layer=LI1_cond $X=4.337 $Y=1.16
+ $X2=4.175 $Y2=1.16
r47 16 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=1.16 $X2=4.265 $Y2=1.16
r48 15 31 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3.91 $Y=1.16
+ $X2=4.175 $Y2=1.16
r49 15 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.16 $X2=3.925 $Y2=1.16
r50 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.055 $Y=1.325
+ $X2=4.055 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.055 $Y=1.325
+ $X2=4.055 $Y2=1.985
r52 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.055 $Y=0.995
+ $X2=4.055 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.055 $Y=0.995
+ $X2=4.055 $Y2=0.56
r54 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.625 $Y=1.325
+ $X2=3.625 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.625 $Y=1.325
+ $X2=3.625 $Y2=1.985
r56 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.625 $Y=0.995
+ $X2=3.625 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.625 $Y=0.995
+ $X2=3.625 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%A_37_297# 1 2 3 12 14 15 18 20 22 24 26
r35 22 28 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=2.075 $Y=2.255
+ $X2=2.075 $Y2=2.355
r36 22 24 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.075 $Y=2.255
+ $X2=2.075 $Y2=2
r37 21 26 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=1.265 $Y=2.355
+ $X2=1.17 $Y2=2.355
r38 20 28 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=1.935 $Y=2.355
+ $X2=2.075 $Y2=2.355
r39 20 21 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=1.935 $Y=2.355
+ $X2=1.265 $Y2=2.355
r40 16 26 1.24671 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=1.17 $Y=2.255 $X2=1.17
+ $Y2=2.355
r41 16 18 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.17 $Y=2.255
+ $X2=1.17 $Y2=1.95
r42 14 26 5.28167 $w=1.85e-07 $l=1.02225e-07 $layer=LI1_cond $X=1.075 $Y=2.37
+ $X2=1.17 $Y2=2.355
r43 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.075 $Y=2.37
+ $X2=0.405 $Y2=2.37
r44 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.275 $Y=2.285
+ $X2=0.405 $Y2=2.37
r45 10 12 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.275 $Y=2.285
+ $X2=0.275 $Y2=1.95
r46 3 28 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=2.34
r47 3 24 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.485 $X2=2.03 $Y2=2
r48 2 18 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.485 $X2=1.17 $Y2=1.95
r49 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%Y 1 2 3 4 13 17 20 21 22 23 24 25 26 37
c53 17 0 1.13948e-19 $X=2.98 $Y=0.755
r54 25 62 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.74 $Y=1.87 $X2=0.74
+ $Y2=1.99
r55 25 49 5.28534 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.715 $Y=1.785
+ $X2=0.715 $Y2=1.65
r56 24 49 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.715 $Y=1.53
+ $X2=0.715 $Y2=1.65
r57 23 24 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=0.715 $Y=1.19
+ $X2=0.715 $Y2=1.53
r58 22 35 3.99737 $w=2.7e-07 $l=1.04881e-07 $layer=LI1_cond $X=0.715 $Y=0.755
+ $X2=0.705 $Y2=0.655
r59 22 41 3.99737 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=0.715 $Y=0.755
+ $X2=0.715 $Y2=0.855
r60 22 23 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=0.895
+ $X2=0.715 $Y2=1.19
r61 22 41 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=0.715 $Y=0.895
+ $X2=0.715 $Y2=0.855
r62 21 35 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=0.705 $Y=0.51
+ $X2=0.705 $Y2=0.655
r63 21 37 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=0.705 $Y=0.51
+ $X2=0.705 $Y2=0.42
r64 19 26 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.6 $Y=0.655
+ $X2=1.6 $Y2=0.51
r65 19 20 1.5279 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=1.6 $Y=0.655 $X2=1.6
+ $Y2=0.755
r66 15 20 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.695 $Y=0.755 $X2=1.6
+ $Y2=0.755
r67 15 17 71.2591 $w=1.98e-07 $l=1.285e-06 $layer=LI1_cond $X=1.695 $Y=0.755
+ $X2=2.98 $Y2=0.755
r68 14 22 2.4424 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=0.855 $Y=0.755 $X2=0.715
+ $Y2=0.755
r69 13 20 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.505 $Y=0.755 $X2=1.6
+ $Y2=0.755
r70 13 14 36.0455 $w=1.98e-07 $l=6.5e-07 $layer=LI1_cond $X=1.505 $Y=0.755
+ $X2=0.855 $Y2=0.755
r71 4 62 600 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.74 $Y2=1.99
r72 4 49 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.74 $Y2=1.65
r73 3 17 182 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.235 $X2=2.98 $Y2=0.755
r74 2 26 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.235 $X2=1.6 $Y2=0.57
r75 1 22 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.76
r76 1 37 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%A_292_297# 1 2 3 12 16 18 20 22 25 27
c44 25 0 1.66419e-19 $X=1.6 $Y=1.65
r45 20 29 2.98511 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=3.84 $Y=1.655 $X2=3.84
+ $Y2=1.555
r46 20 22 27.5306 $w=2.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.84 $Y=1.655
+ $X2=3.84 $Y2=2.3
r47 19 27 6.58019 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=3.115 $Y=1.555
+ $X2=2.98 $Y2=1.555
r48 18 29 4.0299 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=3.705 $Y=1.555 $X2=3.84
+ $Y2=1.555
r49 18 19 32.7182 $w=1.98e-07 $l=5.9e-07 $layer=LI1_cond $X=3.705 $Y=1.555
+ $X2=3.115 $Y2=1.555
r50 14 27 0.287739 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=2.98 $Y=1.655 $X2=2.98
+ $Y2=1.555
r51 14 16 27.5306 $w=2.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.98 $Y=1.655
+ $X2=2.98 $Y2=2.3
r52 13 25 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=1.555 $X2=1.6
+ $Y2=1.555
r53 12 27 6.58019 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=2.845 $Y=1.555
+ $X2=2.98 $Y2=1.555
r54 12 13 59.8909 $w=1.98e-07 $l=1.08e-06 $layer=LI1_cond $X=2.845 $Y=1.555
+ $X2=1.765 $Y2=1.555
r55 3 29 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.485 $X2=3.84 $Y2=1.62
r56 3 22 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.485 $X2=3.84 $Y2=2.3
r57 2 27 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.485 $X2=2.98 $Y2=1.62
r58 2 16 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.485 $X2=2.98 $Y2=2.3
r59 1 25 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=1.46
+ $Y=1.485 $X2=1.6 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%VPWR 1 2 3 12 16 18 20 23 24 25 27 39 44 48
+ 52
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r64 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r65 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 39 47 3.76321 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.377 $Y2=2.72
r67 39 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 38 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r70 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 35 44 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.55 $Y2=2.72
r72 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.665 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 34 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 34 52 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=0.23 $Y2=2.72
r75 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 29 33 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 29 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 27 44 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.55 $Y2=2.72
r79 27 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.435 $Y=2.72
+ $X2=2.07 $Y2=2.72
r80 25 52 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 23 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 23 24 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.41 $Y2=2.72
r83 22 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.525 $Y=2.72
+ $X2=3.91 $Y2=2.72
r84 22 24 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.525 $Y=2.72
+ $X2=3.41 $Y2=2.72
r85 18 47 3.25467 $w=2.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=4.27 $Y=2.635
+ $X2=4.377 $Y2=2.72
r86 18 20 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.27 $Y=2.635
+ $X2=4.27 $Y2=2
r87 14 24 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=2.635
+ $X2=3.41 $Y2=2.72
r88 14 16 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.41 $Y=2.635
+ $X2=3.41 $Y2=2
r89 10 44 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=2.635
+ $X2=2.55 $Y2=2.72
r90 10 12 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.55 $Y=2.635
+ $X2=2.55 $Y2=2
r91 3 20 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=4.13
+ $Y=1.485 $X2=4.27 $Y2=2
r92 2 16 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=1.485 $X2=3.41 $Y2=2
r93 1 12 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.425
+ $Y=1.485 $X2=2.55 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%VGND 1 2 3 4 13 15 19 23 27 29 31 36 41 51
+ 52 58 61 64 69
r73 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r74 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r75 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r76 55 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 52 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r78 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r79 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.84
+ $Y2=0
r80 49 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.37
+ $Y2=0
r81 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r82 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r83 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r84 45 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r85 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r86 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r87 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.03
+ $Y2=0
r88 42 44 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.53
+ $Y2=0
r89 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.84
+ $Y2=0
r90 41 47 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.45
+ $Y2=0
r91 40 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r92 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r93 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r94 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.17
+ $Y2=0
r95 37 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.61
+ $Y2=0
r96 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.03
+ $Y2=0
r97 36 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.61
+ $Y2=0
r98 35 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r99 35 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r100 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r101 32 55 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r102 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r103 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.17
+ $Y2=0
r104 31 34 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=0.69 $Y2=0
r105 29 69 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r106 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0
r107 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0.36
r108 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r109 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.38
r110 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r111 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.38
r112 13 55 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r113 13 15 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.59
r114 4 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.7
+ $Y=0.235 $X2=3.84 $Y2=0.36
r115 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.235 $X2=2.03 $Y2=0.38
r116 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.38
r117 1 15 182 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__A211OI_2%A_485_47# 1 2 3 10 18 19 20
r28 20 22 4.148 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=0.635 $X2=4.31
+ $Y2=0.55
r29 18 20 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=4.185 $Y=0.745
+ $X2=4.31 $Y2=0.635
r30 18 19 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=4.185 $Y=0.745
+ $X2=3.495 $Y2=0.745
r31 15 19 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.41 $Y=0.635
+ $X2=3.495 $Y2=0.745
r32 15 17 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.41 $Y=0.635 $X2=3.41
+ $Y2=0.535
r33 14 17 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.41 $Y=0.475 $X2=3.41
+ $Y2=0.535
r34 10 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.325 $Y=0.37
+ $X2=3.41 $Y2=0.475
r35 10 12 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=3.325 $Y=0.37
+ $X2=2.55 $Y2=0.37
r36 3 22 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.235 $X2=4.27 $Y2=0.55
r37 2 17 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.235 $X2=3.41 $Y2=0.535
r38 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.55 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__sdfrbp_2.pex.spice
* Created: Thu Aug 27 14:45:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%CLK 1 3 6 8 9 15
c31 8 0 1.72041e-20 $X=0.215 $Y=1.19
c32 6 0 9.25139e-20 $X=0.47 $Y=1.985
r33 13 15 31.2282 $w=3.55e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.162
+ $X2=0.47 $Y2=1.162
r34 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.16 $X2=0.315
+ $Y2=1.53
r35 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r36 4 15 22.9692 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.47 $Y=1.345
+ $X2=0.47 $Y2=1.162
r37 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.47 $Y=1.345 $X2=0.47
+ $Y2=1.985
r38 1 15 22.9692 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.47 $Y=0.98
+ $X2=0.47 $Y2=1.162
r39 1 3 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=0.98 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_27_47# 1 2 7 9 12 16 18 20 23 25 27 31 35
+ 41 43 44 45 50 52 53 54 55 56 63 65 69 70 73 75 80 88
c263 80 0 1.04182e-19 $X=8.49 $Y=1.11
c264 70 0 1.18829e-19 $X=0.89 $Y=1.16
c265 69 0 1.34476e-19 $X=0.89 $Y=1.16
c266 54 0 1.14825e-19 $X=1.035 $Y=1.19
c267 50 0 9.88712e-20 $X=0.762 $Y=1.795
c268 45 0 7.54351e-20 $X=0.66 $Y=1.88
c269 35 0 1.24571e-19 $X=5.36 $Y=0.745
c270 27 0 6.68425e-20 $X=8.285 $Y=2.275
c271 16 0 1.63397e-19 $X=5.805 $Y=1.32
c272 7 0 1.72041e-20 $X=0.89 $Y=0.995
r273 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.49
+ $Y=1.11 $X2=8.49 $Y2=1.11
r274 73 76 16.4869 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=4.987 $Y=1.23
+ $X2=4.987 $Y2=1.32
r275 73 75 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=4.987 $Y=1.23
+ $X2=4.987 $Y2=1.065
r276 70 89 7.44021 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.817 $Y=1.16
+ $X2=0.817 $Y2=1.325
r277 70 88 8.29536 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.817 $Y=1.16
+ $X2=0.817 $Y2=0.995
r278 69 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.89 $Y2=1.325
r279 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.89
+ $Y=1.16 $X2=0.89 $Y2=1.16
r280 65 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.49 $Y=1.19
+ $X2=8.49 $Y2=1.19
r281 63 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.23 $X2=4.99 $Y2=1.23
r282 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.99 $Y=1.19
+ $X2=4.99 $Y2=1.19
r283 58 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.89 $Y=1.19
+ $X2=0.89 $Y2=1.19
r284 56 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.135 $Y=1.19
+ $X2=4.99 $Y2=1.19
r285 55 65 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.345 $Y=1.19
+ $X2=8.49 $Y2=1.19
r286 55 56 3.97276 $w=1.4e-07 $l=3.21e-06 $layer=MET1_cond $X=8.345 $Y=1.19
+ $X2=5.135 $Y2=1.19
r287 54 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.035 $Y=1.19
+ $X2=0.89 $Y2=1.19
r288 53 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.845 $Y=1.19
+ $X2=4.99 $Y2=1.19
r289 53 54 4.71534 $w=1.4e-07 $l=3.81e-06 $layer=MET1_cond $X=4.845 $Y=1.19
+ $X2=1.035 $Y2=1.19
r290 50 89 25.4279 $w=2.03e-07 $l=4.7e-07 $layer=LI1_cond $X=0.762 $Y=1.795
+ $X2=0.762 $Y2=1.325
r291 47 88 12.0416 $w=1.73e-07 $l=1.9e-07 $layer=LI1_cond $X=0.747 $Y=0.805
+ $X2=0.747 $Y2=0.995
r292 46 52 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.217 $Y2=1.88
r293 45 50 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.762 $Y2=1.795
r294 45 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r295 43 47 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.747 $Y2=0.805
r296 43 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r297 39 44 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.345 $Y2=0.72
r298 39 41 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.22 $Y=0.635
+ $X2=0.22 $Y2=0.51
r299 33 35 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.07 $Y=0.745
+ $X2=5.36 $Y2=0.745
r300 29 79 38.666 $w=2.85e-07 $l=1.71377e-07 $layer=POLY_cond $X=8.43 $Y=0.945
+ $X2=8.417 $Y2=1.11
r301 29 31 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.43 $Y=0.945
+ $X2=8.43 $Y2=0.415
r302 25 79 58.9607 $w=2.85e-07 $l=3.44739e-07 $layer=POLY_cond $X=8.285 $Y=1.395
+ $X2=8.417 $Y2=1.11
r303 25 27 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=8.285 $Y=1.395
+ $X2=8.285 $Y2=2.275
r304 21 23 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.88 $Y=1.395
+ $X2=5.88 $Y2=2.275
r305 18 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.36 $Y=0.67
+ $X2=5.36 $Y2=0.745
r306 18 20 81.94 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.36 $Y=0.67
+ $X2=5.36 $Y2=0.415
r307 17 76 20.1192 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=5.145 $Y=1.32
+ $X2=4.987 $Y2=1.32
r308 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.805 $Y=1.32
+ $X2=5.88 $Y2=1.395
r309 16 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.805 $Y=1.32
+ $X2=5.145 $Y2=1.32
r310 14 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.07 $Y=0.82
+ $X2=5.07 $Y2=0.745
r311 14 75 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.07 $Y=0.82
+ $X2=5.07 $Y2=1.065
r312 12 71 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.985
+ $X2=0.905 $Y2=1.325
r313 7 69 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r314 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r315 2 52 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r316 1 41 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_299_66# 1 2 7 9 10 12 16 18 19 20 22 25
+ 26 27 30 34 35 41
c137 26 0 1.05347e-19 $X=3.68 $Y=0.34
c138 12 0 1.99718e-19 $X=3.825 $Y=2.215
c139 10 0 1.99654e-19 $X=3.825 $Y=1.685
r140 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.29 $X2=2.385 $Y2=1.29
r141 38 40 7.07246 $w=3.45e-07 $l=2e-07 $layer=LI1_cond $X=2.225 $Y=1.09
+ $X2=2.225 $Y2=1.29
r142 34 35 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.22
+ $X2=2.025 $Y2=2.055
r143 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.765
+ $Y=1.52 $X2=3.765 $Y2=1.52
r144 28 30 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=3.765 $Y=0.425
+ $X2=3.765 $Y2=1.52
r145 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.68 $Y=0.34
+ $X2=3.765 $Y2=0.425
r146 26 27 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.68 $Y=0.34
+ $X2=3.085 $Y2=0.34
r147 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3 $Y=0.425
+ $X2=3.085 $Y2=0.34
r148 24 25 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3 $Y=0.425 $X2=3
+ $Y2=0.995
r149 23 38 4.22896 $w=1.9e-07 $l=2.45e-07 $layer=LI1_cond $X=2.47 $Y=1.09
+ $X2=2.225 $Y2=1.09
r150 22 25 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.915 $Y=1.09
+ $X2=3 $Y2=0.995
r151 22 23 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=2.915 $Y=1.09
+ $X2=2.47 $Y2=1.09
r152 20 40 8.97647 $w=3.45e-07 $l=2.31571e-07 $layer=LI1_cond $X=2.065 $Y=1.455
+ $X2=2.225 $Y2=1.29
r153 20 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.065 $Y=1.455
+ $X2=2.065 $Y2=2.055
r154 18 38 9.72464 $w=3.45e-07 $l=2.75e-07 $layer=LI1_cond $X=2.225 $Y=0.815
+ $X2=2.225 $Y2=1.09
r155 18 19 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.055 $Y=0.815
+ $X2=1.705 $Y2=0.815
r156 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=0.73
+ $X2=1.705 $Y2=0.815
r157 14 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.62 $Y=0.73
+ $X2=1.62 $Y2=0.56
r158 10 31 38.9235 $w=2.69e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.825 $Y=1.685
+ $X2=3.765 $Y2=1.52
r159 10 12 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.825 $Y=1.685
+ $X2=3.825 $Y2=2.215
r160 7 41 75.1296 $w=2.47e-07 $l=4.60999e-07 $layer=POLY_cond $X=2.77 $Y=1.09
+ $X2=2.385 $Y2=1.257
r161 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.77 $Y=1.09 $X2=2.77
+ $Y2=0.805
r162 2 34 600 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.945 $X2=1.985 $Y2=2.22
r163 1 16 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.33 $X2=1.62 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%D 3 7 9 10 14
c46 14 0 1.99654e-19 $X=3.035 $Y=1.62
c47 10 0 1.99718e-19 $X=2.925 $Y=2.125
r48 15 25 6.2547 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.927 $Y=1.62
+ $X2=2.927 $Y2=1.785
r49 14 17 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.62
+ $X2=3.052 $Y2=1.785
r50 14 16 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=3.052 $Y=1.62
+ $X2=3.052 $Y2=1.455
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.62 $X2=3.035 $Y2=1.62
r52 10 25 19.2074 $w=2.53e-07 $l=4.25e-07 $layer=LI1_cond $X=2.992 $Y=2.21
+ $X2=2.992 $Y2=1.785
r53 9 15 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=2.927 $Y=1.53 $X2=2.927
+ $Y2=1.62
r54 7 16 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.13 $Y=0.805
+ $X2=3.13 $Y2=1.455
r55 3 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.025 $Y=2.215
+ $X2=3.025 $Y2=1.785
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%SCE 4 5 6 7 11 13 17 19 21 22 24 26 27 31
+ 32
c99 32 0 4.13626e-20 $X=1.645 $Y=1.31
c100 31 0 2.66381e-19 $X=1.645 $Y=1.31
c101 19 0 1.79332e-19 $X=3.835 $Y=0.255
r102 31 33 43.918 $w=4.39e-07 $l=4e-07 $layer=POLY_cond $X=1.652 $Y=1.31
+ $X2=1.652 $Y2=1.71
r103 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.31 $X2=1.645 $Y2=1.31
r104 26 32 10.3485 $w=2.43e-07 $l=2.2e-07 $layer=LI1_cond $X=1.607 $Y=1.53
+ $X2=1.607 $Y2=1.31
r105 25 26 21.4025 $w=2.43e-07 $l=4.55e-07 $layer=LI1_cond $X=1.607 $Y=1.985
+ $X2=1.607 $Y2=1.53
r106 24 27 4.04442 $w=2.63e-07 $l=9.3e-08 $layer=LI1_cond $X=1.597 $Y=2.117
+ $X2=1.597 $Y2=2.21
r107 24 25 5.82496 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=1.597 $Y=2.117
+ $X2=1.597 $Y2=1.985
r108 19 21 27.474 $w=5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.835 $Y=0.255
+ $X2=3.835 $Y2=0.54
r109 15 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.615 $Y=1.785
+ $X2=2.615 $Y2=2.215
r110 14 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.71
+ $X2=2.195 $Y2=1.71
r111 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.54 $Y=1.71
+ $X2=2.615 $Y2=1.785
r112 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.54 $Y=1.71
+ $X2=2.27 $Y2=1.71
r113 9 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.785
+ $X2=2.195 $Y2=1.71
r114 9 11 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.785
+ $X2=2.195 $Y2=2.215
r115 8 33 28.1521 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=1.905 $Y=1.71
+ $X2=1.652 $Y2=1.71
r116 7 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.71
+ $X2=2.195 $Y2=1.71
r117 7 8 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.12 $Y=1.71
+ $X2=1.905 $Y2=1.71
r118 5 19 38.6381 $w=1.5e-07 $l=2.85044e-07 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.835 $Y2=0.255
r119 5 6 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=1.905 $Y2=0.18
r120 2 31 40.4229 $w=4.39e-07 $l=2.47091e-07 $layer=POLY_cond $X=1.83 $Y=1.145
+ $X2=1.652 $Y2=1.31
r121 2 4 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=1.83 $Y=1.145
+ $X2=1.83 $Y2=0.54
r122 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.83 $Y=0.255
+ $X2=1.905 $Y2=0.18
r123 1 4 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.255
+ $X2=1.83 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%SCD 3 7 13 16
c44 13 0 4.16547e-19 $X=4.165 $Y=1.53
c45 7 0 1.05347e-19 $X=4.385 $Y=0.54
r46 16 19 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.535
+ $X2=4.325 $Y2=1.7
r47 16 18 42.5162 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.535
+ $X2=4.325 $Y2=1.37
r48 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.31
+ $Y=1.535 $X2=4.31 $Y2=1.535
r49 13 17 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=4.207 $Y=1.53
+ $X2=4.207 $Y2=1.535
r50 7 18 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=4.385 $Y=0.54
+ $X2=4.385 $Y2=1.37
r51 3 19 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.255 $Y=2.215
+ $X2=4.255 $Y2=1.7
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_193_47# 1 2 9 13 14 16 19 23 26 29 31 32
+ 36 37 39 40 44 46 51 54 55 56 57 58 67 71 72 76 88 91
c270 88 0 1.95569e-19 $X=1.23 $Y=1.815
c271 76 0 1.25175e-19 $X=5.8 $Y=0.705
c272 71 0 1.38309e-19 $X=5.33 $Y=1.74
c273 56 0 9.25139e-20 $X=1.27 $Y=1.87
c274 55 0 3.51014e-19 $X=5.265 $Y=1.87
c275 54 0 6.24992e-20 $X=8.705 $Y=1.74
c276 51 0 8.14383e-20 $X=8.69 $Y=1.805
c277 46 0 8.4081e-20 $X=8.415 $Y=1.58
c278 36 0 1.25072e-19 $X=8.01 $Y=0.87
c279 32 0 4.31332e-21 $X=5.8 $Y=0.87
r280 72 91 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.74
+ $X2=5.37 $Y2=1.575
r281 71 74 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.33 $Y=1.74
+ $X2=5.33 $Y2=1.875
r282 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.33
+ $Y=1.74 $X2=5.33 $Y2=1.74
r283 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.53 $Y=1.87
+ $X2=8.53 $Y2=1.87
r284 64 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.41 $Y=1.87
+ $X2=5.41 $Y2=1.87
r285 61 88 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.12 $Y=1.815
+ $X2=1.23 $Y2=1.815
r286 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.12 $Y=1.87
+ $X2=1.12 $Y2=1.87
r287 58 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.555 $Y=1.87
+ $X2=5.41 $Y2=1.87
r288 57 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.385 $Y=1.87
+ $X2=8.53 $Y2=1.87
r289 57 58 3.50247 $w=1.4e-07 $l=2.83e-06 $layer=MET1_cond $X=8.385 $Y=1.87
+ $X2=5.555 $Y2=1.87
r290 56 60 0.118675 $w=2.3e-07 $l=1.5e-07 $layer=MET1_cond $X=1.27 $Y=1.87
+ $X2=1.12 $Y2=1.87
r291 55 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.265 $Y=1.87
+ $X2=5.41 $Y2=1.87
r292 55 56 4.9443 $w=1.4e-07 $l=3.995e-06 $layer=MET1_cond $X=5.265 $Y=1.87
+ $X2=1.27 $Y2=1.87
r293 54 84 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.705 $Y=1.74
+ $X2=8.705 $Y2=1.905
r294 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=1.74 $X2=8.705 $Y2=1.74
r295 51 68 6.14636 $w=2.98e-07 $l=1.6e-07 $layer=LI1_cond $X=8.69 $Y=1.805
+ $X2=8.53 $Y2=1.805
r296 51 53 0.61 $w=3e-07 $l=1.5e-08 $layer=LI1_cond $X=8.69 $Y=1.805 $X2=8.705
+ $Y2=1.805
r297 49 68 0.384148 $w=2.98e-07 $l=1e-08 $layer=LI1_cond $X=8.52 $Y=1.805
+ $X2=8.53 $Y2=1.805
r298 46 49 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=8.415 $Y=1.58
+ $X2=8.415 $Y2=1.805
r299 42 44 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.23 $Y2=0.51
r300 39 46 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.31 $Y=1.58
+ $X2=8.415 $Y2=1.58
r301 39 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.31 $Y=1.58
+ $X2=8.095 $Y2=1.58
r302 37 78 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=8.01 $Y=0.87
+ $X2=7.885 $Y2=0.87
r303 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.01
+ $Y=0.87 $X2=8.01 $Y2=0.87
r304 34 40 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.99 $Y=1.495
+ $X2=8.095 $Y2=1.58
r305 34 36 33.0087 $w=2.08e-07 $l=6.25e-07 $layer=LI1_cond $X=7.99 $Y=1.495
+ $X2=7.99 $Y2=0.87
r306 32 76 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=0.87
+ $X2=5.8 $Y2=0.705
r307 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.8
+ $Y=0.87 $X2=5.8 $Y2=0.87
r308 29 31 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.495 $Y=0.87
+ $X2=5.8 $Y2=0.87
r309 27 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.41 $Y=1.035
+ $X2=5.495 $Y2=0.87
r310 27 91 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.41 $Y=1.035
+ $X2=5.41 $Y2=1.575
r311 26 88 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=1.73
+ $X2=1.23 $Y2=1.815
r312 25 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0.675
+ $X2=1.23 $Y2=0.51
r313 25 26 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=1.23 $Y=0.675
+ $X2=1.23 $Y2=1.73
r314 21 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.9
+ $X2=1.12 $Y2=1.815
r315 21 23 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.12 $Y=1.9 $X2=1.12
+ $Y2=1.96
r316 19 84 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.715 $Y=2.275
+ $X2=8.715 $Y2=1.905
r317 14 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.885 $Y=0.705
+ $X2=7.885 $Y2=0.87
r318 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.885 $Y=0.705
+ $X2=7.885 $Y2=0.415
r319 13 76 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.86 $Y=0.415
+ $X2=5.86 $Y2=0.705
r320 9 74 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.32 $Y=2.275 $X2=5.32
+ $Y2=1.875
r321 2 23 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=1.96
r322 1 42 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_1245_303# 1 2 9 13 15 18 21 24 28 31 34
+ 35 36
c112 36 0 6.68425e-20 $X=7.585 $Y=1.595
c113 34 0 1.40308e-19 $X=7.585 $Y=0.835
c114 1 0 1.64006e-19 $X=7.485 $Y=0.235
r115 35 37 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=7.585 $Y=1.68
+ $X2=7.585 $Y2=1.92
r116 35 36 5.14764 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=7.585 $Y=1.68
+ $X2=7.585 $Y2=1.595
r117 34 36 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.63 $Y=0.835
+ $X2=7.63 $Y2=1.595
r118 31 33 3.51899 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=0.36
+ $X2=7.62 $Y2=0.445
r119 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.055 $Y=2.005
+ $X2=8.055 $Y2=2.3
r120 25 37 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.715 $Y=1.92
+ $X2=7.585 $Y2=1.92
r121 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.97 $Y=1.92
+ $X2=8.055 $Y2=2.005
r122 24 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.97 $Y=1.92
+ $X2=7.715 $Y2=1.92
r123 21 34 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=7.585 $Y=0.705
+ $X2=7.585 $Y2=0.835
r124 21 33 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=7.585 $Y=0.705
+ $X2=7.585 $Y2=0.445
r125 18 41 48.1856 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=6.405 $Y=1.68
+ $X2=6.405 $Y2=1.855
r126 18 40 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=6.405 $Y=1.68
+ $X2=6.405 $Y2=1.515
r127 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.68 $X2=6.45 $Y2=1.68
r128 15 35 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.455 $Y=1.68
+ $X2=7.585 $Y2=1.68
r129 15 17 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=7.455 $Y=1.68
+ $X2=6.45 $Y2=1.68
r130 13 40 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=6.39 $Y=0.445
+ $X2=6.39 $Y2=1.515
r131 9 41 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=6.3 $Y=2.275 $X2=6.3
+ $Y2=1.855
r132 2 28 600 $w=1.7e-07 $l=7.35102e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.645 $X2=8.055 $Y2=2.3
r133 1 31 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=7.485
+ $Y=0.235 $X2=7.62 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%RESET_B 3 6 8 9 12 14 16 17 19 20 24 27 29
+ 30 31 38 40 48
c169 48 0 1.42544e-19 $X=9.97 $Y=1.065
c170 38 0 1.40308e-19 $X=6.81 $Y=0.96
c171 31 0 1.38838e-19 $X=9.775 $Y=0.965
c172 29 0 1.64006e-19 $X=9.63 $Y=0.85
c173 20 0 2.28755e-20 $X=10.03 $Y=0.85
c174 12 0 4.33854e-20 $X=9.655 $Y=0.445
c175 6 0 1.1086e-19 $X=6.87 $Y=2.275
r176 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=1.15 $X2=9.69 $Y2=1.15
r177 38 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=0.96
+ $X2=6.81 $Y2=1.125
r178 38 40 57.3029 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=6.81 $Y=0.96
+ $X2=6.81 $Y2=0.755
r179 31 35 0.153245 $w=2.08e-07 $l=2.55e-07 $layer=MET1_cond $X=9.775 $Y=0.85
+ $X2=10.03 $Y2=0.85
r180 29 31 0.100553 $w=2.08e-07 $l=1.45e-07 $layer=MET1_cond $X=9.63 $Y=0.85
+ $X2=9.775 $Y2=0.85
r181 29 30 3.13737 $w=1.4e-07 $l=2.535e-06 $layer=MET1_cond $X=9.63 $Y=0.85
+ $X2=7.095 $Y2=0.85
r182 27 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.81
+ $Y=0.96 $X2=6.81 $Y2=0.96
r183 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.95 $Y=0.85
+ $X2=6.95 $Y2=0.85
r184 24 30 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=6.98 $Y=0.85
+ $X2=7.095 $Y2=0.85
r185 24 26 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=6.98 $Y=0.85
+ $X2=6.95 $Y2=0.85
r186 20 48 8.54397 $w=2.88e-07 $l=2.15e-07 $layer=LI1_cond $X=9.97 $Y=0.85
+ $X2=9.97 $Y2=1.065
r187 20 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.03 $Y=0.85
+ $X2=10.03 $Y2=0.85
r188 19 48 2.95929 $w=2.9e-07 $l=1.05e-07 $layer=LI1_cond $X=9.97 $Y=1.17
+ $X2=9.97 $Y2=1.065
r189 19 44 6.38319 $w=3.78e-07 $l=1.35e-07 $layer=LI1_cond $X=9.825 $Y=1.17
+ $X2=9.69 $Y2=1.17
r190 17 18 59.8102 $w=1.37e-07 $l=1.7e-07 $layer=POLY_cond $X=9.485 $Y=1.915
+ $X2=9.655 $Y2=1.915
r191 14 18 0.6158 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.655 $Y=1.99
+ $X2=9.655 $Y2=1.915
r192 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.655 $Y=1.99
+ $X2=9.655 $Y2=2.275
r193 10 43 38.8259 $w=2.74e-07 $l=1.83016e-07 $layer=POLY_cond $X=9.655 $Y=0.985
+ $X2=9.617 $Y2=1.15
r194 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.655 $Y=0.985
+ $X2=9.655 $Y2=0.445
r195 9 17 0.6158 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.485 $Y=1.84
+ $X2=9.485 $Y2=1.915
r196 8 43 59.9354 $w=2.74e-07 $l=3.44739e-07 $layer=POLY_cond $X=9.485 $Y=1.435
+ $X2=9.617 $Y2=1.15
r197 8 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.485 $Y=1.435
+ $X2=9.485 $Y2=1.84
r198 6 41 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=6.87 $Y=2.275
+ $X2=6.87 $Y2=1.125
r199 3 40 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.75 $Y=0.445
+ $X2=6.75 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_1079_413# 1 2 9 11 13 15 16 22 23 25 26
+ 29 30 32 34 35
c139 34 0 1.1086e-19 $X=7.29 $Y=1.17
c140 32 0 1.87801e-19 $X=6.25 $Y=1.3
c141 29 0 1.38309e-19 $X=5.67 $Y=2.33
c142 11 0 8.4081e-20 $X=7.735 $Y=1.495
c143 9 0 1.25072e-19 $X=7.41 $Y=0.555
r144 34 37 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.29 $Y=1.17
+ $X2=7.29 $Y2=1.3
r145 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.29
+ $Y=1.17 $X2=7.29 $Y2=1.17
r146 29 30 9.47152 $w=3.63e-07 $l=1.95e-07 $layer=LI1_cond $X=5.652 $Y=2.33
+ $X2=5.652 $Y2=2.135
r147 27 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=1.3
+ $X2=6.25 $Y2=1.3
r148 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.205 $Y=1.3
+ $X2=7.29 $Y2=1.3
r149 26 27 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.205 $Y=1.3
+ $X2=6.335 $Y2=1.3
r150 25 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=1.215
+ $X2=6.25 $Y2=1.3
r151 24 25 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.25 $Y=0.475
+ $X2=6.25 $Y2=1.215
r152 22 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=1.3
+ $X2=6.25 $Y2=1.3
r153 22 23 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.165 $Y=1.3
+ $X2=5.835 $Y2=1.3
r154 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.75 $Y=1.385
+ $X2=5.835 $Y2=1.3
r155 20 30 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.75 $Y=1.385
+ $X2=5.75 $Y2=2.135
r156 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.165 $Y=0.39
+ $X2=6.25 $Y2=0.475
r157 16 18 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.165 $Y=0.39
+ $X2=5.65 $Y2=0.39
r158 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.81 $Y=1.57
+ $X2=7.81 $Y2=2.065
r159 12 35 61.4314 $w=2.55e-07 $l=3.99061e-07 $layer=POLY_cond $X=7.485 $Y=1.495
+ $X2=7.32 $Y2=1.17
r160 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.735 $Y=1.495
+ $X2=7.81 $Y2=1.57
r161 11 12 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=7.735 $Y=1.495
+ $X2=7.485 $Y2=1.495
r162 7 35 39.2931 $w=2.55e-07 $l=2.05122e-07 $layer=POLY_cond $X=7.41 $Y=1.005
+ $X2=7.32 $Y2=1.17
r163 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=7.41 $Y=1.005
+ $X2=7.41 $Y2=0.555
r164 2 29 600 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=2.065 $X2=5.67 $Y2=2.33
r165 1 18 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.235 $X2=5.65 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_1767_21# 1 2 9 13 17 21 23 25 28 30 32 35
+ 39 42 43 45 46 47 52 54 55 57 59 62 65 67 74
c188 74 0 2.27161e-19 $X=11.95 $Y=1.16
c189 67 0 2.28902e-19 $X=9.125 $Y=0.98
c190 42 0 1.85044e-19 $X=9.485 $Y=0.78
c191 35 0 1.62009e-19 $X=11.95 $Y=1.985
c192 21 0 1.52702e-19 $X=11.015 $Y=2.125
c193 13 0 1.58056e-19 $X=9.125 $Y=2.275
r194 73 74 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=11.49 $Y=1.16
+ $X2=11.95 $Y2=1.16
r195 72 73 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=11.015 $Y=1.16
+ $X2=11.49 $Y2=1.16
r196 71 72 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=11.01 $Y=1.16
+ $X2=11.015 $Y2=1.16
r197 63 71 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=10.895 $Y=1.16
+ $X2=11.01 $Y2=1.16
r198 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.895
+ $Y=1.16 $X2=10.895 $Y2=1.16
r199 60 65 0.256868 $w=2.7e-07 $l=2.58844e-07 $layer=LI1_cond $X=10.545 $Y=1.19
+ $X2=10.345 $Y2=1.055
r200 60 62 14.9391 $w=2.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.545 $Y=1.19
+ $X2=10.895 $Y2=1.19
r201 58 65 7.44763 $w=1.7e-07 $l=3.22413e-07 $layer=LI1_cond $X=10.46 $Y=1.325
+ $X2=10.345 $Y2=1.055
r202 58 59 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.46 $Y=1.325
+ $X2=10.46 $Y2=1.915
r203 57 65 7.44763 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.43 $Y=1.055
+ $X2=10.345 $Y2=1.055
r204 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.43 $Y=0.465
+ $X2=10.43 $Y2=1.055
r205 54 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.375 $Y=2
+ $X2=10.46 $Y2=1.915
r206 54 55 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.375 $Y=2
+ $X2=9.95 $Y2=2
r207 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.865 $Y=2.085
+ $X2=9.95 $Y2=2
r208 50 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.865 $Y=2.085
+ $X2=9.865 $Y2=2.21
r209 47 49 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.655 $Y=0.38
+ $X2=10.26 $Y2=0.38
r210 46 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.345 $Y=0.38
+ $X2=10.43 $Y2=0.465
r211 46 49 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.38
+ $X2=10.26 $Y2=0.38
r212 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.57 $Y=0.465
+ $X2=9.655 $Y2=0.38
r213 44 45 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.57 $Y=0.465
+ $X2=9.57 $Y2=0.695
r214 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.485 $Y=0.78
+ $X2=9.57 $Y2=0.695
r215 42 43 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.485 $Y=0.78
+ $X2=9.295 $Y2=0.78
r216 40 67 16.1937 $w=2.53e-07 $l=8.5e-08 $layer=POLY_cond $X=9.21 $Y=0.98
+ $X2=9.125 $Y2=0.98
r217 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.21
+ $Y=0.98 $X2=9.21 $Y2=0.98
r218 37 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.21 $Y=0.865
+ $X2=9.295 $Y2=0.78
r219 37 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.21 $Y=0.865
+ $X2=9.21 $Y2=0.98
r220 33 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.95 $Y=1.325
+ $X2=11.95 $Y2=1.16
r221 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.95 $Y=1.325
+ $X2=11.95 $Y2=1.985
r222 30 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.95 $Y=0.995
+ $X2=11.95 $Y2=1.16
r223 30 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.95 $Y=0.995
+ $X2=11.95 $Y2=0.56
r224 26 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.49 $Y=1.325
+ $X2=11.49 $Y2=1.16
r225 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.49 $Y=1.325
+ $X2=11.49 $Y2=1.985
r226 23 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.49 $Y=0.995
+ $X2=11.49 $Y2=1.16
r227 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.49 $Y=0.995
+ $X2=11.49 $Y2=0.56
r228 19 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.015 $Y=1.325
+ $X2=11.015 $Y2=1.16
r229 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=11.015 $Y=1.325
+ $X2=11.015 $Y2=2.125
r230 15 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.01 $Y=0.995
+ $X2=11.01 $Y2=1.16
r231 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=11.01 $Y=0.995
+ $X2=11.01 $Y2=0.445
r232 11 67 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.145
+ $X2=9.125 $Y2=0.98
r233 11 13 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=9.125 $Y=1.145
+ $X2=9.125 $Y2=2.275
r234 7 67 40.9605 $w=2.53e-07 $l=2.85832e-07 $layer=POLY_cond $X=8.91 $Y=0.815
+ $X2=9.125 $Y2=0.98
r235 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.91 $Y=0.815
+ $X2=8.91 $Y2=0.445
r236 2 52 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.73
+ $Y=2.065 $X2=9.865 $Y2=2.21
r237 1 49 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=10.125
+ $Y=0.235 $X2=10.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_1592_47# 1 2 7 9 10 12 15 16 20 25 27 28
+ 30
c117 25 0 1.41552e-19 $X=8.83 $Y=1.315
c118 16 0 4.33854e-20 $X=8.745 $Y=0.395
c119 15 0 1.82308e-20 $X=10.11 $Y=1.495
c120 7 0 1.66814e-19 $X=10.05 $Y=0.73
r121 33 34 13.5811 $w=2.65e-07 $l=2.95e-07 $layer=LI1_cond $X=8.83 $Y=1.485
+ $X2=9.125 $Y2=1.485
r122 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.04
+ $Y=1.66 $X2=10.04 $Y2=1.66
r123 28 34 5.47642 $w=2.65e-07 $l=2.13307e-07 $layer=LI1_cond $X=9.21 $Y=1.66
+ $X2=9.125 $Y2=1.485
r124 28 30 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.21 $Y=1.66
+ $X2=10.04 $Y2=1.66
r125 26 34 3.33486 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=9.125 $Y=1.745
+ $X2=9.125 $Y2=1.485
r126 26 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.125 $Y=1.745
+ $X2=9.125 $Y2=2.035
r127 25 33 3.33486 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.83 $Y=1.315
+ $X2=8.83 $Y2=1.485
r128 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=8.83 $Y=0.535
+ $X2=8.83 $Y2=1.315
r129 20 27 3.88471 $w=5.15e-07 $l=3.10161e-07 $layer=LI1_cond $X=9.015 $Y=2.295
+ $X2=9.125 $Y2=2.035
r130 20 22 17.2866 $w=3.38e-07 $l=5.1e-07 $layer=LI1_cond $X=9.015 $Y=2.295
+ $X2=8.505 $Y2=2.295
r131 16 24 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=8.745 $Y=0.395
+ $X2=8.83 $Y2=0.535
r132 16 18 23.6662 $w=2.78e-07 $l=5.75e-07 $layer=LI1_cond $X=8.745 $Y=0.395
+ $X2=8.17 $Y2=0.395
r133 15 31 38.7444 $w=2.79e-07 $l=1.94808e-07 $layer=POLY_cond $X=10.11 $Y=1.495
+ $X2=10.045 $Y2=1.66
r134 14 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.11 $Y=0.85
+ $X2=10.11 $Y2=1.495
r135 10 31 38.7444 $w=2.79e-07 $l=1.79374e-07 $layer=POLY_cond $X=10.075
+ $Y=1.825 $X2=10.045 $Y2=1.66
r136 10 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.075 $Y=1.825
+ $X2=10.075 $Y2=2.275
r137 7 14 28.3529 $w=2.04e-07 $l=1.46969e-07 $layer=POLY_cond $X=10.05 $Y=0.73
+ $X2=10.11 $Y2=0.85
r138 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.05 $Y=0.73
+ $X2=10.05 $Y2=0.445
r139 2 22 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=8.36
+ $Y=2.065 $X2=8.505 $Y2=2.335
r140 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.96
+ $Y=0.235 $X2=8.17 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_2135_47# 1 2 7 9 12 14 16 19 23 27 28 29
+ 32 34 36 37 42 47
c110 47 0 1.91378e-19 $X=12.82 $Y=1.16
c111 37 0 1.52702e-19 $X=11.317 $Y=1.94
r112 43 47 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=12.4 $Y=1.16
+ $X2=12.82 $Y2=1.16
r113 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.4
+ $Y=1.16 $X2=12.4 $Y2=1.16
r114 39 42 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=12.18 $Y=1.16
+ $X2=12.4 $Y2=1.16
r115 34 37 48.7435 $w=2.16e-07 $l=8.63e-07 $layer=LI1_cond $X=12.18 $Y=1.94
+ $X2=11.317 $Y2=1.94
r116 33 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=1.325
+ $X2=12.18 $Y2=1.16
r117 33 34 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=12.18 $Y=1.325
+ $X2=12.18 $Y2=1.865
r118 32 37 2.00054 $w=1.75e-07 $l=1.45e-07 $layer=LI1_cond $X=11.317 $Y=1.795
+ $X2=11.317 $Y2=1.94
r119 31 32 57.6727 $w=1.73e-07 $l=9.1e-07 $layer=LI1_cond $X=11.317 $Y=0.885
+ $X2=11.317 $Y2=1.795
r120 30 36 2.97688 $w=2.4e-07 $l=8.8e-08 $layer=LI1_cond $X=10.89 $Y=1.915
+ $X2=10.802 $Y2=1.915
r121 29 37 4.57109 $w=2.4e-07 $l=9.87117e-08 $layer=LI1_cond $X=11.23 $Y=1.915
+ $X2=11.317 $Y2=1.94
r122 29 30 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=11.23 $Y=1.915
+ $X2=10.89 $Y2=1.915
r123 27 31 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=11.23 $Y=0.8
+ $X2=11.317 $Y2=0.885
r124 27 28 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.23 $Y=0.8
+ $X2=10.885 $Y2=0.8
r125 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.8 $Y=0.715
+ $X2=10.885 $Y2=0.8
r126 21 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.8 $Y=0.715
+ $X2=10.8 $Y2=0.51
r127 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.82 $Y=1.325
+ $X2=12.82 $Y2=1.16
r128 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.82 $Y=1.325
+ $X2=12.82 $Y2=1.985
r129 14 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.82 $Y=0.995
+ $X2=12.82 $Y2=1.16
r130 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.82 $Y=0.995
+ $X2=12.82 $Y2=0.56
r131 10 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.4 $Y=1.325
+ $X2=12.4 $Y2=1.16
r132 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.4 $Y=1.325
+ $X2=12.4 $Y2=1.985
r133 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.4 $Y=0.995
+ $X2=12.4 $Y2=1.16
r134 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.4 $Y=0.995
+ $X2=12.4 $Y2=0.56
r135 2 36 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=10.68
+ $Y=1.805 $X2=10.805 $Y2=1.96
r136 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=10.675
+ $Y=0.235 $X2=10.8 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 61 63 65 70 71 73 76 79 81 93 104 108 113 118 123 128 134 137 140 143 146
+ 149 152 156 159
c217 70 0 6.21315e-20 $X=2.32 $Y=2.72
r218 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r219 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r220 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r221 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r222 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r223 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r224 137 138 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r225 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r226 132 156 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r227 132 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r228 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r229 129 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.355 $Y=2.72
+ $X2=12.19 $Y2=2.72
r230 129 131 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.355 $Y=2.72
+ $X2=12.65 $Y2=2.72
r231 128 155 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.995 $Y=2.72
+ $X2=13.167 $Y2=2.72
r232 128 131 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.995 $Y=2.72
+ $X2=12.65 $Y2=2.72
r233 127 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r234 127 150 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r235 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r236 124 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.42 $Y=2.72
+ $X2=11.255 $Y2=2.72
r237 124 126 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.42 $Y=2.72
+ $X2=11.73 $Y2=2.72
r238 123 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=12.19 $Y2=2.72
r239 123 126 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=11.73 $Y2=2.72
r240 122 150 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r241 122 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r242 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r243 119 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=2.72
+ $X2=10.285 $Y2=2.72
r244 119 121 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=10.45 $Y=2.72
+ $X2=10.81 $Y2=2.72
r245 118 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.09 $Y=2.72
+ $X2=11.255 $Y2=2.72
r246 118 121 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.09 $Y=2.72
+ $X2=10.81 $Y2=2.72
r247 117 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r248 117 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r249 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r250 114 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.61 $Y=2.72
+ $X2=9.485 $Y2=2.72
r251 114 116 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=9.61 $Y=2.72
+ $X2=9.89 $Y2=2.72
r252 113 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.12 $Y=2.72
+ $X2=10.285 $Y2=2.72
r253 113 116 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=10.12 $Y=2.72
+ $X2=9.89 $Y2=2.72
r254 112 144 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=9.43 $Y2=2.72
r255 112 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r256 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r257 109 140 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.745 $Y=2.72
+ $X2=7.56 $Y2=2.72
r258 109 111 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=2.72
+ $X2=8.05 $Y2=2.72
r259 108 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=9.485 $Y2=2.72
r260 108 111 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=9.36 $Y=2.72
+ $X2=8.05 $Y2=2.72
r261 107 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r262 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r263 104 140 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=7.375 $Y=2.72
+ $X2=7.56 $Y2=2.72
r264 104 106 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.375 $Y=2.72
+ $X2=7.13 $Y2=2.72
r265 103 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r266 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r267 100 103 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r268 100 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r269 99 102 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r270 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r271 97 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=2.72
+ $X2=4.465 $Y2=2.72
r272 97 99 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.63 $Y=2.72 $X2=4.83
+ $Y2=2.72
r273 96 138 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.37 $Y2=2.72
r274 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r275 93 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=2.72
+ $X2=4.465 $Y2=2.72
r276 93 95 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=4.3 $Y=2.72
+ $X2=2.53 $Y2=2.72
r277 92 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r278 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r279 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r280 89 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r281 88 91 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r282 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r283 86 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=2.72
+ $X2=0.695 $Y2=2.72
r284 86 88 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=2.72
+ $X2=1.15 $Y2=2.72
r285 83 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r286 81 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=2.72
+ $X2=0.695 $Y2=2.72
r287 81 83 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.53 $Y=2.72 $X2=0.23
+ $Y2=2.72
r288 79 135 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r289 79 159 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r290 77 106 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.74 $Y=2.72
+ $X2=7.13 $Y2=2.72
r291 76 102 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.41 $Y=2.72
+ $X2=6.21 $Y2=2.72
r292 75 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.74 $Y2=2.72
r293 75 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.41 $Y2=2.72
r294 73 75 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.575 $Y=2.44
+ $X2=6.575 $Y2=2.72
r295 70 91 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.32 $Y=2.72
+ $X2=2.07 $Y2=2.72
r296 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.32 $Y=2.72
+ $X2=2.405 $Y2=2.72
r297 69 95 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.49 $Y=2.72 $X2=2.53
+ $Y2=2.72
r298 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=2.72
+ $X2=2.405 $Y2=2.72
r299 65 68 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=13.12 $Y=1.66
+ $X2=13.12 $Y2=2.34
r300 63 155 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=13.12 $Y=2.635
+ $X2=13.167 $Y2=2.72
r301 63 68 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.12 $Y=2.635
+ $X2=13.12 $Y2=2.34
r302 59 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.19 $Y=2.635
+ $X2=12.19 $Y2=2.72
r303 59 61 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.19 $Y=2.635
+ $X2=12.19 $Y2=2.34
r304 55 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.255 $Y=2.635
+ $X2=11.255 $Y2=2.72
r305 55 57 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=11.255 $Y=2.635
+ $X2=11.255 $Y2=2.29
r306 51 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=2.635
+ $X2=10.285 $Y2=2.72
r307 51 53 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.285 $Y=2.635
+ $X2=10.285 $Y2=2.34
r308 47 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.485 $Y=2.635
+ $X2=9.485 $Y2=2.72
r309 47 49 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=9.485 $Y=2.635
+ $X2=9.485 $Y2=2.36
r310 43 140 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.56 $Y=2.635
+ $X2=7.56 $Y2=2.72
r311 43 45 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.56 $Y=2.635
+ $X2=7.56 $Y2=2.34
r312 39 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=2.635
+ $X2=4.465 $Y2=2.72
r313 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.465 $Y=2.635
+ $X2=4.465 $Y2=2.36
r314 35 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=2.635
+ $X2=2.405 $Y2=2.72
r315 35 37 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.405 $Y=2.635
+ $X2=2.405 $Y2=2.225
r316 31 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.72
r317 31 33 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.695 $Y=2.635
+ $X2=0.695 $Y2=2.22
r318 10 68 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=12.895
+ $Y=1.485 $X2=13.08 $Y2=2.34
r319 10 65 400 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=1 $X=12.895
+ $Y=1.485 $X2=13.08 $Y2=1.66
r320 9 61 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=12.025
+ $Y=1.485 $X2=12.19 $Y2=2.34
r321 8 57 600 $w=1.7e-07 $l=5.61471e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.805 $X2=11.255 $Y2=2.29
r322 7 53 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.15
+ $Y=2.065 $X2=10.285 $Y2=2.34
r323 6 49 600 $w=1.7e-07 $l=3.99124e-07 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=2.065 $X2=9.445 $Y2=2.36
r324 5 45 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=7.475
+ $Y=1.645 $X2=7.6 $Y2=2.34
r325 4 73 600 $w=1.7e-07 $l=4.64354e-07 $layer=licon1_PDIFF $count=1 $X=6.375
+ $Y=2.065 $X2=6.575 $Y2=2.44
r326 3 41 600 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_PDIFF $count=1 $X=4.33
+ $Y=1.945 $X2=4.465 $Y2=2.36
r327 2 37 600 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.945 $X2=2.405 $Y2=2.225
r328 1 33 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.695 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_620_389# 1 2 3 4 15 18 21 23 24 26 27 28
+ 30 32 42
c103 32 0 1.87617e-19 $X=3.357 $Y=1.185
c104 30 0 2.63145e-19 $X=5.06 $Y=0.715
r105 39 42 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.06 $Y=0.42 $X2=5.15
+ $Y2=0.42
r106 33 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.375 $Y=2.02
+ $X2=3.545 $Y2=2.02
r107 31 32 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=3.357 $Y=1.015
+ $X2=3.357 $Y2=1.185
r108 29 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.505
+ $X2=5.06 $Y2=0.42
r109 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.06 $Y=0.505
+ $X2=5.06 $Y2=0.715
r110 27 30 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.975 $Y=0.805
+ $X2=5.06 $Y2=0.715
r111 27 28 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=4.975 $Y=0.805
+ $X2=4.735 $Y2=0.805
r112 26 38 20.7085 $w=2.71e-07 $l=5.71489e-07 $layer=LI1_cond $X=4.65 $Y=1.935
+ $X2=5.11 $Y2=2.185
r113 25 28 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.65 $Y=0.895
+ $X2=4.735 $Y2=0.805
r114 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.65 $Y=0.895
+ $X2=4.65 $Y2=1.935
r115 24 35 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=2.02
+ $X2=3.545 $Y2=2.02
r116 23 26 5.51241 $w=2.71e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.565 $Y=2.02
+ $X2=4.65 $Y2=1.935
r117 23 24 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=4.565 $Y=2.02 $X2=3.63
+ $Y2=2.02
r118 19 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=2.105
+ $X2=3.545 $Y2=2.02
r119 19 21 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.545 $Y=2.105
+ $X2=3.545 $Y2=2.3
r120 18 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=1.935
+ $X2=3.375 $Y2=2.02
r121 18 32 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.375 $Y=1.935
+ $X2=3.375 $Y2=1.185
r122 15 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=0.89
+ $X2=3.34 $Y2=1.015
r123 4 38 600 $w=1.7e-07 $l=3.16307e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=2.065 $X2=5.11 $Y2=2.27
r124 3 21 600 $w=1.7e-07 $l=5.96657e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=1.945 $X2=3.545 $Y2=2.3
r125 2 42 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.235 $X2=5.15 $Y2=0.42
r126 1 15 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.595 $X2=3.34 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%A_1191_413# 1 2 7 9 14
c31 9 0 1.87801e-19 $X=6.09 $Y=2.02
r32 14 17 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.08 $Y=2.02
+ $X2=7.08 $Y2=2.21
r33 9 12 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.09 $Y=2.02 $X2=6.09
+ $Y2=2.21
r34 8 9 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=2.02 $X2=6.09
+ $Y2=2.02
r35 7 14 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=2.02
+ $X2=7.08 $Y2=2.02
r36 7 8 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.995 $Y=2.02
+ $X2=6.175 $Y2=2.02
r37 2 17 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=2.065 $X2=7.08 $Y2=2.21
r38 1 12 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=2.065 $X2=6.09 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%Q 1 2 7 10 14
r19 14 16 14.4879 $w=3.48e-07 $l=4.4e-07 $layer=LI1_cond $X=11.75 $Y=1.17
+ $X2=11.75 $Y2=1.61
r20 7 14 0.0987808 $w=3.48e-07 $l=3e-09 $layer=LI1_cond $X=11.75 $Y=1.167
+ $X2=11.75 $Y2=1.17
r21 7 10 17.6818 $w=3.48e-07 $l=5.37e-07 $layer=LI1_cond $X=11.75 $Y=1.167
+ $X2=11.75 $Y2=0.63
r22 2 16 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=11.565
+ $Y=1.485 $X2=11.74 $Y2=1.61
r23 1 10 182 $w=1.7e-07 $l=4.745e-07 $layer=licon1_NDIFF $count=1 $X=11.565
+ $Y=0.235 $X2=11.74 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%Q_N 1 2 9 13 18 21
c30 21 0 6.17411e-20 $X=12.745 $Y=1.15
c31 13 0 1.62009e-19 $X=12.61 $Y=1.62
r32 20 21 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.74 $Y=0.825
+ $X2=12.74 $Y2=1.15
r33 18 20 16.4563 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=12.635 $Y=0.4
+ $X2=12.635 $Y2=0.825
r34 14 21 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.74 $Y=1.535
+ $X2=12.74 $Y2=1.15
r35 13 15 14.2361 $w=3.88e-07 $l=4.6e-07 $layer=LI1_cond $X=12.63 $Y=1.62
+ $X2=12.63 $Y2=2.08
r36 13 14 6.24364 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=12.63 $Y=1.62
+ $X2=12.63 $Y2=1.535
r37 9 15 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=12.675 $Y=2.3
+ $X2=12.675 $Y2=2.08
r38 2 13 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=12.475
+ $Y=1.485 $X2=12.61 $Y2=1.62
r39 2 9 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.61 $Y2=2.3
r40 1 18 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=12.475
+ $Y=0.235 $X2=12.61 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__SDFRBP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 36 40 44 48 52
+ 56 60 62 64 67 68 70 71 72 74 79 91 105 112 117 123 126 129 132 135 138 142
+ 145
c218 60 0 1.91378e-19 $X=12.19 $Y=0.565
c219 44 0 1.79332e-19 $X=4.61 $Y=0.455
c220 30 0 1.34476e-19 $X=0.68 $Y=0.38
r221 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r222 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r223 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r224 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r225 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r226 127 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.53 $Y2=0
r227 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r228 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r229 121 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r230 121 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r231 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r232 118 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.275 $Y=0
+ $X2=12.19 $Y2=0
r233 118 120 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.275 $Y=0
+ $X2=12.65 $Y2=0
r234 117 141 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=13.167 $Y2=0
r235 117 120 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.995 $Y=0
+ $X2=12.65 $Y2=0
r236 116 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r237 116 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r238 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r239 113 135 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=11.365 $Y=0
+ $X2=11.227 $Y2=0
r240 113 115 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.365 $Y=0
+ $X2=11.73 $Y2=0
r241 112 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.19 $Y2=0
r242 112 115 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.73 $Y2=0
r243 111 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r244 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r245 108 111 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r246 107 110 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.43 $Y=0
+ $X2=10.81 $Y2=0
r247 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r248 105 135 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=11.09 $Y=0
+ $X2=11.227 $Y2=0
r249 105 110 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.09 $Y=0
+ $X2=10.81 $Y2=0
r250 104 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r251 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r252 101 104 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.97 $Y2=0
r253 101 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r254 100 103 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=8.97 $Y2=0
r255 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r256 98 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.08 $Y2=0
r257 98 100 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.59 $Y2=0
r258 97 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r259 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r260 94 97 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.67 $Y2=0
r261 93 96 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.67
+ $Y2=0
r262 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r263 91 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=7.08 $Y2=0
r264 91 96 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=6.67
+ $Y2=0
r265 90 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r266 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r267 87 90 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.37 $Y2=0
r268 87 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.53 $Y2=0
r269 86 89 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r270 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r271 84 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=2.56 $Y2=0
r272 84 86 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=2.99 $Y2=0
r273 83 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.07 $Y2=0
r274 83 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=0.69 $Y2=0
r275 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r276 80 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r277 80 82 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r278 79 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.04 $Y2=0
r279 79 82 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r280 76 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r281 74 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r282 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r283 72 124 0.128044 $w=4.8e-07 $l=4.5e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.69 $Y2=0
r284 72 145 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.23 $Y2=0
r285 70 103 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=9.085 $Y=0
+ $X2=8.97 $Y2=0
r286 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.085 $Y=0 $X2=9.17
+ $Y2=0
r287 69 107 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.255 $Y=0
+ $X2=9.43 $Y2=0
r288 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=0 $X2=9.17
+ $Y2=0
r289 67 89 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.37
+ $Y2=0
r290 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.61
+ $Y2=0
r291 66 93 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.83
+ $Y2=0
r292 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.61
+ $Y2=0
r293 62 141 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=13.08 $Y=0.085
+ $X2=13.167 $Y2=0
r294 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.08 $Y=0.085
+ $X2=13.08 $Y2=0.4
r295 58 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.19 $Y=0.085
+ $X2=12.19 $Y2=0
r296 58 60 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=12.19 $Y=0.085
+ $X2=12.19 $Y2=0.565
r297 54 135 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.227 $Y=0.085
+ $X2=11.227 $Y2=0
r298 54 56 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=11.227 $Y=0.085
+ $X2=11.227 $Y2=0.38
r299 50 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.17 $Y=0.085
+ $X2=9.17 $Y2=0
r300 50 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.17 $Y=0.085
+ $X2=9.17 $Y2=0.36
r301 46 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0
r302 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.08 $Y=0.085
+ $X2=7.08 $Y2=0.38
r303 42 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=0.085
+ $X2=4.61 $Y2=0
r304 42 44 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.61 $Y=0.085
+ $X2=4.61 $Y2=0.455
r305 38 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r306 38 40 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.74
r307 37 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.04 $Y2=0
r308 36 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.56 $Y2=0
r309 36 37 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.205 $Y2=0
r310 32 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r311 32 34 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.475
r312 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r313 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r314 9 64 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=12.895
+ $Y=0.235 $X2=13.08 $Y2=0.4
r315 8 60 182 $w=1.7e-07 $l=4.04166e-07 $layer=licon1_NDIFF $count=1 $X=12.025
+ $Y=0.235 $X2=12.19 $Y2=0.565
r316 7 56 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=11.085
+ $Y=0.235 $X2=11.255 $Y2=0.38
r317 6 52 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=8.985
+ $Y=0.235 $X2=9.17 $Y2=0.36
r318 5 48 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=6.825
+ $Y=0.235 $X2=7.08 $Y2=0.38
r319 4 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.33 $X2=4.61 $Y2=0.455
r320 3 40 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.595 $X2=2.56 $Y2=0.74
r321 2 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.33 $X2=2.04 $Y2=0.475
r322 1 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND CLK a_643_369# VNB nshort w=420000u l=150000u
+  ad=1.2874e+12p pd=1.423e+07u as=1.092e+11p ps=1.36e+06u
M1001 a_27_369# a_319_21# a_181_47# VPB phighvt w=640000u l=150000u
+  ad=3.328e+11p pd=3.6e+06u as=2.82e+11p ps=3.18e+06u
M1002 a_193_369# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.8575e+12p ps=1.806e+07u
M1003 Q a_2412_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1004 a_181_47# D a_193_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Q_N a_1587_329# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1006 a_1587_329# a_809_369# a_1514_47# VNB nshort w=640000u l=150000u
+  ad=2.524e+11p pd=2.22e+06u as=4.448e+11p ps=2.67e+06u
M1007 a_997_413# a_809_369# a_181_47# VPB phighvt w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1008 a_1129_21# a_997_413# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1009 a_1347_47# a_997_413# a_1129_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.092e+11p ps=1.36e+06u
M1010 VGND SET_B a_1879_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.058e+11p ps=1.82e+06u
M1011 VPWR a_1770_295# a_1712_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.218e+11p ps=1.42e+06u
M1012 a_181_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=8.82e+10p ps=1.26e+06u
M1013 VGND SCE a_319_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1014 a_1514_47# a_997_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1807_47# a_643_369# a_1587_329# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1016 a_1514_329# a_997_413# VPWR VPB phighvt w=840000u l=150000u
+  ad=1.806e+11p pd=2.11e+06u as=0p ps=0u
M1017 a_1587_329# a_643_369# a_1514_329# VPB phighvt w=840000u l=150000u
+  ad=4.137e+11p pd=3.99e+06u as=0p ps=0u
M1018 a_1879_47# a_1770_295# a_1807_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_2412_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1020 a_1770_295# a_1587_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1021 VPWR SCD a_27_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_265_47# D a_181_47# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1023 a_997_413# a_643_369# a_181_47# VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1024 a_1087_47# a_809_369# a_997_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1025 VGND a_1129_21# a_1087_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR SCE a_319_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1027 VPWR a_1587_329# a_2412_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1028 a_1587_329# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q_N a_1587_329# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1030 a_809_369# a_643_369# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1031 VGND a_319_21# a_265_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR SET_B a_1129_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1587_329# a_2412_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1034 VPWR CLK a_643_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1035 a_1081_413# a_643_369# a_997_413# VPB phighvt w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1036 a_809_369# a_643_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1037 VPWR a_1129_21# a_1081_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1770_295# a_1587_329# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1039 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1712_413# a_809_369# a_1587_329# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND SET_B a_1347_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

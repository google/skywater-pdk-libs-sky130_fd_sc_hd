* File: sky130_fd_sc_hd__a41o_1.spice
* Created: Thu Aug 27 14:06:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a41o_1.spice.pex"
.subckt sky130_fd_sc_hd__a41o_1  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_79_21#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.160875 AS=0.169 PD=1.145 PS=1.82 NRD=13.836 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1004 N_A_79_21#_M1004_d N_B1_M1004_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.183625 AS=0.160875 PD=1.215 PS=1.145 NRD=6.456 NRS=25.836 M=1 R=4.33333
+ SA=75000.8 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1002 A_381_47# N_A1_M1002_g N_A_79_21#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.183625 PD=0.92 PS=1.215 NRD=14.76 NRS=46.152 M=1 R=4.33333
+ SA=75001.5 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 A_465_47# N_A2_M1005_g A_381_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75002
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 A_561_47# N_A3_M1006_g A_465_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.10725 PD=0.98 PS=0.98 NRD=20.304 NRS=20.304 M=1 R=4.33333 SA=75002.4
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A4_M1009_g A_561_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.10725 PD=1.82 PS=0.98 NRD=0 NRS=20.304 M=1 R=4.33333 SA=75002.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_79_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1001 N_A_297_297#_M1001_d N_B1_M1001_g N_A_79_21#_M1001_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_297_297#_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_297_297#_M1008_d N_A2_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A3_M1003_g N_A_297_297#_M1008_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.165 PD=1.33 PS=1.33 NRD=4.9053 NRS=10.8153 M=1 R=6.66667
+ SA=75001.5 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1000 N_A_297_297#_M1000_d N_A4_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.165 PD=2.52 PS=1.33 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75002
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a41o_1.spice.SKY130_FD_SC_HD__A41O_1.pxi"
*
.ends
*
*

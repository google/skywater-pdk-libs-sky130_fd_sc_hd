* File: sky130_fd_sc_hd__o41ai_2.pex.spice
* Created: Tue Sep  1 19:26:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41AI_2%B1 1 3 6 8 10 13 15 21
r43 20 21 66.8119 $w=3.03e-07 $l=4.2e-07 $layer=POLY_cond $X=0.47 $Y=1.155
+ $X2=0.89 $Y2=1.155
r44 18 20 31.0198 $w=3.03e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.155
+ $X2=0.47 $Y2=1.155
r45 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r46 11 21 19.2026 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.89 $Y=1.31
+ $X2=0.89 $Y2=1.155
r47 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.89 $Y=1.31
+ $X2=0.89 $Y2=1.985
r48 8 21 19.2026 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.89 $Y=1 $X2=0.89
+ $Y2=1.155
r49 8 10 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.89 $Y=1 $X2=0.89
+ $Y2=0.56
r50 4 20 19.2026 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.47 $Y=1.31
+ $X2=0.47 $Y2=1.155
r51 4 6 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.47 $Y=1.31 $X2=0.47
+ $Y2=1.985
r52 1 20 19.2026 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.47 $Y=1 $X2=0.47
+ $Y2=1.155
r53 1 3 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.47 $Y=1 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A4 3 7 9 11 15 17 18
r51 21 23 53.4613 $w=2.84e-07 $l=3.15e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=2.145 $Y2=1.16
r52 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.145
+ $Y=1.16 $X2=2.145 $Y2=1.16
r53 17 18 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=1.635 $Y=1.175
+ $X2=2.095 $Y2=1.175
r54 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.25 $Y=1.305
+ $X2=2.25 $Y2=1.985
r55 9 13 17.6835 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.25 $Y2=1.305
r56 9 23 17.8204 $w=2.84e-07 $l=1.05e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.145 $Y2=1.16
r57 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r58 5 21 17.6835 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.83 $Y=1.305
+ $X2=1.83 $Y2=1.16
r59 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.83 $Y=1.305 $X2=1.83
+ $Y2=1.985
r60 1 21 17.6835 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.83 $Y=1.015
+ $X2=1.83 $Y2=1.16
r61 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.83 $Y=1.015
+ $X2=1.83 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A3 1 3 6 8 10 13 15 16 23
c51 23 0 1.77369e-19 $X=3.18 $Y=1.16
c52 6 0 6.60366e-20 $X=2.67 $Y=1.985
r53 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.18
+ $Y=1.16 $X2=3.18 $Y2=1.16
r54 21 23 17.9961 $w=3e-07 $l=9e-08 $layer=POLY_cond $X=3.09 $Y=1.16 $X2=3.18
+ $Y2=1.16
r55 19 21 83.9817 $w=3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.67 $Y=1.16 $X2=3.09
+ $Y2=1.16
r56 16 24 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.18 $Y2=1.175
r57 15 24 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.18 $Y2=1.175
r58 11 21 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.09 $Y=1.31
+ $X2=3.09 $Y2=1.16
r59 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.09 $Y=1.31
+ $X2=3.09 $Y2=1.985
r60 8 21 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.09 $Y=1.01 $X2=3.09
+ $Y2=1.16
r61 8 10 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.09 $Y=1.01 $X2=3.09
+ $Y2=0.56
r62 4 19 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.67 $Y=1.31 $X2=2.67
+ $Y2=1.16
r63 4 6 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.67 $Y=1.31 $X2=2.67
+ $Y2=1.985
r64 1 19 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.67 $Y=1.01 $X2=2.67
+ $Y2=1.16
r65 1 3 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.67 $Y=1.01 $X2=2.67
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A2 1 3 6 8 10 13 15 16
c52 16 0 3.71905e-19 $X=4.415 $Y=1.19
r53 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.32
+ $Y=1.16 $X2=4.32 $Y2=1.16
r54 16 23 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=4.415 $Y=1.175
+ $X2=4.32 $Y2=1.175
r55 15 23 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=3.955 $Y=1.175
+ $X2=4.32 $Y2=1.175
r56 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.49 $Y=1.295
+ $X2=4.49 $Y2=1.985
r57 8 11 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=4.49 $Y=1.142
+ $X2=4.49 $Y2=1.295
r58 8 22 33.4353 $w=3.05e-07 $l=1.7e-07 $layer=POLY_cond $X=4.49 $Y=1.142
+ $X2=4.32 $Y2=1.142
r59 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.49 $Y=0.99 $X2=4.49
+ $Y2=0.56
r60 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.07 $Y=1.295 $X2=4.07
+ $Y2=1.985
r61 1 22 49.1696 $w=3.05e-07 $l=2.5e-07 $layer=POLY_cond $X=4.07 $Y=1.142
+ $X2=4.32 $Y2=1.142
r62 1 4 19.3576 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=4.07 $Y=1.142
+ $X2=4.07 $Y2=1.295
r63 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.07 $Y=0.99 $X2=4.07
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A1 3 7 11 15 17 21 22 23 28
c45 17 0 1.94535e-19 $X=5.405 $Y=1.16
r46 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.57
+ $Y=1.16 $X2=5.57 $Y2=1.16
r47 23 29 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=5.795 $Y=1.175
+ $X2=5.57 $Y2=1.175
r48 22 29 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.335 $Y=1.175
+ $X2=5.57 $Y2=1.175
r49 21 22 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.875 $Y=1.175
+ $X2=5.335 $Y2=1.175
r50 18 20 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.91 $Y=1.16 $X2=5.33
+ $Y2=1.16
r51 17 28 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.16
+ $X2=5.57 $Y2=1.16
r52 17 20 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.405 $Y=1.16
+ $X2=5.33 $Y2=1.16
r53 13 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.33 $Y=1.295
+ $X2=5.33 $Y2=1.16
r54 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.33 $Y=1.295
+ $X2=5.33 $Y2=1.985
r55 9 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.33 $Y=1.025
+ $X2=5.33 $Y2=1.16
r56 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.33 $Y=1.025
+ $X2=5.33 $Y2=0.56
r57 5 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.91 $Y=1.295
+ $X2=4.91 $Y2=1.16
r58 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.91 $Y=1.295 $X2=4.91
+ $Y2=1.985
r59 1 18 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.91 $Y=1.025
+ $X2=4.91 $Y2=1.16
r60 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.91 $Y=1.025
+ $X2=4.91 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%VPWR 1 2 3 10 12 18 22 25 26 27 29 42 43 49
r72 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r74 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r75 39 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 37 40 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=4.83 $Y2=2.72
r77 37 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 36 39 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=4.83 $Y2=2.72
r79 36 37 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r80 34 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.14 $Y2=2.72
r81 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r82 33 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r84 30 46 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r85 30 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 29 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.14 $Y2=2.72
r87 29 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 27 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 27 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r90 25 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=4.83 $Y2=2.72
r91 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.955 $Y=2.72
+ $X2=5.12 $Y2=2.72
r92 24 42 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.75 $Y2=2.72
r93 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.12 $Y2=2.72
r94 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.635
+ $X2=5.12 $Y2=2.72
r95 20 22 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.12 $Y=2.635
+ $X2=5.12 $Y2=2
r96 16 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2.72
r97 16 18 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.14 $Y=2.635
+ $X2=1.14 $Y2=2
r98 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r99 10 46 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r100 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r101 3 22 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.985
+ $Y=1.485 $X2=5.12 $Y2=2
r102 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r103 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r104 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%Y 1 2 3 12 14 19 20 21 22 35 39
c46 35 0 1.15518e-19 $X=0.68 $Y=0.72
c47 19 0 6.60366e-20 $X=2.04 $Y=1.66
r48 39 40 2.19385 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.68 $Y=0.85
+ $X2=0.68 $Y2=0.885
r49 21 22 9.2696 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=0.727 $Y=1.19
+ $X2=0.727 $Y2=1.445
r50 20 39 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.68 $Y2=0.85
r51 20 35 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.68 $Y=0.825
+ $X2=0.68 $Y2=0.72
r52 20 21 13.7312 $w=2.33e-07 $l=2.8e-07 $layer=LI1_cond $X=0.727 $Y=0.91
+ $X2=0.727 $Y2=1.19
r53 20 40 1.226 $w=2.33e-07 $l=2.5e-08 $layer=LI1_cond $X=0.727 $Y=0.91
+ $X2=0.727 $Y2=0.885
r54 15 22 2.25663 $w=2.2e-07 $l=3.54119e-07 $layer=LI1_cond $X=0.845 $Y=1.555
+ $X2=0.515 $Y2=1.505
r55 14 19 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.555
+ $X2=2.04 $Y2=1.555
r56 14 15 53.9553 $w=2.18e-07 $l=1.03e-06 $layer=LI1_cond $X=1.875 $Y=1.555
+ $X2=0.845 $Y2=1.555
r57 10 22 4.1757 $w=2.82e-07 $l=2.31571e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.515 $Y2=1.505
r58 10 12 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.68 $Y=1.665
+ $X2=0.68 $Y2=2.34
r59 3 19 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.66
r60 2 22 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r61 2 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r62 1 35 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A_299_297# 1 2 3 12 14 15 17 20 21 24
r38 22 24 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.34 $Y=1.615
+ $X2=3.34 $Y2=1.62
r39 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.215 $Y=1.53
+ $X2=3.34 $Y2=1.615
r40 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.215 $Y=1.53
+ $X2=2.545 $Y2=1.53
r41 17 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.295
+ $X2=2.46 $Y2=2.38
r42 17 19 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.46 $Y=2.295
+ $X2=2.46 $Y2=1.62
r43 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.46 $Y=1.615
+ $X2=2.545 $Y2=1.53
r44 16 19 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.46 $Y=1.615
+ $X2=2.46 $Y2=1.62
r45 14 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=2.46 $Y2=2.38
r46 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.375 $Y=2.38
+ $X2=1.705 $Y2=2.38
r47 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.58 $Y=2.295
+ $X2=1.705 $Y2=2.38
r48 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=2.295
+ $X2=1.58 $Y2=2
r49 3 24 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.62
r50 2 27 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.3
r51 2 19 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.62
r52 1 12 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.485 $X2=1.62 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A_549_297# 1 2 9 11 12 15
r24 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.28 $Y=2.295
+ $X2=4.28 $Y2=2
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.115 $Y=2.38
+ $X2=4.28 $Y2=2.295
r26 11 12 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.115 $Y=2.38
+ $X2=3.045 $Y2=2.38
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.88 $Y=2.295
+ $X2=3.045 $Y2=2.38
r28 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.88 $Y=2.295
+ $X2=2.88 $Y2=2
r29 2 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.145
+ $Y=1.485 $X2=4.28 $Y2=2
r30 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A_743_297# 1 2 3 12 16 18 20 22 25 27
r39 20 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=1.615
+ $X2=5.58 $Y2=1.53
r40 20 22 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.58 $Y=1.615
+ $X2=5.58 $Y2=2.29
r41 19 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=1.53 $X2=4.7
+ $Y2=1.53
r42 18 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.455 $Y=1.53
+ $X2=5.58 $Y2=1.53
r43 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.455 $Y=1.53
+ $X2=4.785 $Y2=1.53
r44 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=1.615 $X2=4.7
+ $Y2=1.53
r45 14 16 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.7 $Y=1.615
+ $X2=4.7 $Y2=2.29
r46 13 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=1.53
+ $X2=3.82 $Y2=1.53
r47 12 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.615 $Y=1.53 $X2=4.7
+ $Y2=1.53
r48 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.615 $Y=1.53
+ $X2=3.945 $Y2=1.53
r49 3 29 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=1.485 $X2=5.54 $Y2=1.61
r50 3 22 400 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=1.485 $X2=5.54 $Y2=2.29
r51 2 27 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.7 $Y2=1.61
r52 2 16 400 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.7 $Y2=2.29
r53 1 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.715
+ $Y=1.485 $X2=3.86 $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%A_27_47# 1 2 3 4 5 6 7 22 24 26 28 31 32 33
+ 36 38 42 44 48 50 54 56 60 66 67 68 69
r136 58 60 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.54 $Y=0.735
+ $X2=5.54 $Y2=0.38
r137 57 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=0.82
+ $X2=4.7 $Y2=0.82
r138 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.375 $Y=0.82
+ $X2=5.54 $Y2=0.735
r139 56 57 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.375 $Y=0.82
+ $X2=4.865 $Y2=0.82
r140 52 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=0.735 $X2=4.7
+ $Y2=0.82
r141 52 54 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.7 $Y=0.735
+ $X2=4.7 $Y2=0.38
r142 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=0.82
+ $X2=3.86 $Y2=0.82
r143 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=0.82
+ $X2=4.7 $Y2=0.82
r144 50 51 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.535 $Y=0.82
+ $X2=4.025 $Y2=0.82
r145 46 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=0.735
+ $X2=3.86 $Y2=0.82
r146 46 48 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.86 $Y=0.735
+ $X2=3.86 $Y2=0.38
r147 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0.82
+ $X2=2.88 $Y2=0.82
r148 44 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=0.82
+ $X2=3.86 $Y2=0.82
r149 44 45 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.695 $Y=0.82
+ $X2=3.045 $Y2=0.82
r150 40 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=2.88 $Y2=0.82
r151 40 42 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.88 $Y=0.735
+ $X2=2.88 $Y2=0.38
r152 39 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0.82
+ $X2=2.04 $Y2=0.82
r153 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=0.82
+ $X2=2.88 $Y2=0.82
r154 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.715 $Y=0.82
+ $X2=2.205 $Y2=0.82
r155 34 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.735
+ $X2=2.04 $Y2=0.82
r156 34 36 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.04 $Y=0.735
+ $X2=2.04 $Y2=0.38
r157 32 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=2.04 $Y2=0.82
r158 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.875 $Y=0.82
+ $X2=1.265 $Y2=0.82
r159 29 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.14 $Y=0.735
+ $X2=1.265 $Y2=0.82
r160 29 31 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.14 $Y=0.735
+ $X2=1.14 $Y2=0.72
r161 28 65 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.14 $Y=0.465
+ $X2=1.14 $Y2=0.36
r162 28 31 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.14 $Y=0.465
+ $X2=1.14 $Y2=0.72
r163 27 63 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=0.215 $Y2=0.36
r164 26 65 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=0.36
+ $X2=1.14 $Y2=0.36
r165 26 27 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.36
+ $X2=0.345 $Y2=0.36
r166 22 63 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.36
r167 22 24 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.72
r168 7 60 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.405
+ $Y=0.235 $X2=5.54 $Y2=0.38
r169 6 54 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.565
+ $Y=0.235 $X2=4.7 $Y2=0.38
r170 5 48 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.715
+ $Y=0.235 $X2=3.86 $Y2=0.38
r171 4 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.38
r172 3 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r173 2 65 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r174 2 31 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.72
r175 1 63 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r176 1 24 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_2%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 46 47 48 50 72 73 76
r99 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r100 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r101 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r102 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r103 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r104 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r105 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r106 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r107 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r108 61 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r109 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r110 58 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.58
+ $Y2=0
r111 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.705 $Y=0
+ $X2=2.07 $Y2=0
r112 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r113 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r114 52 56 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r115 50 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.58
+ $Y2=0
r116 50 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r117 48 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r118 48 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r119 46 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.035 $Y=0
+ $X2=4.83 $Y2=0
r120 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.12
+ $Y2=0
r121 45 72 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.205 $Y=0
+ $X2=5.75 $Y2=0
r122 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=0 $X2=5.12
+ $Y2=0
r123 43 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.195 $Y=0
+ $X2=3.91 $Y2=0
r124 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=0 $X2=4.28
+ $Y2=0
r125 42 69 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.365 $Y=0
+ $X2=4.83 $Y2=0
r126 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=0 $X2=4.28
+ $Y2=0
r127 40 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=2.99 $Y2=0
r128 40 41 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=3.332 $Y2=0
r129 39 66 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r130 39 41 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=3.332
+ $Y2=0
r131 37 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.07 $Y2=0
r132 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.46
+ $Y2=0
r133 36 63 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.545 $Y=0
+ $X2=2.99 $Y2=0
r134 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.46
+ $Y2=0
r135 32 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=0.085
+ $X2=5.12 $Y2=0
r136 32 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.12 $Y=0.085
+ $X2=5.12 $Y2=0.38
r137 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0
r138 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.28 $Y=0.085
+ $X2=4.28 $Y2=0.38
r139 24 41 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.332 $Y=0.085
+ $X2=3.332 $Y2=0
r140 24 26 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=3.332 $Y=0.085
+ $X2=3.332 $Y2=0.38
r141 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r142 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.38
r143 16 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r144 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.38
r145 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=0.235 $X2=5.12 $Y2=0.38
r146 4 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.38
r147 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.38
r148 2 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.38
r149 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__a2111oi_0.spice.SKY130_FD_SC_HD__A2111OI_0.pxi
* Created: Thu Aug 27 13:58:51 2020
* 
x_PM_SKY130_FD_SC_HD__A2111OI_0%D1 N_D1_c_72_n N_D1_c_73_n N_D1_c_68_n
+ N_D1_M1008_g N_D1_c_74_n N_D1_M1007_g N_D1_c_69_n D1 D1 D1 N_D1_c_71_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%D1
x_PM_SKY130_FD_SC_HD__A2111OI_0%C1 N_C1_M1002_g N_C1_M1006_g C1 C1 C1 C1
+ N_C1_c_106_n PM_SKY130_FD_SC_HD__A2111OI_0%C1
x_PM_SKY130_FD_SC_HD__A2111OI_0%B1 N_B1_M1001_g N_B1_M1000_g B1 B1 N_B1_c_144_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%B1
x_PM_SKY130_FD_SC_HD__A2111OI_0%A1 N_A1_c_180_n N_A1_M1009_g N_A1_M1003_g
+ N_A1_c_181_n N_A1_c_176_n A1 A1 A1 N_A1_c_179_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%A1
x_PM_SKY130_FD_SC_HD__A2111OI_0%A2 N_A2_c_238_n N_A2_M1004_g N_A2_c_243_n
+ N_A2_M1005_g N_A2_c_239_n N_A2_c_240_n N_A2_c_244_n N_A2_c_245_n A2 A2 A2
+ N_A2_c_242_n PM_SKY130_FD_SC_HD__A2111OI_0%A2
x_PM_SKY130_FD_SC_HD__A2111OI_0%Y N_Y_M1008_d N_Y_M1000_d N_Y_M1007_s
+ N_Y_c_327_p N_Y_c_286_n N_Y_c_287_n N_Y_c_318_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_HD__A2111OI_0%Y
x_PM_SKY130_FD_SC_HD__A2111OI_0%A_313_369# N_A_313_369#_M1001_d
+ N_A_313_369#_M1005_d N_A_313_369#_c_349_n N_A_313_369#_c_342_n
+ N_A_313_369#_c_343_n N_A_313_369#_c_344_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%A_313_369#
x_PM_SKY130_FD_SC_HD__A2111OI_0%VPWR N_VPWR_M1009_d N_VPWR_c_372_n VPWR
+ N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_371_n N_VPWR_c_376_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%VPWR
x_PM_SKY130_FD_SC_HD__A2111OI_0%VGND N_VGND_M1008_s N_VGND_M1002_d
+ N_VGND_M1004_d N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n VGND N_VGND_c_414_n
+ N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n
+ PM_SKY130_FD_SC_HD__A2111OI_0%VGND
cc_1 VNB N_D1_c_68_n 0.0175908f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=0.73
cc_2 VNB N_D1_c_69_n 0.036729f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=0.805
cc_3 VNB D1 0.026041f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_D1_c_71_n 0.0323833f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.93
cc_5 VNB N_C1_M1002_g 0.0326082f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=0.73
cc_6 VNB C1 0.00359528f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.805
cc_7 VNB N_C1_c_106_n 0.0211701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_M1000_g 0.0309783f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=2.165
cc_9 VNB B1 0.00344245f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.805
cc_10 VNB N_B1_c_144_n 0.0220334f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.62
cc_11 VNB N_A1_M1003_g 0.0332964f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.77
cc_12 VNB N_A1_c_176_n 0.00859088f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_13 VNB A1 0.00563536f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB A1 0.00992749f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_15 VNB N_A1_c_179_n 0.0206134f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.93
cc_16 VNB N_A2_c_238_n 0.0165883f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.695
cc_17 VNB N_A2_c_239_n 0.0412299f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=2.165
cc_18 VNB N_A2_c_240_n 0.00653866f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=2.165
cc_19 VNB A2 0.0325179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_242_n 0.0297379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_286_n 0.0123718f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.62
cc_22 VNB N_Y_c_287_n 0.00808114f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_23 VNB Y 0.00744702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_371_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_407_n 0.014085f $X=-0.19 $Y=-0.24 $X2=0.7 $Y2=0.805
cc_26 VNB N_VGND_c_408_n 0.00499893f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_27 VNB N_VGND_c_409_n 0.012216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_410_n 0.0104832f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.93
cc_29 VNB N_VGND_c_411_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.85
cc_30 VNB N_VGND_c_412_n 0.0148983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_413_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=0.93
cc_32 VNB N_VGND_c_414_n 0.0242727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_415_n 0.0140696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_416_n 0.18561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_417_n 0.00510217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_D1_c_72_n 0.0273599f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.695
cc_37 VPB N_D1_c_73_n 0.0227331f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=1.695
cc_38 VPB N_D1_c_74_n 0.0174014f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.77
cc_39 VPB D1 0.0183922f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_40 VPB N_D1_c_71_n 0.0236853f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.93
cc_41 VPB N_C1_M1006_g 0.0287427f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=2.165
cc_42 VPB C1 0.00668905f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.805
cc_43 VPB N_C1_c_106_n 0.0141418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_B1_M1001_g 0.032384f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=0.73
cc_45 VPB B1 0.00670007f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.805
cc_46 VPB N_B1_c_144_n 0.0118425f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.62
cc_47 VPB N_A1_c_180_n 0.0155172f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.695
cc_48 VPB N_A1_c_181_n 0.0372961f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.805
cc_49 VPB N_A1_c_176_n 0.00389076f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_50 VPB A1 5.86836e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_51 VPB A1 0.0047054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A1_c_179_n 0.0151083f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.93
cc_53 VPB N_A2_c_243_n 0.0201805f $X=-0.19 $Y=1.305 $X2=0.7 $Y2=0.445
cc_54 VPB N_A2_c_244_n 0.0458956f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.805
cc_55 VPB N_A2_c_245_n 0.00567663f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.88
cc_56 VPB A2 0.0191029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A2_c_242_n 0.0221662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB Y 0.00677326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB Y 0.0173138f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=0.85
cc_60 VPB Y 0.0107083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_313_369#_c_342_n 0.00781726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_313_369#_c_343_n 0.0149545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_372_n 0.00557173f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.77
cc_64 VPB N_VPWR_c_373_n 0.0560342f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.88
cc_65 VPB N_VPWR_c_374_n 0.0253092f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_66 VPB N_VPWR_c_371_n 0.0658284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_376_n 0.0063111f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.93
cc_68 N_D1_c_68_n N_C1_M1002_g 0.0183957f $X=0.7 $Y=0.73 $X2=0 $Y2=0
cc_69 N_D1_c_71_n N_C1_M1002_g 0.0012297f $X=0.35 $Y=0.93 $X2=0 $Y2=0
cc_70 N_D1_c_72_n N_C1_M1006_g 0.0606851f $X=0.695 $Y=1.695 $X2=0 $Y2=0
cc_71 N_D1_c_71_n N_C1_M1006_g 0.00166782f $X=0.35 $Y=0.93 $X2=0 $Y2=0
cc_72 N_D1_c_72_n C1 0.00450543f $X=0.695 $Y=1.695 $X2=0 $Y2=0
cc_73 N_D1_c_71_n N_C1_c_106_n 0.00827852f $X=0.35 $Y=0.93 $X2=0 $Y2=0
cc_74 N_D1_c_68_n N_Y_c_287_n 0.0071923f $X=0.7 $Y=0.73 $X2=0 $Y2=0
cc_75 N_D1_c_69_n N_Y_c_287_n 0.0109211f $X=0.7 $Y=0.805 $X2=0 $Y2=0
cc_76 D1 N_Y_c_287_n 0.0124103f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_77 N_D1_c_72_n Y 0.0150698f $X=0.695 $Y=1.695 $X2=0 $Y2=0
cc_78 N_D1_c_74_n Y 0.00161223f $X=0.77 $Y=1.77 $X2=0 $Y2=0
cc_79 D1 Y 0.0581772f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_80 N_D1_c_71_n Y 0.0049653f $X=0.35 $Y=0.93 $X2=0 $Y2=0
cc_81 N_D1_c_74_n Y 0.00775495f $X=0.77 $Y=1.77 $X2=0 $Y2=0
cc_82 N_D1_c_73_n Y 0.0105212f $X=0.485 $Y=1.695 $X2=0 $Y2=0
cc_83 N_D1_c_74_n Y 0.00343428f $X=0.77 $Y=1.77 $X2=0 $Y2=0
cc_84 D1 Y 0.00647637f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_85 N_D1_c_74_n N_VPWR_c_373_n 0.00450273f $X=0.77 $Y=1.77 $X2=0 $Y2=0
cc_86 N_D1_c_74_n N_VPWR_c_371_n 0.00849017f $X=0.77 $Y=1.77 $X2=0 $Y2=0
cc_87 N_D1_c_68_n N_VGND_c_407_n 0.00342537f $X=0.7 $Y=0.73 $X2=0 $Y2=0
cc_88 N_D1_c_69_n N_VGND_c_407_n 0.00676693f $X=0.7 $Y=0.805 $X2=0 $Y2=0
cc_89 D1 N_VGND_c_407_n 0.00829011f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_90 N_D1_c_69_n N_VGND_c_410_n 2.42799e-19 $X=0.7 $Y=0.805 $X2=0 $Y2=0
cc_91 D1 N_VGND_c_410_n 0.00319028f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_92 N_D1_c_68_n N_VGND_c_412_n 0.00424946f $X=0.7 $Y=0.73 $X2=0 $Y2=0
cc_93 N_D1_c_68_n N_VGND_c_416_n 0.00673077f $X=0.7 $Y=0.73 $X2=0 $Y2=0
cc_94 D1 N_VGND_c_416_n 0.00624456f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_95 N_C1_c_106_n N_B1_M1001_g 0.0469588f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_96 N_C1_M1002_g N_B1_M1000_g 0.0231028f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_97 N_C1_M1002_g B1 5.95419e-19 $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_98 C1 B1 0.0544958f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_99 N_C1_M1002_g N_B1_c_144_n 0.0469588f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_100 C1 N_B1_c_144_n 0.0118518f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_101 N_C1_M1002_g N_Y_c_286_n 0.0159954f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_102 C1 N_Y_c_286_n 0.0234479f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_103 C1 N_Y_c_287_n 0.00782467f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_104 N_C1_c_106_n N_Y_c_287_n 0.00415784f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_105 N_C1_M1002_g Y 0.00442014f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_106 N_C1_M1006_g Y 0.00156352f $X=1.13 $Y=2.165 $X2=0 $Y2=0
cc_107 C1 Y 0.102244f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_108 N_C1_c_106_n Y 0.00305723f $X=1.04 $Y=1.22 $X2=0 $Y2=0
cc_109 N_C1_M1006_g Y 6.03196e-19 $X=1.13 $Y=2.165 $X2=0 $Y2=0
cc_110 C1 A_169_369# 0.00484557f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 C1 A_241_369# 0.00565829f $X=1.065 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_112 N_C1_M1006_g N_A_313_369#_c_344_n 7.60716e-19 $X=1.13 $Y=2.165 $X2=0
+ $Y2=0
cc_113 C1 N_A_313_369#_c_344_n 0.0304196f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_114 N_C1_M1006_g N_VPWR_c_373_n 0.0037867f $X=1.13 $Y=2.165 $X2=0 $Y2=0
cc_115 C1 N_VPWR_c_373_n 0.0128628f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_116 N_C1_M1006_g N_VPWR_c_371_n 0.00506666f $X=1.13 $Y=2.165 $X2=0 $Y2=0
cc_117 C1 N_VPWR_c_371_n 0.0126597f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_118 N_C1_M1002_g N_VGND_c_408_n 0.00177558f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_119 N_C1_M1002_g N_VGND_c_412_n 0.00422112f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_120 N_C1_M1002_g N_VGND_c_416_n 0.00577107f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_A1_M1003_g 0.0263656f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_122 B1 N_A1_M1003_g 0.00486323f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B1_c_144_n N_A1_M1003_g 0.0219886f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_124 N_B1_M1001_g N_A1_c_181_n 0.0176267f $X=1.49 $Y=2.165 $X2=0 $Y2=0
cc_125 B1 N_A1_c_181_n 0.00210869f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_A1_c_176_n 0.00457386f $X=1.49 $Y=2.165 $X2=0 $Y2=0
cc_127 B1 A1 5.73348e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_128 B1 A1 0.025105f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B1_c_144_n A1 3.24931e-19 $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_130 B1 A1 0.0127533f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B1_M1000_g N_Y_c_286_n 0.0156777f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_132 B1 N_Y_c_286_n 0.0292042f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B1_c_144_n N_Y_c_286_n 0.00448543f $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_134 N_B1_M1001_g N_A_313_369#_c_344_n 0.00733743f $X=1.49 $Y=2.165 $X2=0
+ $Y2=0
cc_135 B1 N_A_313_369#_c_344_n 0.0223874f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_136 N_B1_c_144_n N_A_313_369#_c_344_n 6.98824e-19 $X=1.61 $Y=1.22 $X2=0 $Y2=0
cc_137 N_B1_M1001_g N_VPWR_c_373_n 0.0054895f $X=1.49 $Y=2.165 $X2=0 $Y2=0
cc_138 N_B1_M1001_g N_VPWR_c_371_n 0.00980226f $X=1.49 $Y=2.165 $X2=0 $Y2=0
cc_139 N_B1_M1000_g N_VGND_c_408_n 0.00320636f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_140 N_B1_M1000_g N_VGND_c_414_n 0.00422112f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_141 N_B1_M1000_g N_VGND_c_416_n 0.00584081f $X=1.63 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A1_M1003_g N_A2_c_238_n 0.0472357f $X=2.06 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_143 A1 N_A2_c_238_n 0.00563404f $X=2.445 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_144 N_A1_c_180_n N_A2_c_243_n 0.0210578f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_145 A1 N_A2_c_239_n 0.00673154f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_146 A1 N_A2_c_240_n 0.00403146f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_147 A1 N_A2_c_240_n 4.42326e-19 $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A1_c_179_n N_A2_c_240_n 0.0181539f $X=2.46 $Y=1.235 $X2=0 $Y2=0
cc_149 A1 N_A2_c_244_n 0.00411778f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_150 N_A1_c_181_n N_A2_c_245_n 0.00998278f $X=2.075 $Y=1.595 $X2=0 $Y2=0
cc_151 A1 N_A2_c_245_n 0.00531235f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_152 N_A1_c_179_n N_A2_c_245_n 0.0162052f $X=2.46 $Y=1.235 $X2=0 $Y2=0
cc_153 N_A1_M1003_g A2 2.49469e-19 $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_154 A1 A2 0.0324856f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_155 A1 A2 0.0273754f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_156 A1 A2 0.0265642f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_157 N_A1_c_179_n A2 0.00110148f $X=2.46 $Y=1.235 $X2=0 $Y2=0
cc_158 N_A1_M1003_g N_A2_c_242_n 0.00111419f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A1_c_181_n N_A2_c_242_n 0.00121261f $X=2.075 $Y=1.595 $X2=0 $Y2=0
cc_160 A1 N_A2_c_242_n 4.02603e-19 $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_161 A1 N_A2_c_242_n 4.40277e-19 $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_162 A1 N_A2_c_242_n 4.87727e-19 $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_163 N_A1_c_179_n N_A2_c_242_n 0.0208234f $X=2.46 $Y=1.235 $X2=0 $Y2=0
cc_164 N_A1_M1003_g N_Y_c_286_n 0.00981702f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_165 A1 N_Y_c_286_n 0.0107811f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_166 A1 N_Y_c_286_n 3.70047e-19 $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A1_M1003_g N_Y_c_318_n 0.00661931f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A1_c_180_n N_A_313_369#_c_349_n 0.0125968f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_169 N_A1_c_181_n N_A_313_369#_c_349_n 0.0049549f $X=2.075 $Y=1.595 $X2=0
+ $Y2=0
cc_170 A1 N_A_313_369#_c_349_n 0.0092798f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_171 A1 N_A_313_369#_c_349_n 0.0121181f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_172 N_A1_c_179_n N_A_313_369#_c_349_n 0.00328726f $X=2.46 $Y=1.235 $X2=0
+ $Y2=0
cc_173 A1 N_A_313_369#_c_342_n 0.00503177f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_174 N_A1_c_180_n N_A_313_369#_c_344_n 0.00722207f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_175 N_A1_c_180_n N_VPWR_c_372_n 0.00434795f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_176 N_A1_c_180_n N_VPWR_c_373_n 0.00415375f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_177 N_A1_c_180_n N_VPWR_c_371_n 0.00592734f $X=1.92 $Y=1.77 $X2=0 $Y2=0
cc_178 N_A1_M1003_g N_VGND_c_409_n 0.00187505f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_179 A1 N_VGND_c_409_n 0.00954736f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_180 N_A1_M1003_g N_VGND_c_414_n 0.00505274f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_181 A1 N_VGND_c_414_n 0.00186056f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_182 N_A1_M1003_g N_VGND_c_416_n 0.00873617f $X=2.06 $Y=0.445 $X2=0 $Y2=0
cc_183 A1 N_VGND_c_416_n 0.00345788f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A2_c_238_n N_Y_c_286_n 9.45117e-19 $X=2.42 $Y=0.73 $X2=0 $Y2=0
cc_185 N_A2_c_238_n N_Y_c_318_n 0.00128877f $X=2.42 $Y=0.73 $X2=0 $Y2=0
cc_186 N_A2_c_243_n N_A_313_369#_c_349_n 0.0104776f $X=2.45 $Y=1.77 $X2=0 $Y2=0
cc_187 N_A2_c_244_n N_A_313_369#_c_342_n 0.0104667f $X=2.835 $Y=1.695 $X2=0
+ $Y2=0
cc_188 A2 N_A_313_369#_c_342_n 0.00639937f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_189 N_A2_c_243_n N_A_313_369#_c_344_n 3.15266e-19 $X=2.45 $Y=1.77 $X2=0 $Y2=0
cc_190 N_A2_c_243_n N_VPWR_c_372_n 0.00331648f $X=2.45 $Y=1.77 $X2=0 $Y2=0
cc_191 N_A2_c_243_n N_VPWR_c_374_n 0.00425094f $X=2.45 $Y=1.77 $X2=0 $Y2=0
cc_192 N_A2_c_243_n N_VPWR_c_371_n 0.0069728f $X=2.45 $Y=1.77 $X2=0 $Y2=0
cc_193 N_A2_c_238_n N_VGND_c_409_n 0.0100466f $X=2.42 $Y=0.73 $X2=0 $Y2=0
cc_194 N_A2_c_239_n N_VGND_c_409_n 0.0069583f $X=2.835 $Y=0.805 $X2=0 $Y2=0
cc_195 N_A2_c_238_n N_VGND_c_414_n 0.00367933f $X=2.42 $Y=0.73 $X2=0 $Y2=0
cc_196 N_A2_c_239_n N_VGND_c_415_n 0.00104172f $X=2.835 $Y=0.805 $X2=0 $Y2=0
cc_197 A2 N_VGND_c_415_n 0.00656683f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_198 N_A2_c_238_n N_VGND_c_416_n 0.00440171f $X=2.42 $Y=0.73 $X2=0 $Y2=0
cc_199 A2 N_VGND_c_416_n 0.00998581f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_200 Y N_VPWR_c_373_n 0.0275134f $X=0.605 $Y=2.125 $X2=0 $Y2=0
cc_201 N_Y_M1007_s N_VPWR_c_371_n 0.00238012f $X=0.4 $Y=1.845 $X2=0 $Y2=0
cc_202 Y N_VPWR_c_371_n 0.0157961f $X=0.605 $Y=2.125 $X2=0 $Y2=0
cc_203 N_Y_c_286_n N_VGND_M1002_d 0.00243865f $X=1.71 $Y=0.75 $X2=0 $Y2=0
cc_204 N_Y_c_286_n N_VGND_c_408_n 0.0184417f $X=1.71 $Y=0.75 $X2=0 $Y2=0
cc_205 N_Y_c_318_n N_VGND_c_409_n 0.00708715f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_206 N_Y_c_327_p N_VGND_c_412_n 0.014695f $X=0.915 $Y=0.42 $X2=0 $Y2=0
cc_207 N_Y_c_286_n N_VGND_c_412_n 0.00284415f $X=1.71 $Y=0.75 $X2=0 $Y2=0
cc_208 N_Y_c_287_n N_VGND_c_412_n 0.00288105f $X=1.04 $Y=0.75 $X2=0 $Y2=0
cc_209 N_Y_c_286_n N_VGND_c_414_n 0.00283681f $X=1.71 $Y=0.75 $X2=0 $Y2=0
cc_210 N_Y_c_318_n N_VGND_c_414_n 0.0164206f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_211 N_Y_M1008_d N_VGND_c_416_n 0.00229602f $X=0.775 $Y=0.235 $X2=0 $Y2=0
cc_212 N_Y_M1000_d N_VGND_c_416_n 0.00226885f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_213 N_Y_c_327_p N_VGND_c_416_n 0.00972398f $X=0.915 $Y=0.42 $X2=0 $Y2=0
cc_214 N_Y_c_286_n N_VGND_c_416_n 0.00986951f $X=1.71 $Y=0.75 $X2=0 $Y2=0
cc_215 N_Y_c_287_n N_VGND_c_416_n 0.0043017f $X=1.04 $Y=0.75 $X2=0 $Y2=0
cc_216 N_Y_c_318_n N_VGND_c_416_n 0.0121765f $X=1.845 $Y=0.445 $X2=0 $Y2=0
cc_217 A_169_369# N_VPWR_c_371_n 0.00558195f $X=0.845 $Y=1.845 $X2=1.04 $Y2=1.22
cc_218 A_241_369# N_VPWR_c_371_n 0.00489617f $X=1.205 $Y=1.845 $X2=1.04 $Y2=1.22
cc_219 N_A_313_369#_c_349_n N_VPWR_M1009_d 0.00673881f $X=2.54 $Y=1.995
+ $X2=-0.19 $Y2=1.305
cc_220 N_A_313_369#_c_349_n N_VPWR_c_372_n 0.0203701f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_221 N_A_313_369#_c_349_n N_VPWR_c_373_n 0.00247661f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_222 N_A_313_369#_c_344_n N_VPWR_c_373_n 0.0187174f $X=1.705 $Y=1.99 $X2=0
+ $Y2=0
cc_223 N_A_313_369#_c_349_n N_VPWR_c_374_n 0.00264253f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_224 N_A_313_369#_c_343_n N_VPWR_c_374_n 0.0214045f $X=2.705 $Y=2.33 $X2=0
+ $Y2=0
cc_225 N_A_313_369#_M1001_d N_VPWR_c_371_n 0.00223231f $X=1.565 $Y=1.845 $X2=0
+ $Y2=0
cc_226 N_A_313_369#_M1005_d N_VPWR_c_371_n 0.00250514f $X=2.525 $Y=1.845 $X2=0
+ $Y2=0
cc_227 N_A_313_369#_c_349_n N_VPWR_c_371_n 0.00963148f $X=2.54 $Y=1.995 $X2=0
+ $Y2=0
cc_228 N_A_313_369#_c_343_n N_VPWR_c_371_n 0.0125683f $X=2.705 $Y=2.33 $X2=0
+ $Y2=0
cc_229 N_A_313_369#_c_344_n N_VPWR_c_371_n 0.0122048f $X=1.705 $Y=1.99 $X2=0
+ $Y2=0
cc_230 N_VGND_c_416_n A_427_47# 0.00897657f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

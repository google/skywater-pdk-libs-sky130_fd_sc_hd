* File: sky130_fd_sc_hd__nor2_8.pex.spice
* Created: Tue Sep  1 19:17:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR2_8%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 72 73
r142 71 73 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.32 $Y=1.16
+ $X2=3.43 $Y2=1.16
r143 71 72 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r144 69 71 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.32 $Y2=1.16
r145 68 69 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.59 $Y=1.16
+ $X2=3.01 $Y2=1.16
r146 67 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.17 $Y=1.16
+ $X2=2.59 $Y2=1.16
r147 66 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.75 $Y=1.16
+ $X2=2.17 $Y2=1.16
r148 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.75 $Y2=1.16
r149 64 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r150 62 64 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.6 $Y=1.16 $X2=0.91
+ $Y2=1.16
r151 62 63 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r152 59 62 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.6 $Y2=1.16
r153 57 72 145.845 $w=1.98e-07 $l=2.63e-06 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=3.32 $Y2=1.175
r154 57 63 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=0.69 $Y=1.175 $X2=0.6
+ $Y2=1.175
r155 53 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.16
r156 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.43 $Y=1.325
+ $X2=3.43 $Y2=1.985
r157 50 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.16
r158 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r159 46 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.16
r160 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.01 $Y=1.325
+ $X2=3.01 $Y2=1.985
r161 43 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=1.16
r162 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r163 39 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.16
r164 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.59 $Y=1.325
+ $X2=2.59 $Y2=1.985
r165 36 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=1.16
r166 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.59 $Y=0.995
+ $X2=2.59 $Y2=0.56
r167 32 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.16
r168 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=1.325
+ $X2=2.17 $Y2=1.985
r169 29 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=1.16
r170 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.17 $Y=0.995
+ $X2=2.17 $Y2=0.56
r171 25 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r172 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r173 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r174 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r175 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r176 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r177 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r178 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r179 11 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r180 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r181 8 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r182 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r183 4 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r184 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r185 1 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r186 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_8%B 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 71 73
r143 72 73 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.37 $Y=1.16
+ $X2=6.79 $Y2=1.16
r144 70 72 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.355 $Y=1.16
+ $X2=6.37 $Y2=1.16
r145 70 71 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=6.355
+ $Y=1.16 $X2=6.355 $Y2=1.16
r146 68 70 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=5.95 $Y=1.16
+ $X2=6.355 $Y2=1.16
r147 67 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.53 $Y=1.16
+ $X2=5.95 $Y2=1.16
r148 66 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.11 $Y=1.16
+ $X2=5.53 $Y2=1.16
r149 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.69 $Y=1.16
+ $X2=5.11 $Y2=1.16
r150 64 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.27 $Y=1.16
+ $X2=4.69 $Y2=1.16
r151 62 64 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=3.975 $Y=1.16
+ $X2=4.27 $Y2=1.16
r152 62 63 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=3.975
+ $Y=1.16 $X2=3.975 $Y2=1.16
r153 59 62 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.85 $Y=1.16
+ $X2=3.975 $Y2=1.16
r154 57 71 84.5682 $w=1.98e-07 $l=1.525e-06 $layer=LI1_cond $X=4.83 $Y=1.175
+ $X2=6.355 $Y2=1.175
r155 57 63 47.4136 $w=1.98e-07 $l=8.55e-07 $layer=LI1_cond $X=4.83 $Y=1.175
+ $X2=3.975 $Y2=1.175
r156 53 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.79 $Y=1.325
+ $X2=6.79 $Y2=1.16
r157 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.79 $Y=1.325
+ $X2=6.79 $Y2=1.985
r158 50 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.79 $Y=0.995
+ $X2=6.79 $Y2=1.16
r159 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.79 $Y=0.995
+ $X2=6.79 $Y2=0.56
r160 46 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.325
+ $X2=6.37 $Y2=1.16
r161 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.37 $Y=1.325
+ $X2=6.37 $Y2=1.985
r162 43 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=0.995
+ $X2=6.37 $Y2=1.16
r163 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.37 $Y=0.995
+ $X2=6.37 $Y2=0.56
r164 39 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.16
r165 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.95 $Y=1.325
+ $X2=5.95 $Y2=1.985
r166 36 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=1.16
r167 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.95 $Y=0.995
+ $X2=5.95 $Y2=0.56
r168 32 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.53 $Y=1.325
+ $X2=5.53 $Y2=1.16
r169 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.53 $Y=1.325
+ $X2=5.53 $Y2=1.985
r170 29 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.53 $Y=0.995
+ $X2=5.53 $Y2=1.16
r171 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.53 $Y=0.995
+ $X2=5.53 $Y2=0.56
r172 25 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=1.325
+ $X2=5.11 $Y2=1.16
r173 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.11 $Y=1.325
+ $X2=5.11 $Y2=1.985
r174 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.11 $Y=0.995
+ $X2=5.11 $Y2=1.16
r175 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.11 $Y=0.995
+ $X2=5.11 $Y2=0.56
r176 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.16
r177 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.69 $Y=1.325
+ $X2=4.69 $Y2=1.985
r178 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=1.16
r179 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.69 $Y=0.995
+ $X2=4.69 $Y2=0.56
r180 11 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.325
+ $X2=4.27 $Y2=1.16
r181 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.27 $Y=1.325
+ $X2=4.27 $Y2=1.985
r182 8 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=0.995
+ $X2=4.27 $Y2=1.16
r183 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.27 $Y=0.995
+ $X2=4.27 $Y2=0.56
r184 4 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.325
+ $X2=3.85 $Y2=1.16
r185 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.85 $Y=1.325
+ $X2=3.85 $Y2=1.985
r186 1 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=0.995
+ $X2=3.85 $Y2=1.16
r187 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.85 $Y=0.995
+ $X2=3.85 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_8%A_27_297# 1 2 3 4 5 6 7 8 9 28 30 32 36 38 42
+ 44 48 50 52 53 54 58 60 64 66 70 72 76 81 83 85 90 91 92
r103 74 76 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7 $Y=2.295 $X2=7
+ $Y2=1.96
r104 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.285 $Y=2.38
+ $X2=6.16 $Y2=2.38
r105 72 74 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.875 $Y=2.38
+ $X2=7 $Y2=2.295
r106 72 73 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.875 $Y=2.38
+ $X2=6.285 $Y2=2.38
r107 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=2.295
+ $X2=6.16 $Y2=2.38
r108 68 70 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.16 $Y=2.295
+ $X2=6.16 $Y2=1.96
r109 67 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.445 $Y=2.38
+ $X2=5.32 $Y2=2.38
r110 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.035 $Y=2.38
+ $X2=6.16 $Y2=2.38
r111 66 67 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.035 $Y=2.38
+ $X2=5.445 $Y2=2.38
r112 62 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=2.295
+ $X2=5.32 $Y2=2.38
r113 62 64 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.32 $Y=2.295
+ $X2=5.32 $Y2=1.96
r114 61 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.605 $Y=2.38
+ $X2=4.48 $Y2=2.38
r115 60 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.195 $Y=2.38
+ $X2=5.32 $Y2=2.38
r116 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.195 $Y=2.38
+ $X2=4.605 $Y2=2.38
r117 56 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=2.295
+ $X2=4.48 $Y2=2.38
r118 56 58 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.48 $Y=2.295
+ $X2=4.48 $Y2=1.96
r119 55 89 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.765 $Y=2.38
+ $X2=3.64 $Y2=2.38
r120 54 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.355 $Y=2.38
+ $X2=4.48 $Y2=2.38
r121 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.355 $Y=2.38
+ $X2=3.765 $Y2=2.38
r122 53 89 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.295
+ $X2=3.64 $Y2=2.38
r123 52 87 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.64 $Y=1.665
+ $X2=3.64 $Y2=1.56
r124 52 53 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=3.64 $Y=1.665
+ $X2=3.64 $Y2=2.295
r125 51 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.925 $Y=1.56
+ $X2=2.8 $Y2=1.56
r126 50 87 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.515 $Y=1.56
+ $X2=3.64 $Y2=1.56
r127 50 51 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=3.515 $Y=1.56
+ $X2=2.925 $Y2=1.56
r128 46 85 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.8 $Y=1.665
+ $X2=2.8 $Y2=1.56
r129 46 48 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.8 $Y=1.665
+ $X2=2.8 $Y2=2.3
r130 45 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.56
+ $X2=1.96 $Y2=1.56
r131 44 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=1.56
+ $X2=2.8 $Y2=1.56
r132 44 45 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=2.675 $Y=1.56
+ $X2=2.085 $Y2=1.56
r133 40 83 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=1.56
r134 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.96 $Y=1.665
+ $X2=1.96 $Y2=2.3
r135 39 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=1.56
+ $X2=1.12 $Y2=1.56
r136 38 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.56
+ $X2=1.96 $Y2=1.56
r137 38 39 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=1.56
+ $X2=1.245 $Y2=1.56
r138 34 81 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=1.56
r139 34 36 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.12 $Y=1.665
+ $X2=1.12 $Y2=2.3
r140 33 79 4.31179 $w=2.1e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.56
+ $X2=0.247 $Y2=1.56
r141 32 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.56
+ $X2=1.12 $Y2=1.56
r142 32 33 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.56
+ $X2=0.405 $Y2=1.56
r143 28 79 2.86543 $w=3.15e-07 $l=1.05e-07 $layer=LI1_cond $X=0.247 $Y=1.665
+ $X2=0.247 $Y2=1.56
r144 28 30 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=0.247 $Y=1.665
+ $X2=0.247 $Y2=2.3
r145 9 76 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.865
+ $Y=1.485 $X2=7 $Y2=1.96
r146 8 70 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.025
+ $Y=1.485 $X2=6.16 $Y2=1.96
r147 7 64 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.185
+ $Y=1.485 $X2=5.32 $Y2=1.96
r148 6 58 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.48 $Y2=1.96
r149 5 89 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=2.3
r150 5 87 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.485 $X2=3.64 $Y2=1.62
r151 4 85 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=1.62
r152 4 48 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.8 $Y2=2.3
r153 3 83 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.62
r154 3 42 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.3
r155 2 81 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r156 2 36 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r157 1 79 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r158 1 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_8%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 36 37 38
+ 40 59 60 63
r100 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r101 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r102 57 60 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=7.13 $Y2=2.72
r103 56 59 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=7.13 $Y2=2.72
r104 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r105 54 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r107 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r108 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 48 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r111 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 45 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r113 45 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 40 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r115 40 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r116 38 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 38 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r118 36 53 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=2.72
+ $X2=2.99 $Y2=2.72
r119 36 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=2.72
+ $X2=3.22 $Y2=2.72
r120 35 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=2.72
+ $X2=3.45 $Y2=2.72
r121 35 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=2.72
+ $X2=3.22 $Y2=2.72
r122 33 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.07 $Y2=2.72
r123 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=2.72
+ $X2=2.38 $Y2=2.72
r124 32 53 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.99 $Y2=2.72
r125 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.38 $Y2=2.72
r126 30 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=2.72
+ $X2=1.54 $Y2=2.72
r128 29 50 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=2.07 $Y2=2.72
r129 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.665 $Y=2.72
+ $X2=1.54 $Y2=2.72
r130 25 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r131 25 27 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2
r132 21 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2.72
r133 21 23 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.38 $Y=2.635
+ $X2=2.38 $Y2=2
r134 17 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2.72
r135 17 19 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.54 $Y=2.635
+ $X2=1.54 $Y2=2
r136 13 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r137 13 15 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2
r138 4 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.085
+ $Y=1.485 $X2=3.22 $Y2=2
r139 3 23 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.245
+ $Y=1.485 $X2=2.38 $Y2=2
r140 2 19 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=2
r141 1 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 41 42 45 47
+ 51 53 57 59 63 67 69 70 71 75 79 81 83 87 91 93 95 99 103 105 106 107 108 109
+ 110 111 112 114 115
r225 113 115 9.45786 $w=7.33e-07 $l=5.4e-07 $layer=LI1_cond $X=6.992 $Y=0.905
+ $X2=6.992 $Y2=1.445
r226 113 114 2.2976 $w=4.47e-07 $l=1.86652e-07 $layer=LI1_cond $X=6.992 $Y=0.905
+ $X2=6.845 $Y2=0.815
r227 101 115 2.37703 $w=4.07e-07 $l=3.24731e-07 $layer=LI1_cond $X=6.58 $Y=1.615
+ $X2=6.865 $Y2=1.53
r228 101 103 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.58 $Y=1.615
+ $X2=6.58 $Y2=1.62
r229 97 114 2.2976 $w=4.47e-07 $l=3.06716e-07 $layer=LI1_cond $X=6.58 $Y=0.725
+ $X2=6.845 $Y2=0.815
r230 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.58 $Y=0.725
+ $X2=6.58 $Y2=0.39
r231 96 111 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0.815
+ $X2=5.74 $Y2=0.815
r232 95 114 4.75417 $w=1.8e-07 $l=4.3e-07 $layer=LI1_cond $X=6.415 $Y=0.815
+ $X2=6.845 $Y2=0.815
r233 95 96 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.415 $Y=0.815
+ $X2=5.905 $Y2=0.815
r234 94 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.865 $Y=1.53
+ $X2=5.74 $Y2=1.53
r235 93 115 4.61444 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=6.455 $Y=1.53
+ $X2=6.865 $Y2=1.53
r236 93 94 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.455 $Y=1.53
+ $X2=5.865 $Y2=1.53
r237 89 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.74 $Y=1.615
+ $X2=5.74 $Y2=1.53
r238 89 91 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.74 $Y=1.615
+ $X2=5.74 $Y2=1.62
r239 85 111 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.74 $Y=0.725
+ $X2=5.74 $Y2=0.815
r240 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.74 $Y=0.725
+ $X2=5.74 $Y2=0.39
r241 84 109 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=0.815
+ $X2=4.9 $Y2=0.815
r242 83 111 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=0.815
+ $X2=5.74 $Y2=0.815
r243 83 84 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.575 $Y=0.815
+ $X2=5.065 $Y2=0.815
r244 82 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.025 $Y=1.53
+ $X2=4.9 $Y2=1.53
r245 81 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.615 $Y=1.53
+ $X2=5.74 $Y2=1.53
r246 81 82 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.615 $Y=1.53
+ $X2=5.025 $Y2=1.53
r247 77 110 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.9 $Y=1.615
+ $X2=4.9 $Y2=1.53
r248 77 79 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.9 $Y=1.615 $X2=4.9
+ $Y2=1.62
r249 73 109 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.9 $Y=0.725 $X2=4.9
+ $Y2=0.815
r250 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.9 $Y=0.725
+ $X2=4.9 $Y2=0.39
r251 72 108 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=0.815
+ $X2=4.06 $Y2=0.815
r252 71 109 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=0.815
+ $X2=4.9 $Y2=0.815
r253 71 72 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.735 $Y=0.815
+ $X2=4.225 $Y2=0.815
r254 69 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.775 $Y=1.53
+ $X2=4.9 $Y2=1.53
r255 69 70 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.775 $Y=1.53
+ $X2=4.185 $Y2=1.53
r256 65 70 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.06 $Y=1.615
+ $X2=4.185 $Y2=1.53
r257 65 67 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.06 $Y=1.615
+ $X2=4.06 $Y2=1.62
r258 61 108 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.06 $Y=0.725
+ $X2=4.06 $Y2=0.815
r259 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.06 $Y=0.725
+ $X2=4.06 $Y2=0.39
r260 60 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=3.22 $Y2=0.815
r261 59 108 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0.815
+ $X2=4.06 $Y2=0.815
r262 59 60 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.895 $Y=0.815
+ $X2=3.385 $Y2=0.815
r263 55 107 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.815
r264 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.22 $Y=0.725
+ $X2=3.22 $Y2=0.39
r265 54 106 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0.815
+ $X2=2.38 $Y2=0.815
r266 53 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=3.22 $Y2=0.815
r267 53 54 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.055 $Y=0.815
+ $X2=2.545 $Y2=0.815
r268 49 106 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.815
r269 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=0.725
+ $X2=2.38 $Y2=0.39
r270 48 105 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=0.815
+ $X2=1.54 $Y2=0.815
r271 47 106 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=2.38 $Y2=0.815
r272 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.215 $Y=0.815
+ $X2=1.705 $Y2=0.815
r273 43 105 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.815
r274 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.39
r275 41 105 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=1.54 $Y2=0.815
r276 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.815
+ $X2=0.865 $Y2=0.815
r277 37 42 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.815
r278 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.7 $Y2=0.39
r279 12 103 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.445
+ $Y=1.485 $X2=6.58 $Y2=1.62
r280 11 91 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.605
+ $Y=1.485 $X2=5.74 $Y2=1.62
r281 10 79 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=1.485 $X2=4.9 $Y2=1.62
r282 9 67 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.485 $X2=4.06 $Y2=1.62
r283 8 99 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.445
+ $Y=0.235 $X2=6.58 $Y2=0.39
r284 7 87 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.605
+ $Y=0.235 $X2=5.74 $Y2=0.39
r285 6 75 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.765
+ $Y=0.235 $X2=4.9 $Y2=0.39
r286 5 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.925
+ $Y=0.235 $X2=4.06 $Y2=0.39
r287 4 57 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.39
r288 3 51 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.235 $X2=2.38 $Y2=0.39
r289 2 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r290 1 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2_8%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 52 56 60 62 64 67 68 70 71 73 74 76 77 78 79 81 82 83 105 113 117
r141 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r142 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r143 108 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r144 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r145 105 116 4.3 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.915 $Y=0 $X2=7.137
+ $Y2=0
r146 105 107 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.915 $Y=0
+ $X2=6.67 $Y2=0
r147 104 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r148 104 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r149 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r150 101 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=0
+ $X2=5.32 $Y2=0
r151 101 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=0
+ $X2=5.75 $Y2=0
r152 100 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r153 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r154 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r155 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r156 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r157 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r158 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r159 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r160 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r161 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r162 85 110 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r163 85 87 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.69 $Y2=0
r164 83 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r165 83 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r166 81 103 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=5.75 $Y2=0
r167 81 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=0 $X2=6.16
+ $Y2=0
r168 80 107 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.245 $Y=0
+ $X2=6.67 $Y2=0
r169 80 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=0 $X2=6.16
+ $Y2=0
r170 78 99 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r171 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.48
+ $Y2=0
r172 76 96 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r173 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.64
+ $Y2=0
r174 75 99 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.725 $Y=0
+ $X2=4.37 $Y2=0
r175 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.64
+ $Y2=0
r176 73 93 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=2.53 $Y2=0
r177 73 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.8
+ $Y2=0
r178 72 96 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r179 72 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.8
+ $Y2=0
r180 70 90 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r181 70 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r182 69 93 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.53 $Y2=0
r183 69 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r184 67 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r185 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r186 66 90 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.61 $Y2=0
r187 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r188 62 116 3.13784 $w=2.9e-07 $l=1.17346e-07 $layer=LI1_cond $X=7.06 $Y=0.085
+ $X2=7.137 $Y2=0
r189 62 64 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=7.06 $Y=0.085
+ $X2=7.06 $Y2=0.39
r190 58 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=0.085
+ $X2=6.16 $Y2=0
r191 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.16 $Y=0.085
+ $X2=6.16 $Y2=0.39
r192 54 113 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0
r193 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.32 $Y=0.085
+ $X2=5.32 $Y2=0.39
r194 53 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0 $X2=4.48
+ $Y2=0
r195 52 113 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0 $X2=5.32
+ $Y2=0
r196 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.235 $Y=0
+ $X2=4.565 $Y2=0
r197 48 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0
r198 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0.39
r199 44 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0
r200 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.64 $Y=0.085
+ $X2=3.64 $Y2=0.39
r201 40 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r202 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.39
r203 36 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r204 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r205 32 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r206 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r207 28 110 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r208 28 30 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r209 9 64 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.865
+ $Y=0.235 $X2=7 $Y2=0.39
r210 8 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.235 $X2=6.16 $Y2=0.39
r211 7 56 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.185
+ $Y=0.235 $X2=5.32 $Y2=0.39
r212 6 50 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.345
+ $Y=0.235 $X2=4.48 $Y2=0.39
r213 5 46 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.39
r214 4 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.8 $Y2=0.39
r215 3 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r216 2 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r217 1 30 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__mux2_1.spice.pex
* Created: Thu Aug 27 14:27:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__MUX2_1%A_76_199# 1 2 9 12 16 17 19 20 22 25 26 27 29
+ 33
c77 29 0 1.9931e-19 $X=1.36 $Y=0.54
r78 29 31 10.0255 $w=4.32e-07 $l=3.55e-07 $layer=LI1_cond $X=1.36 $Y=0.54
+ $X2=1.715 $Y2=0.54
r79 26 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r80 26 33 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r81 25 27 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.557 $Y=1.16
+ $X2=0.557 $Y2=0.995
r82 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r83 20 22 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.445 $Y=2.04
+ $X2=2.235 $Y2=2.04
r84 19 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.36 $Y=1.955
+ $X2=1.445 $Y2=2.04
r85 18 29 6.24874 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.36 $Y=0.825
+ $X2=1.36 $Y2=0.54
r86 18 19 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.36 $Y=0.825
+ $X2=1.36 $Y2=1.955
r87 16 29 7.19232 $w=4.32e-07 $l=2.40832e-07 $layer=LI1_cond $X=1.27 $Y=0.74
+ $X2=1.36 $Y2=0.54
r88 16 17 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.27 $Y=0.74
+ $X2=0.685 $Y2=0.74
r89 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.825
+ $X2=0.685 $Y2=0.74
r90 14 27 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.6 $Y=0.825 $X2=0.6
+ $Y2=0.995
r91 12 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r92 9 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
r93 2 22 300 $w=1.7e-07 $l=7.0993e-07 $layer=licon1_PDIFF $count=2 $X=1.605
+ $Y=1.87 $X2=2.235 $Y2=2.04
r94 1 31 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.715 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%S 3 7 11 15 18 19 20 21 22 24 25 28 29 37 43
c92 24 0 1.44221e-19 $X=0.995 $Y=1.16
c93 3 0 4.3721e-20 $X=1.015 $Y=0.445
r94 41 43 1.7512 $w=1.88e-07 $l=3e-08 $layer=LI1_cond $X=2.965 $Y=1.535
+ $X2=2.995 $Y2=1.535
r95 37 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.545
+ $X2=3.38 $Y2=1.71
r96 37 39 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.545
+ $X2=3.38 $Y2=1.38
r97 29 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.545 $X2=3.38 $Y2=1.545
r98 28 41 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.535
+ $X2=2.965 $Y2=1.535
r99 28 29 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=3.022 $Y=1.535
+ $X2=3.38 $Y2=1.535
r100 28 43 1.57608 $w=1.88e-07 $l=2.7e-08 $layer=LI1_cond $X=3.022 $Y=1.535
+ $X2=2.995 $Y2=1.535
r101 25 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=1.325
r102 25 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.16
+ $X2=0.995 $Y2=0.995
r103 24 27 9.59627 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.007 $Y=1.16
+ $X2=1.007 $Y2=1.325
r104 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r105 21 28 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.88 $Y=1.63
+ $X2=2.88 $Y2=1.535
r106 21 22 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.88 $Y=1.63
+ $X2=2.88 $Y2=2.295
r107 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.795 $Y=2.38
+ $X2=2.88 $Y2=2.295
r108 19 20 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=2.795 $Y=2.38
+ $X2=1.105 $Y2=2.38
r109 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.02 $Y=2.295
+ $X2=1.105 $Y2=2.38
r110 18 27 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.02 $Y=2.295
+ $X2=1.02 $Y2=1.325
r111 15 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.44 $Y=2.08
+ $X2=3.44 $Y2=1.71
r112 11 39 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=3.44 $Y=0.445
+ $X2=3.44 $Y2=1.38
r113 7 35 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.015 $Y=2.08
+ $X2=1.015 $Y2=1.325
r114 3 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.015 $Y=0.445
+ $X2=1.015 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%A1 3 7 11 12 14 15 17 18 26
c63 14 0 1.6555e-19 $X=2.435 $Y=1.7
c64 12 0 1.44221e-19 $X=1.7 $Y=0.98
c65 11 0 4.3721e-20 $X=1.7 $Y=0.98
r66 26 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.545
+ $X2=2.54 $Y2=1.71
r67 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.545 $X2=2.54 $Y2=1.545
r68 18 27 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.545
r69 17 18 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.53 $Y=0.85
+ $X2=2.53 $Y2=1.19
r70 16 27 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=2.53 $Y=1.615 $X2=2.53
+ $Y2=1.545
r71 14 16 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.435 $Y=1.7
+ $X2=2.53 $Y2=1.615
r72 14 15 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.435 $Y=1.7
+ $X2=1.785 $Y2=1.7
r73 12 21 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.7 $Y=0.98
+ $X2=1.495 $Y2=0.98
r74 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=0.98 $X2=1.7 $Y2=0.98
r75 9 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=1.615
+ $X2=1.785 $Y2=1.7
r76 9 11 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.7 $Y=1.615 $X2=1.7
+ $Y2=0.98
r77 7 29 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.6 $Y=2.08 $X2=2.6
+ $Y2=1.71
r78 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=0.815
+ $X2=1.495 $Y2=0.98
r79 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.495 $Y=0.815
+ $X2=1.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%A0 1 3 4 5 8 11 12 15 16
r51 15 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=0.98
+ $X2=2.18 $Y2=1.145
r52 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=0.98
+ $X2=2.18 $Y2=0.815
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.18
+ $Y=0.98 $X2=2.18 $Y2=0.98
r54 12 16 8.80047 $w=2.73e-07 $l=2.1e-07 $layer=LI1_cond $X=2.127 $Y=1.19
+ $X2=2.127 $Y2=0.98
r55 11 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.12 $Y=1.645 $X2=2.12
+ $Y2=1.145
r56 8 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.12 $Y=0.445
+ $X2=2.12 $Y2=0.815
r57 4 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.045 $Y=1.72
+ $X2=2.12 $Y2=1.645
r58 4 5 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.045 $Y=1.72
+ $X2=1.605 $Y2=1.72
r59 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.53 $Y=1.795
+ $X2=1.605 $Y2=1.72
r60 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.53 $Y=1.795 $X2=1.53
+ $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%A_505_21# 1 2 9 13 15 22 25 26 30 33
c56 13 0 1.6555e-19 $X=2.96 $Y=2.08
r57 32 33 81.8491 $w=2.12e-07 $l=3.6e-07 $layer=POLY_cond $X=2.6 $Y=0.98
+ $X2=2.96 $Y2=0.98
r58 28 30 6.60547 $w=4.08e-07 $l=2.35e-07 $layer=LI1_cond $X=3.65 $Y=2.08
+ $X2=3.885 $Y2=2.08
r59 25 30 1.83547 $w=3.4e-07 $l=2.05e-07 $layer=LI1_cond $X=3.885 $Y=1.875
+ $X2=3.885 $Y2=2.08
r60 24 26 3.22182 $w=2.92e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.885 $Y=1.065
+ $X2=3.795 $Y2=0.98
r61 24 25 27.4553 $w=3.38e-07 $l=8.1e-07 $layer=LI1_cond $X=3.885 $Y=1.065
+ $X2=3.885 $Y2=1.875
r62 20 26 3.22182 $w=2.92e-07 $l=1.75425e-07 $layer=LI1_cond $X=3.657 $Y=0.895
+ $X2=3.795 $Y2=0.98
r63 20 22 20.6969 $w=2.43e-07 $l=4.4e-07 $layer=LI1_cond $X=3.657 $Y=0.895
+ $X2=3.657 $Y2=0.455
r64 18 33 6.82075 $w=2.12e-07 $l=3e-08 $layer=POLY_cond $X=2.99 $Y=0.98 $X2=2.96
+ $Y2=0.98
r65 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=0.98 $X2=2.99 $Y2=0.98
r66 15 26 3.35233 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.535 $Y=0.98
+ $X2=3.795 $Y2=0.98
r67 15 17 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.535 $Y=0.98
+ $X2=2.99 $Y2=0.98
r68 11 33 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.96 $Y=1.115
+ $X2=2.96 $Y2=0.98
r69 11 13 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=2.96 $Y=1.115
+ $X2=2.96 $Y2=2.08
r70 7 32 10.9192 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.6 $Y=0.845 $X2=2.6
+ $Y2=0.98
r71 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.6 $Y=0.845 $X2=2.6
+ $Y2=0.445
r72 2 28 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.87 $X2=3.65 $Y2=2.04
r73 1 22 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%X 1 2 10 13 14 15 16 17
r20 17 30 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.34
r21 16 17 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=2.21
r22 13 14 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=1.495
r23 11 16 7.15547 $w=3.33e-07 $l=2.08e-07 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.87
r24 11 13 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.66
r25 10 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.175 $Y=0.825
+ $X2=0.175 $Y2=1.495
r26 9 15 10.0782 $w=2.53e-07 $l=2.23e-07 $layer=LI1_cond $X=0.217 $Y=0.698
+ $X2=0.217 $Y2=0.475
r27 9 10 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=0.217 $Y=0.698
+ $X2=0.217 $Y2=0.825
r28 2 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r29 2 13 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r30 1 15 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%VPWR 1 2 9 15 18 19 20 22 32 33 36
r40 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r42 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r43 30 37 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=0.68 $Y2=2.72
r46 27 29 145.16 $w=1.68e-07 $l=2.225e-06 $layer=LI1_cond $X=0.765 $Y=2.72
+ $X2=2.99 $Y2=2.72
r47 22 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.68 $Y2=2.72
r48 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 20 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 20 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 18 29 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.22 $Y2=2.72
r53 17 32 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.305 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=2.72
+ $X2=3.22 $Y2=2.72
r55 13 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r56 13 15 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.04
r57 9 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.66 $X2=0.68
+ $Y2=2.34
r58 7 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635 $X2=0.68
+ $Y2=2.72
r59 7 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r60 2 15 600 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.87 $X2=3.22 $Y2=2.04
r61 1 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r62 1 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__MUX2_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 33 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r58 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r59 30 39 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.06
+ $Y2=0
r60 30 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.91
+ $Y2=0
r61 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r62 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r63 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r64 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r65 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r66 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r68 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r69 22 39 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=3.06
+ $Y2=0
r70 22 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.53
+ $Y2=0
r71 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r72 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r73 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 11 39 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.06 $Y2=0
r76 11 13 8.67743 $w=5.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.06 $Y2=0.455
r77 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r78 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r79 2 13 91 $w=1.7e-07 $l=6.55839e-07 $layer=licon1_NDIFF $count=2 $X=2.675
+ $Y=0.235 $X2=3.23 $Y2=0.455
r80 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* NGSPICE file created from sky130_fd_sc_hd__o2111ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_1163_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.40285e+12p pd=2.282e+07u as=1.08e+12p ps=1.016e+07u
M1001 VPWR C1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.63335e+12p ps=2.328e+07u
M1002 Y A2 a_1163_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR D1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1163_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=1.27725e+12p ps=1.303e+07u
M1006 a_803_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1163_297# A2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A2 a_1163_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_803_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_445_47# B1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=7.02e+11p pd=7.36e+06u as=0p ps=0u
M1015 VPWR B1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_47# D1 Y VNB nshort w=650000u l=150000u
+  ad=8.645e+11p pd=9.16e+06u as=3.51e+11p ps=3.68e+06u
M1017 a_445_47# B1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A1 a_1163_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_27_47# D1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_445_47# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_803_47# B1 a_445_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Y D1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_803_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR D1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_47# C1 a_445_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_803_47# B1 a_445_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_803_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND A2 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR C1 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND A2 a_803_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_445_47# C1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_47# C1 a_445_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1163_297# A2 Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1163_297# A1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Y D1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Y C1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Y B1 VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 Y D1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__clkdlybuf4s18_2.pxi.spice
* Created: Tue Sep  1 19:00:46 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A N_A_M1000_g N_A_c_75_n N_A_M1004_g A
+ N_A_c_76_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_27_47# N_A_27_47#_M1000_s
+ N_A_27_47#_M1004_s N_A_27_47#_M1003_g N_A_27_47#_M1009_g N_A_27_47#_c_106_n
+ N_A_27_47#_c_112_n N_A_27_47#_c_107_n N_A_27_47#_c_108_n N_A_27_47#_c_113_n
+ N_A_27_47#_c_114_n N_A_27_47#_c_109_n N_A_27_47#_c_110_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_227_47# N_A_227_47#_M1003_d
+ N_A_227_47#_M1009_d N_A_227_47#_M1005_g N_A_227_47#_M1007_g
+ N_A_227_47#_c_175_n N_A_227_47#_c_168_n N_A_227_47#_c_169_n
+ N_A_227_47#_c_170_n N_A_227_47#_c_171_n N_A_227_47#_c_172_n
+ N_A_227_47#_c_173_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_227_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_334_47# N_A_334_47#_M1005_s
+ N_A_334_47#_M1007_s N_A_334_47#_M1001_g N_A_334_47#_M1002_g
+ N_A_334_47#_c_231_n N_A_334_47#_M1008_g N_A_334_47#_M1006_g
+ N_A_334_47#_c_234_n N_A_334_47#_c_235_n N_A_334_47#_c_244_n
+ N_A_334_47#_c_236_n N_A_334_47#_c_237_n N_A_334_47#_c_245_n
+ N_A_334_47#_c_246_n N_A_334_47#_c_238_n N_A_334_47#_c_239_n
+ N_A_334_47#_c_295_p N_A_334_47#_c_240_n N_A_334_47#_c_241_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%A_334_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VPWR N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_M1006_d N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n VPWR N_VPWR_c_333_n N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_326_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%X N_X_M1001_s N_X_M1002_s N_X_c_370_n
+ N_X_c_374_n N_X_c_371_n N_X_c_372_n X X X N_X_c_376_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VGND N_VGND_M1000_d N_VGND_M1005_d
+ N_VGND_M1008_d N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n VGND N_VGND_c_418_n N_VGND_c_419_n
+ N_VGND_c_420_n N_VGND_c_421_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_2%VGND
cc_1 VNB N_A_M1000_g 0.0392118f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.445
cc_2 VNB N_A_c_75_n 0.02846f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.305
cc_3 VNB N_A_c_76_n 0.0123232f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_4 VNB N_A_27_47#_M1003_g 0.0235085f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_M1009_g 5.30872e-19 $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_6 VNB N_A_27_47#_c_106_n 0.0187625f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.182
cc_7 VNB N_A_27_47#_c_107_n 0.0034131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_108_n 0.0101565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_109_n 0.00322944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_110_n 0.0275331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_227_47#_M1005_g 0.0255972f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_12 VNB N_A_227_47#_M1007_g 6.5763e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_227_47#_c_168_n 0.00646638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_227_47#_c_169_n 0.00767495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_227_47#_c_170_n 0.0567465f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_227_47#_c_171_n 9.51146e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_227_47#_c_172_n 0.00323153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_227_47#_c_173_n 0.00173909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_334_47#_M1001_g 0.0330137f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_20 VNB N_A_334_47#_M1002_g 5.21807e-19 $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_21 VNB N_A_334_47#_c_231_n 0.0130324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_334_47#_M1008_g 0.0368784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_334_47#_M1006_g 5.20615e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_334_47#_c_234_n 0.0120052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_334_47#_c_235_n 0.00443493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_334_47#_c_236_n 0.00471131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_334_47#_c_237_n 0.00338658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_334_47#_c_238_n 0.00266415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_334_47#_c_239_n 6.26893e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_334_47#_c_240_n 0.016953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_334_47#_c_241_n 0.001023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_326_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_370_n 0.0131408f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_34 VNB N_X_c_371_n 0.00117225f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.182
cc_35 VNB N_X_c_372_n 0.0079518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_412_n 0.00557365f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_37 VNB N_VGND_c_413_n 0.00579861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_414_n 0.0102019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_415_n 0.0228552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_416_n 0.0329153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_417_n 0.00708926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_418_n 0.0171347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_419_n 0.0208366f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_420_n 0.00632006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_421_n 0.207654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_A_c_75_n 0.00413708f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.305
cc_47 VPB N_A_M1004_g 0.028617f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.985
cc_48 VPB N_A_27_47#_M1009_g 0.036778f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_49 VPB N_A_27_47#_c_112_n 0.0331199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_113_n 0.00454327f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_47#_c_114_n 0.00970379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_109_n 0.00160595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_227_47#_M1007_g 0.0409174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_227_47#_c_175_n 0.00621365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_227_47#_c_171_n 0.00884179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_334_47#_M1002_g 0.0217151f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_57 VPB N_A_334_47#_M1006_g 0.0236223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_334_47#_c_244_n 0.00783868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_334_47#_c_245_n 0.00580323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_334_47#_c_246_n 0.00405362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_334_47#_c_239_n 0.002759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_327_n 0.00557247f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_63 VPB N_VPWR_c_328_n 0.00600372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_329_n 0.0101727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_330_n 0.0400699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_331_n 0.0316997f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_332_n 0.00794987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_333_n 0.0178855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_334_n 0.0202676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_335_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_326_n 0.0517767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_370_n 0.00495107f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_73 VPB N_X_c_374_n 0.00639874f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_74 N_A_M1000_g N_A_27_47#_M1003_g 0.0204132f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_c_75_n N_A_27_47#_M1009_g 0.0252071f $X=0.48 $Y=1.305 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_A_27_47#_c_106_n 0.00814049f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_M1004_g N_A_27_47#_c_112_n 0.0132942f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_A_27_47#_c_107_n 0.0102304f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_c_76_n N_A_27_47#_c_107_n 0.00999367f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_A_27_47#_c_108_n 0.00376303f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_A_27_47#_c_108_n 0.00425739f $X=0.48 $Y=1.305 $X2=0 $Y2=0
cc_82 N_A_c_76_n N_A_27_47#_c_108_n 0.0274014f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_A_27_47#_c_113_n 0.011714f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_c_76_n N_A_27_47#_c_113_n 0.0089583f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_75_n N_A_27_47#_c_114_n 0.00404637f $X=0.48 $Y=1.305 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_A_27_47#_c_114_n 0.00423547f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_c_76_n N_A_27_47#_c_114_n 0.0287201f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_A_27_47#_c_109_n 0.00292861f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_c_75_n N_A_27_47#_c_109_n 0.00610333f $X=0.48 $Y=1.305 $X2=0 $Y2=0
cc_90 N_A_c_76_n N_A_27_47#_c_109_n 0.0173767f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_c_75_n N_A_27_47#_c_110_n 0.0143452f $X=0.48 $Y=1.305 $X2=0 $Y2=0
cc_92 N_A_c_76_n N_A_27_47#_c_110_n 2.33591e-19 $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_M1004_g N_VPWR_c_327_n 0.00708566f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_M1004_g N_VPWR_c_333_n 0.0054895f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_M1004_g N_VPWR_c_326_n 0.0110389f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_M1000_g N_VGND_c_412_n 0.00318627f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_M1000_g N_VGND_c_418_n 0.00435476f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_M1000_g N_VGND_c_421_n 0.00714481f $X=0.48 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1009_g N_A_227_47#_c_175_n 0.00887531f $X=1.045 $Y=2.075 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_M1003_g N_A_227_47#_c_168_n 0.0109006f $X=1.045 $Y=0.56 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_107_n N_A_227_47#_c_168_n 0.0111634f $X=0.73 $Y=0.82 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_109_n N_A_227_47#_c_168_n 0.0106055f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_110_n N_A_227_47#_c_170_n 0.00689859f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_113_n N_A_227_47#_c_171_n 0.0113718f $X=0.73 $Y=1.545 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_109_n N_A_227_47#_c_171_n 0.0128084f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_110_n N_A_227_47#_c_171_n 0.0130383f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_109_n N_A_227_47#_c_173_n 0.0127166f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_110_n N_A_227_47#_c_173_n 0.00178354f $X=0.97 $Y=1.16 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_113_n N_VPWR_M1004_d 0.00239473f $X=0.73 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_27_47#_M1009_g N_VPWR_c_327_n 0.00323342f $X=1.045 $Y=2.075 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_113_n N_VPWR_c_327_n 0.0263277f $X=0.73 $Y=1.545 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_110_n N_VPWR_c_327_n 4.33882e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_27_47#_M1009_g N_VPWR_c_331_n 0.00666027f $X=1.045 $Y=2.075 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_112_n N_VPWR_c_333_n 0.0221174f $X=0.265 $Y=1.965 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1004_s N_VPWR_c_326_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_M1009_g N_VPWR_c_326_n 0.013117f $X=1.045 $Y=2.075 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_112_n N_VPWR_c_326_n 0.0130273f $X=0.265 $Y=1.965 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_c_107_n N_VGND_M1000_d 0.00272434f $X=0.73 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_27_47#_M1003_g N_VGND_c_412_n 0.00516205f $X=1.045 $Y=0.56 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_c_107_n N_VGND_c_412_n 0.0247699f $X=0.73 $Y=0.82 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_110_n N_VGND_c_412_n 4.28992e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1003_g N_VGND_c_416_n 0.00604919f $X=1.045 $Y=0.56 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_107_n N_VGND_c_416_n 0.00174068f $X=0.73 $Y=0.82 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_106_n N_VGND_c_418_n 0.0191713f $X=0.265 $Y=0.435 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_107_n N_VGND_c_418_n 0.0022703f $X=0.73 $Y=0.82 $X2=0 $Y2=0
cc_126 N_A_27_47#_M1000_s N_VGND_c_421_n 0.00218082f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_M1003_g N_VGND_c_421_n 0.011047f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_106_n N_VGND_c_421_n 0.0124046f $X=0.265 $Y=0.435 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_107_n N_VGND_c_421_n 0.00843414f $X=0.73 $Y=0.82 $X2=0 $Y2=0
cc_130 N_A_227_47#_M1005_g N_A_334_47#_M1001_g 0.0181287f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_131 N_A_227_47#_M1007_g N_A_334_47#_M1002_g 0.0239768f $X=2.025 $Y=2.075
+ $X2=0 $Y2=0
cc_132 N_A_227_47#_M1005_g N_A_334_47#_c_235_n 0.00954382f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_133 N_A_227_47#_c_172_n N_A_334_47#_c_235_n 0.0349233f $X=1.275 $Y=0.435
+ $X2=0 $Y2=0
cc_134 N_A_227_47#_M1007_g N_A_334_47#_c_244_n 0.0141015f $X=2.025 $Y=2.075
+ $X2=0 $Y2=0
cc_135 N_A_227_47#_c_171_n N_A_334_47#_c_244_n 0.0635588f $X=1.275 $Y=1.8 $X2=0
+ $Y2=0
cc_136 N_A_227_47#_M1005_g N_A_334_47#_c_236_n 0.0111577f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_137 N_A_227_47#_c_169_n N_A_334_47#_c_236_n 0.0169822f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_227_47#_c_170_n N_A_334_47#_c_236_n 0.00205431f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_227_47#_M1005_g N_A_334_47#_c_237_n 0.00418166f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_140 N_A_227_47#_c_168_n N_A_334_47#_c_237_n 0.0132713f $X=1.355 $Y=1.075
+ $X2=0 $Y2=0
cc_141 N_A_227_47#_c_169_n N_A_334_47#_c_237_n 0.0264204f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_227_47#_c_170_n N_A_334_47#_c_237_n 0.0072072f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_227_47#_M1007_g N_A_334_47#_c_245_n 0.0142437f $X=2.025 $Y=2.075
+ $X2=0 $Y2=0
cc_144 N_A_227_47#_c_169_n N_A_334_47#_c_245_n 0.0146737f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_227_47#_c_170_n N_A_334_47#_c_245_n 0.00198517f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_227_47#_M1007_g N_A_334_47#_c_246_n 0.00423476f $X=2.025 $Y=2.075
+ $X2=0 $Y2=0
cc_147 N_A_227_47#_c_169_n N_A_334_47#_c_246_n 0.0230874f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_A_227_47#_c_170_n N_A_334_47#_c_246_n 0.00702766f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_227_47#_c_171_n N_A_334_47#_c_246_n 0.0132713f $X=1.275 $Y=1.8 $X2=0
+ $Y2=0
cc_150 N_A_227_47#_M1005_g N_A_334_47#_c_238_n 0.00242676f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_151 N_A_227_47#_c_170_n N_A_334_47#_c_238_n 0.00110315f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_227_47#_M1007_g N_A_334_47#_c_239_n 0.00334444f $X=2.025 $Y=2.075
+ $X2=0 $Y2=0
cc_153 N_A_227_47#_c_169_n N_A_334_47#_c_239_n 6.81451e-19 $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_227_47#_c_170_n N_A_334_47#_c_239_n 9.45436e-19 $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_227_47#_c_170_n N_A_334_47#_c_240_n 0.0110408f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_227_47#_c_169_n N_A_334_47#_c_241_n 0.0146301f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_227_47#_c_170_n N_A_334_47#_c_241_n 6.36921e-19 $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_227_47#_M1007_g N_VPWR_c_328_n 0.00856683f $X=2.025 $Y=2.075 $X2=0
+ $Y2=0
cc_159 N_A_227_47#_M1007_g N_VPWR_c_331_n 0.00666027f $X=2.025 $Y=2.075 $X2=0
+ $Y2=0
cc_160 N_A_227_47#_c_175_n N_VPWR_c_331_n 0.0210373f $X=1.275 $Y=1.965 $X2=0
+ $Y2=0
cc_161 N_A_227_47#_M1009_d N_VPWR_c_326_n 0.00213418f $X=1.135 $Y=1.665 $X2=0
+ $Y2=0
cc_162 N_A_227_47#_M1007_g N_VPWR_c_326_n 0.0133223f $X=2.025 $Y=2.075 $X2=0
+ $Y2=0
cc_163 N_A_227_47#_c_175_n N_VPWR_c_326_n 0.0124461f $X=1.275 $Y=1.965 $X2=0
+ $Y2=0
cc_164 N_A_227_47#_M1007_g X 8.87225e-19 $X=2.025 $Y=2.075 $X2=0 $Y2=0
cc_165 N_A_227_47#_M1005_g N_X_c_376_n 3.97021e-19 $X=2.025 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_227_47#_M1005_g N_VGND_c_413_n 0.00549393f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_167 N_A_227_47#_M1005_g N_VGND_c_416_n 0.00515476f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_168 N_A_227_47#_c_172_n N_VGND_c_416_n 0.0166557f $X=1.275 $Y=0.435 $X2=0
+ $Y2=0
cc_169 N_A_227_47#_M1003_d N_VGND_c_421_n 0.00300709f $X=1.135 $Y=0.235 $X2=0
+ $Y2=0
cc_170 N_A_227_47#_M1005_g N_VGND_c_421_n 0.00860111f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_171 N_A_227_47#_c_172_n N_VGND_c_421_n 0.0105515f $X=1.275 $Y=0.435 $X2=0
+ $Y2=0
cc_172 N_A_334_47#_c_245_n N_VPWR_M1007_d 0.00364896f $X=2.375 $Y=1.545 $X2=0
+ $Y2=0
cc_173 N_A_334_47#_M1002_g N_VPWR_c_328_n 0.00785658f $X=2.665 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_334_47#_c_245_n N_VPWR_c_328_n 0.0324986f $X=2.375 $Y=1.545 $X2=0
+ $Y2=0
cc_175 N_A_334_47#_M1006_g N_VPWR_c_330_n 0.02111f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_334_47#_c_244_n N_VPWR_c_331_n 0.0210489f $X=1.795 $Y=1.965 $X2=0
+ $Y2=0
cc_177 N_A_334_47#_M1002_g N_VPWR_c_334_n 0.0054895f $X=2.665 $Y=1.985 $X2=0
+ $Y2=0
cc_178 N_A_334_47#_M1006_g N_VPWR_c_334_n 0.00389548f $X=3.095 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_334_47#_M1007_s N_VPWR_c_326_n 0.00213418f $X=1.67 $Y=1.665 $X2=0
+ $Y2=0
cc_180 N_A_334_47#_M1002_g N_VPWR_c_326_n 0.0102438f $X=2.665 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_A_334_47#_M1006_g N_VPWR_c_326_n 0.00711603f $X=3.095 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_334_47#_c_244_n N_VPWR_c_326_n 0.0124497f $X=1.795 $Y=1.965 $X2=0
+ $Y2=0
cc_183 N_A_334_47#_M1001_g N_X_c_370_n 5.6795e-19 $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_334_47#_M1002_g N_X_c_370_n 8.91465e-19 $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_334_47#_c_231_n N_X_c_370_n 0.00487596f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_334_47#_M1008_g N_X_c_370_n 0.00243579f $X=3.095 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_334_47#_M1006_g N_X_c_370_n 0.00384105f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_334_47#_c_234_n N_X_c_370_n 0.00758359f $X=3.095 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_334_47#_c_238_n N_X_c_370_n 0.00445012f $X=2.46 $Y=1.075 $X2=0 $Y2=0
cc_190 N_A_334_47#_c_239_n N_X_c_370_n 0.00612992f $X=2.46 $Y=1.46 $X2=0 $Y2=0
cc_191 N_A_334_47#_c_295_p N_X_c_370_n 0.0123998f $X=2.675 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_334_47#_M1002_g N_X_c_374_n 0.00266781f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_334_47#_c_231_n N_X_c_374_n 0.00435155f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_334_47#_M1006_g N_X_c_374_n 0.0052416f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_195 N_A_334_47#_c_245_n N_X_c_374_n 0.0077915f $X=2.375 $Y=1.545 $X2=0 $Y2=0
cc_196 N_A_334_47#_c_239_n N_X_c_374_n 0.00304905f $X=2.46 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A_334_47#_c_295_p N_X_c_374_n 0.00964897f $X=2.675 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_334_47#_M1001_g N_X_c_371_n 0.00319838f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A_334_47#_M1008_g N_X_c_371_n 0.00729481f $X=3.095 $Y=0.445 $X2=0 $Y2=0
cc_200 N_A_334_47#_c_236_n N_X_c_371_n 0.00771024f $X=2.375 $Y=0.82 $X2=0 $Y2=0
cc_201 N_A_334_47#_M1008_g N_X_c_372_n 0.00592877f $X=3.095 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A_334_47#_c_238_n N_X_c_372_n 0.0016135f $X=2.46 $Y=1.075 $X2=0 $Y2=0
cc_203 N_A_334_47#_M1002_g X 0.0148115f $X=2.665 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_334_47#_M1006_g X 0.0239821f $X=3.095 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_334_47#_M1001_g N_X_c_376_n 0.00618879f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A_334_47#_c_231_n N_X_c_376_n 0.00307003f $X=3.02 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_334_47#_M1008_g N_X_c_376_n 0.00777605f $X=3.095 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A_334_47#_c_295_p N_X_c_376_n 0.00360088f $X=2.675 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_334_47#_c_236_n N_VGND_M1005_d 0.00484875f $X=2.375 $Y=0.82 $X2=0
+ $Y2=0
cc_210 N_A_334_47#_M1001_g N_VGND_c_413_n 0.0053316f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_334_47#_c_236_n N_VGND_c_413_n 0.0296837f $X=2.375 $Y=0.82 $X2=0
+ $Y2=0
cc_212 N_A_334_47#_M1008_g N_VGND_c_415_n 0.0124506f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_213 N_A_334_47#_c_235_n N_VGND_c_416_n 0.0191269f $X=1.795 $Y=0.435 $X2=0
+ $Y2=0
cc_214 N_A_334_47#_c_236_n N_VGND_c_416_n 0.00239634f $X=2.375 $Y=0.82 $X2=0
+ $Y2=0
cc_215 N_A_334_47#_M1001_g N_VGND_c_419_n 0.00534477f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_334_47#_M1008_g N_VGND_c_419_n 0.00392237f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_334_47#_M1005_s N_VGND_c_421_n 0.00213973f $X=1.67 $Y=0.235 $X2=0
+ $Y2=0
cc_218 N_A_334_47#_M1001_g N_VGND_c_421_n 0.00993061f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_334_47#_M1008_g N_VGND_c_421_n 0.00649335f $X=3.095 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_334_47#_c_235_n N_VGND_c_421_n 0.0123353f $X=1.795 $Y=0.435 $X2=0
+ $Y2=0
cc_221 N_A_334_47#_c_236_n N_VGND_c_421_n 0.00633292f $X=2.375 $Y=0.82 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_326_n N_X_M1002_s 0.00223231f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_330_n X 0.0656615f $X=3.405 $Y=1.965 $X2=0 $Y2=0
cc_224 N_VPWR_c_334_n X 0.0260842f $X=3.32 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_326_n X 0.015831f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_226 N_X_c_376_n N_VGND_c_415_n 0.0293052f $X=2.88 $Y=0.435 $X2=0 $Y2=0
cc_227 N_X_c_376_n N_VGND_c_419_n 0.0238818f $X=2.88 $Y=0.435 $X2=0 $Y2=0
cc_228 N_X_M1001_s N_VGND_c_421_n 0.00223815f $X=2.74 $Y=0.235 $X2=0 $Y2=0
cc_229 N_X_c_372_n N_VGND_c_421_n 0.00104252f $X=3.072 $Y=0.945 $X2=0 $Y2=0
cc_230 N_X_c_376_n N_VGND_c_421_n 0.0158854f $X=2.88 $Y=0.435 $X2=0 $Y2=0

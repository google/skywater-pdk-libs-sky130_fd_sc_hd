* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_394_47# a_256_243# a_286_413# VNB nshort w=360000u l=150000u
+  ad=1.806e+11p pd=1.76e+06u as=1.35e+11p ps=1.47e+06u
M1001 a_464_315# a_286_413# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.533e+11p pd=2.52e+06u as=1.3369e+12p ps=1.205e+07u
M1002 a_1094_47# a_464_315# a_1012_47# VNB nshort w=420000u l=150000u
+  ad=1.722e+11p pd=1.66e+06u as=1.092e+11p ps=1.36e+06u
M1003 a_464_315# a_286_413# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=6.8955e+11p ps=6.89e+06u
M1004 VGND CLK a_1094_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_47# GATE a_109_369# VPB phighvt w=640000u l=150000u
+  ad=2.235e+11p pd=2.03e+06u as=1.344e+11p ps=1.7e+06u
M1006 a_256_147# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1007 a_382_413# a_256_147# a_286_413# VPB phighvt w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=1.386e+11p ps=1.5e+06u
M1008 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=2.433e+11p pd=2.86e+06u as=0p ps=0u
M1009 GCLK a_1012_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1010 a_109_369# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_256_147# a_256_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1012 VPWR CLK a_1012_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 GCLK a_1012_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1014 a_256_147# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1015 VPWR a_256_147# a_256_243# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.629e+11p ps=1.8e+06u
M1016 a_1012_47# a_464_315# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_464_315# a_382_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_464_315# a_394_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_286_413# a_256_147# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_286_413# a_256_243# a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_16.spice.SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16.pxi
* Created: Thu Aug 27 14:23:14 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A N_A_M1012_g N_A_c_124_n
+ N_A_M1009_g N_A_M1022_g N_A_c_125_n N_A_M1019_g N_A_M1026_g N_A_c_126_n
+ N_A_M1021_g N_A_M1039_g N_A_c_127_n N_A_M1038_g A A N_A_c_123_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A_110_47# N_A_110_47#_M1012_d
+ N_A_110_47#_M1026_d N_A_110_47#_M1009_s N_A_110_47#_M1021_s
+ N_A_110_47#_M1002_g N_A_110_47#_M1000_g N_A_110_47#_M1003_g
+ N_A_110_47#_M1001_g N_A_110_47#_M1004_g N_A_110_47#_M1005_g
+ N_A_110_47#_M1007_g N_A_110_47#_M1006_g N_A_110_47#_M1008_g
+ N_A_110_47#_M1010_g N_A_110_47#_M1015_g N_A_110_47#_M1011_g
+ N_A_110_47#_M1017_g N_A_110_47#_M1013_g N_A_110_47#_M1018_g
+ N_A_110_47#_M1014_g N_A_110_47#_M1020_g N_A_110_47#_M1016_g
+ N_A_110_47#_M1023_g N_A_110_47#_M1024_g N_A_110_47#_M1029_g
+ N_A_110_47#_M1025_g N_A_110_47#_M1031_g N_A_110_47#_M1027_g
+ N_A_110_47#_M1032_g N_A_110_47#_M1028_g N_A_110_47#_M1033_g
+ N_A_110_47#_M1030_g N_A_110_47#_M1036_g N_A_110_47#_M1034_g
+ N_A_110_47#_c_201_n N_A_110_47#_M1037_g N_A_110_47#_M1035_g
+ N_A_110_47#_c_203_n N_A_110_47#_c_223_n N_A_110_47#_c_236_n
+ N_A_110_47#_c_204_n N_A_110_47#_c_224_n N_A_110_47#_c_205_n
+ N_A_110_47#_c_244_n N_A_110_47#_c_246_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%A_110_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%KAPWR N_KAPWR_M1009_d
+ N_KAPWR_M1019_d N_KAPWR_M1038_d N_KAPWR_M1001_s N_KAPWR_M1006_s
+ N_KAPWR_M1011_s N_KAPWR_M1014_s N_KAPWR_M1024_s N_KAPWR_M1027_s
+ N_KAPWR_M1030_s N_KAPWR_M1035_s N_KAPWR_c_521_n N_KAPWR_c_522_n
+ N_KAPWR_c_525_n N_KAPWR_c_541_n N_KAPWR_c_527_n N_KAPWR_c_545_n
+ N_KAPWR_c_546_n N_KAPWR_c_548_n N_KAPWR_c_550_n N_KAPWR_c_551_n
+ N_KAPWR_c_553_n N_KAPWR_c_555_n N_KAPWR_c_556_n N_KAPWR_c_558_n
+ N_KAPWR_c_560_n N_KAPWR_c_561_n N_KAPWR_c_563_n N_KAPWR_c_565_n
+ N_KAPWR_c_567_n N_KAPWR_c_569_n N_KAPWR_c_571_n N_KAPWR_c_572_n
+ N_KAPWR_c_574_n N_KAPWR_c_576_n N_KAPWR_c_578_n N_KAPWR_c_581_n
+ N_KAPWR_c_583_n N_KAPWR_c_523_n KAPWR N_KAPWR_c_524_n N_KAPWR_c_532_n
+ N_KAPWR_c_535_n KAPWR PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%X N_X_M1002_s N_X_M1004_s
+ N_X_M1008_s N_X_M1017_s N_X_M1020_s N_X_M1029_s N_X_M1032_s N_X_M1036_s
+ N_X_M1000_d N_X_M1005_d N_X_M1010_d N_X_M1013_d N_X_M1016_d N_X_M1025_d
+ N_X_M1028_d N_X_M1034_d N_X_c_719_n N_X_c_720_n N_X_c_721_n N_X_c_755_n
+ N_X_c_722_n N_X_c_723_n N_X_c_765_n N_X_c_724_n N_X_c_725_n N_X_c_775_n
+ N_X_c_726_n N_X_c_727_n N_X_c_786_n N_X_c_728_n N_X_c_729_n N_X_c_796_n
+ N_X_c_730_n N_X_c_731_n N_X_c_806_n N_X_c_732_n N_X_c_733_n N_X_c_734_n
+ N_X_c_816_n N_X_c_735_n N_X_c_822_n N_X_c_736_n N_X_c_828_n N_X_c_737_n
+ N_X_c_835_n N_X_c_738_n N_X_c_842_n N_X_c_739_n N_X_c_848_n N_X_c_740_n X X X
+ X N_X_c_743_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%X
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VGND N_VGND_M1012_s N_VGND_M1022_s
+ N_VGND_M1039_s N_VGND_M1003_d N_VGND_M1007_d N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1023_d N_VGND_M1031_d N_VGND_M1033_d N_VGND_M1037_d N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n
+ N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n N_VGND_c_1031_n
+ N_VGND_c_1032_n N_VGND_c_1033_n N_VGND_c_1034_n N_VGND_c_1035_n
+ N_VGND_c_1036_n N_VGND_c_1037_n N_VGND_c_1038_n N_VGND_c_1039_n
+ N_VGND_c_1040_n N_VGND_c_1041_n N_VGND_c_1042_n N_VGND_c_1043_n VGND
+ N_VGND_c_1044_n N_VGND_c_1045_n N_VGND_c_1046_n N_VGND_c_1047_n
+ N_VGND_c_1048_n N_VGND_c_1049_n N_VGND_c_1050_n N_VGND_c_1051_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VPWR VPWR N_VPWR_c_1180_n
+ N_VPWR_c_1179_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_16%VPWR
cc_1 VNB N_A_M1012_g 0.0293912f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_M1022_g 0.0229781f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_3 VNB N_A_M1026_g 0.0229774f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.445
cc_4 VNB N_A_M1039_g 0.0234436f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.445
cc_5 VNB A 0.0236658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_123_n 0.109553f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.155
cc_7 VNB N_A_110_47#_M1002_g 0.0260664f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.9
cc_8 VNB N_A_110_47#_M1003_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.445
cc_9 VNB N_A_110_47#_M1004_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_110_47#_M1007_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.155
cc_11 VNB N_A_110_47#_M1008_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_110_47#_M1015_g 0.0241428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1017_g 0.0238169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_M1018_g 0.0240545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_M1020_g 0.0240466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_110_47#_M1023_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_110_47#_M1029_g 0.0241355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_110_47#_M1031_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_110_47#_M1032_g 0.0241328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_110_47#_M1033_g 0.0241116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_110_47#_M1036_g 0.0237673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_110_47#_c_201_n 0.300055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_110_47#_M1037_g 0.0320587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_110_47#_c_203_n 0.00436501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_110_47#_c_204_n 0.00481736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_110_47#_c_205_n 0.00429043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_719_n 0.00160391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_720_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_721_n 0.00419804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_722_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_723_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_724_n 0.00125415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_725_n 0.00501892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_726_n 6.22964e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_727_n 0.00491776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_728_n 0.00125437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_729_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_730_n 0.00126258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_731_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_732_n 0.00126798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_733_n 4.84646e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_734_n 0.00137779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_735_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_736_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_737_n 0.00217463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_X_c_738_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_739_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_740_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB X 0.0318745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_1019_n 0.0107531f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_51 VNB N_VGND_c_1020_n 0.0190761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_1021_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.155
cc_53 VNB N_VGND_c_1022_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1023_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1024_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1025_n 0.00390627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1026_n 0.0157899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1027_n 0.00395785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1028_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1029_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1030_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1031_n 0.00402207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1032_n 0.0135264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1033_n 0.0178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1034_n 0.0167416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1035_n 0.00500104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1036_n 0.0160902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1037_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1038_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1039_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1040_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1041_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1042_n 0.0157075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1043_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1044_n 0.0169722f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1045_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1046_n 0.0154599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1047_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1048_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1049_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1050_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1051_n 0.430355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VPWR_c_1179_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_84 VPB N_A_c_124_n 0.0192412f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.41
cc_85 VPB N_A_c_125_n 0.0143984f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.41
cc_86 VPB N_A_c_126_n 0.0143984f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.41
cc_87 VPB N_A_c_127_n 0.0145807f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.41
cc_88 VPB A 0.00122297f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_89 VPB N_A_c_123_n 0.0418698f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.155
cc_90 VPB N_A_110_47#_M1000_g 0.0190636f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.41
cc_91 VPB N_A_110_47#_M1001_g 0.0187483f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_92 VPB N_A_110_47#_M1005_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_93 VPB N_A_110_47#_M1006_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_110_47#_M1010_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_110_47#_M1011_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_110_47#_M1013_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_110_47#_M1014_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_110_47#_M1016_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_110_47#_M1024_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_110_47#_M1025_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_110_47#_M1027_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_110_47#_M1028_g 0.0187387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_110_47#_M1030_g 0.0186963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_110_47#_M1034_g 0.0173762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_110_47#_c_201_n 0.0522358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_110_47#_M1035_g 0.0224494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_110_47#_c_223_n 0.00131518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_110_47#_c_224_n 0.00131518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_110_47#_c_205_n 0.00258437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_KAPWR_c_521_n 0.00916947f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_111 VPB N_KAPWR_c_522_n 0.0124499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_KAPWR_c_523_n 0.0178729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_KAPWR_c_524_n 0.0332027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB X 0.0102708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_X_c_743_n 0.00990633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_1180_n 0.245418f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.9
cc_117 VPB N_VPWR_c_1179_n 0.0439056f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=0.445
cc_118 N_A_M1039_g N_A_110_47#_M1002_g 0.0178631f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_c_127_n N_A_110_47#_M1000_g 0.0178631f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_123_n N_A_110_47#_c_201_n 0.0178631f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_121 N_A_M1012_g N_A_110_47#_c_203_n 0.00388687f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_M1022_g N_A_110_47#_c_203_n 0.00353563f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_123 A N_A_110_47#_c_203_n 0.0212325f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_124 N_A_c_123_n N_A_110_47#_c_203_n 0.0132823f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_125 N_A_c_124_n N_A_110_47#_c_223_n 0.00207315f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_125_n N_A_110_47#_c_223_n 0.00124674f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_123_n N_A_110_47#_c_223_n 0.00991177f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_128 N_A_c_123_n N_A_110_47#_c_236_n 0.0527608f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_129 N_A_M1026_g N_A_110_47#_c_204_n 0.00352135f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_M1039_g N_A_110_47#_c_204_n 0.00356184f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_c_123_n N_A_110_47#_c_204_n 0.0139367f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_132 N_A_c_126_n N_A_110_47#_c_224_n 0.00124674f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_127_n N_A_110_47#_c_224_n 0.00207315f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_123_n N_A_110_47#_c_224_n 0.00774413f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_135 N_A_c_123_n N_A_110_47#_c_205_n 0.0206088f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_136 A N_A_110_47#_c_244_n 0.0178087f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_137 N_A_c_123_n N_A_110_47#_c_244_n 0.010956f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_138 N_A_c_123_n N_A_110_47#_c_246_n 0.00889636f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_139 N_A_c_124_n N_KAPWR_c_525_n 0.00604839f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_125_n N_KAPWR_c_525_n 0.00604839f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_126_n N_KAPWR_c_527_n 0.00604839f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_127_n N_KAPWR_c_527_n 0.00604839f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_124_n N_KAPWR_c_524_n 0.0105462f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_144 A N_KAPWR_c_524_n 0.0236933f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_145 N_A_c_123_n N_KAPWR_c_524_n 0.00809407f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_146 N_A_c_125_n N_KAPWR_c_532_n 0.00968558f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_126_n N_KAPWR_c_532_n 0.00972223f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_123_n N_KAPWR_c_532_n 0.00281536f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_149 N_A_c_127_n N_KAPWR_c_535_n 0.0097223f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_M1012_g N_VGND_c_1020_n 0.0038241f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_151 A N_VGND_c_1020_n 0.0245931f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_152 N_A_c_123_n N_VGND_c_1020_n 0.00149294f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_153 N_A_M1022_g N_VGND_c_1021_n 0.00168046f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_M1026_g N_VGND_c_1021_n 0.00168046f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_c_123_n N_VGND_c_1021_n 0.00255763f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_156 N_A_M1039_g N_VGND_c_1022_n 0.00170359f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_M1026_g N_VGND_c_1034_n 0.00585385f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_M1039_g N_VGND_c_1034_n 0.00585385f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_M1012_g N_VGND_c_1044_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_M1022_g N_VGND_c_1044_n 0.00585385f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_M1012_g N_VGND_c_1051_n 0.011499f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_M1022_g N_VGND_c_1051_n 0.010643f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_M1026_g N_VGND_c_1051_n 0.010643f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_M1039_g N_VGND_c_1051_n 0.0106694f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_165 A N_VGND_c_1051_n 0.00157507f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A_c_124_n N_VPWR_c_1180_n 0.0054895f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_125_n N_VPWR_c_1180_n 0.0054895f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_126_n N_VPWR_c_1180_n 0.0054895f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_127_n N_VPWR_c_1180_n 0.0054895f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_124_n N_VPWR_c_1179_n 0.00605725f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_125_n N_VPWR_c_1179_n 0.00512464f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_126_n N_VPWR_c_1179_n 0.00512464f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_127_n N_VPWR_c_1179_n 0.00514998f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_110_47#_c_223_n N_KAPWR_c_521_n 4.33193e-19 $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_175 N_A_110_47#_M1034_g N_KAPWR_c_522_n 0.00272513f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_176 N_A_110_47#_M1035_g N_KAPWR_c_522_n 0.0023812f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A_110_47#_M1009_s N_KAPWR_c_525_n 0.00380222f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_110_47#_c_223_n N_KAPWR_c_525_n 0.0200676f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_179 N_A_110_47#_c_223_n N_KAPWR_c_541_n 4.33193e-19 $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_180 N_A_110_47#_c_224_n N_KAPWR_c_541_n 4.33193e-19 $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_181 N_A_110_47#_M1021_s N_KAPWR_c_527_n 0.00380222f $X=1.41 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A_110_47#_c_224_n N_KAPWR_c_527_n 0.0200378f $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_183 N_A_110_47#_c_224_n N_KAPWR_c_545_n 4.39484e-19 $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_184 N_A_110_47#_M1001_g N_KAPWR_c_546_n 0.00114528f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_110_47#_M1005_g N_KAPWR_c_546_n 0.00114528f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_110_47#_M1000_g N_KAPWR_c_548_n 0.00604839f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_110_47#_M1001_g N_KAPWR_c_548_n 0.00233003f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_110_47#_M1001_g N_KAPWR_c_550_n 6.91139e-19 $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_110_47#_M1006_g N_KAPWR_c_551_n 0.00115346f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_110_47#_M1010_g N_KAPWR_c_551_n 0.00115346f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_110_47#_M1005_g N_KAPWR_c_553_n 0.0026941f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_110_47#_M1006_g N_KAPWR_c_553_n 0.0026941f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_110_47#_M1010_g N_KAPWR_c_555_n 6.44793e-19 $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_110_47#_M1011_g N_KAPWR_c_556_n 0.00115346f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_110_47#_M1013_g N_KAPWR_c_556_n 0.00115346f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_110_47#_M1010_g N_KAPWR_c_558_n 0.00251207f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_110_47#_M1011_g N_KAPWR_c_558_n 0.0026941f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_198 N_A_110_47#_M1013_g N_KAPWR_c_560_n 6.44793e-19 $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_110_47#_M1014_g N_KAPWR_c_561_n 0.00113845f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_110_47#_M1016_g N_KAPWR_c_561_n 0.00111208f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_110_47#_M1013_g N_KAPWR_c_563_n 0.00251207f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_110_47#_M1014_g N_KAPWR_c_563_n 0.00260308f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_110_47#_M1014_g N_KAPWR_c_565_n 4.8879e-19 $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_110_47#_M1016_g N_KAPWR_c_565_n 6.40226e-19 $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_110_47#_M1024_g N_KAPWR_c_567_n 0.00116608f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_110_47#_M1025_g N_KAPWR_c_567_n 0.00112416f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_110_47#_M1016_g N_KAPWR_c_569_n 0.00251207f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_110_47#_M1024_g N_KAPWR_c_569_n 0.0026941f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_110_47#_M1025_g N_KAPWR_c_571_n 6.40226e-19 $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_110_47#_M1027_g N_KAPWR_c_572_n 0.00116608f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_110_47#_M1028_g N_KAPWR_c_572_n 0.00112416f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_110_47#_M1025_g N_KAPWR_c_574_n 0.00251207f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_110_47#_M1027_g N_KAPWR_c_574_n 0.00260308f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_110_47#_M1027_g N_KAPWR_c_576_n 4.93728e-19 $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_110_47#_M1028_g N_KAPWR_c_576_n 3.61486e-19 $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_110_47#_M1030_g N_KAPWR_c_578_n 0.00116801f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_110_47#_M1034_g N_KAPWR_c_578_n 0.00115258f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_110_47#_c_201_n N_KAPWR_c_578_n 3.46041e-19 $X=8.64 $Y=0.95 $X2=0
+ $Y2=0
cc_219 N_A_110_47#_M1028_g N_KAPWR_c_581_n 0.00260308f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_110_47#_M1030_g N_KAPWR_c_581_n 0.00244893f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_110_47#_M1030_g N_KAPWR_c_583_n 6.11058e-19 $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_110_47#_M1035_g N_KAPWR_c_523_n 0.00394183f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_110_47#_c_223_n N_KAPWR_c_524_n 0.0388243f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_224 N_A_110_47#_c_223_n N_KAPWR_c_532_n 0.0388243f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_225 N_A_110_47#_c_236_n N_KAPWR_c_532_n 0.0212385f $X=1.43 $Y=1.2 $X2=0 $Y2=0
cc_226 N_A_110_47#_c_224_n N_KAPWR_c_532_n 0.0386342f $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_227 N_A_110_47#_M1000_g N_KAPWR_c_535_n 0.00962434f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_110_47#_c_224_n N_KAPWR_c_535_n 0.0386367f $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_229 N_A_110_47#_c_205_n N_KAPWR_c_535_n 0.0223469f $X=7.505 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_110_47#_M1002_g N_X_c_719_n 0.00120255f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_110_47#_M1003_g N_X_c_719_n 0.00120255f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A_110_47#_c_204_n N_X_c_719_n 0.00257148f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A_110_47#_M1003_g N_X_c_720_n 0.0119364f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A_110_47#_M1004_g N_X_c_720_n 0.0122327f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_235 N_A_110_47#_c_201_n N_X_c_720_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_236 N_A_110_47#_c_205_n N_X_c_720_n 0.0429599f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_110_47#_M1002_g N_X_c_721_n 0.00289158f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_238 N_A_110_47#_c_201_n N_X_c_721_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_239 N_A_110_47#_c_204_n N_X_c_721_n 0.00599637f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A_110_47#_c_205_n N_X_c_721_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_110_47#_M1001_g N_X_c_755_n 0.0113432f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_110_47#_M1005_g N_X_c_755_n 0.0113034f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_243 N_A_110_47#_c_201_n N_X_c_755_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_244 N_A_110_47#_c_205_n N_X_c_755_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_110_47#_M1004_g N_X_c_722_n 0.00120255f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_246 N_A_110_47#_M1007_g N_X_c_722_n 0.00120255f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_247 N_A_110_47#_M1007_g N_X_c_723_n 0.0122792f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_248 N_A_110_47#_M1008_g N_X_c_723_n 0.0122792f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A_110_47#_c_201_n N_X_c_723_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_250 N_A_110_47#_c_205_n N_X_c_723_n 0.0429599f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_110_47#_M1006_g N_X_c_765_n 0.0113694f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_110_47#_M1010_g N_X_c_765_n 0.0113563f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_253 N_A_110_47#_c_201_n N_X_c_765_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_254 N_A_110_47#_c_205_n N_X_c_765_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_110_47#_M1008_g N_X_c_724_n 0.00120255f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_256 N_A_110_47#_M1015_g N_X_c_724_n 0.00118828f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_257 N_A_110_47#_M1015_g N_X_c_725_n 0.0122792f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A_110_47#_M1017_g N_X_c_725_n 0.00994201f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_110_47#_c_201_n N_X_c_725_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_260 N_A_110_47#_c_205_n N_X_c_725_n 0.0418783f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_110_47#_M1011_g N_X_c_775_n 0.0113694f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_110_47#_M1013_g N_X_c_775_n 0.0113007f $X=4.775 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_110_47#_c_201_n N_X_c_775_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_264 N_A_110_47#_c_205_n N_X_c_775_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_110_47#_M1015_g N_X_c_726_n 5.05907e-19 $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_266 N_A_110_47#_M1017_g N_X_c_726_n 0.0062908f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_267 N_A_110_47#_M1018_g N_X_c_726_n 0.00119799f $X=5.205 $Y=0.445 $X2=0 $Y2=0
cc_268 N_A_110_47#_M1018_g N_X_c_727_n 0.0122482f $X=5.205 $Y=0.445 $X2=0 $Y2=0
cc_269 N_A_110_47#_M1020_g N_X_c_727_n 0.0101865f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_110_47#_c_201_n N_X_c_727_n 0.00253724f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_271 N_A_110_47#_c_205_n N_X_c_727_n 0.0418596f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_110_47#_M1014_g N_X_c_786_n 0.0113189f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_110_47#_M1016_g N_X_c_786_n 0.0113123f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_110_47#_c_201_n N_X_c_786_n 0.00220405f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_275 N_A_110_47#_c_205_n N_X_c_786_n 0.0378421f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_110_47#_M1020_g N_X_c_728_n 0.00121272f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A_110_47#_M1023_g N_X_c_728_n 0.00117849f $X=6.06 $Y=0.445 $X2=0 $Y2=0
cc_278 N_A_110_47#_M1023_g N_X_c_729_n 0.0122792f $X=6.06 $Y=0.445 $X2=0 $Y2=0
cc_279 N_A_110_47#_M1029_g N_X_c_729_n 0.0102175f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_110_47#_c_201_n N_X_c_729_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_281 N_A_110_47#_c_205_n N_X_c_729_n 0.0429636f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_110_47#_M1024_g N_X_c_796_n 0.0113694f $X=6.06 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_110_47#_M1025_g N_X_c_796_n 0.0113563f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_110_47#_c_201_n N_X_c_796_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_285 N_A_110_47#_c_205_n N_X_c_796_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_110_47#_M1029_g N_X_c_730_n 0.00122723f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_287 N_A_110_47#_M1031_g N_X_c_730_n 0.00117849f $X=6.92 $Y=0.445 $X2=0 $Y2=0
cc_288 N_A_110_47#_M1031_g N_X_c_731_n 0.0122792f $X=6.92 $Y=0.445 $X2=0 $Y2=0
cc_289 N_A_110_47#_M1032_g N_X_c_731_n 0.0102175f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_290 N_A_110_47#_c_201_n N_X_c_731_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_291 N_A_110_47#_c_205_n N_X_c_731_n 0.0429636f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_110_47#_M1027_g N_X_c_806_n 0.011359f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A_110_47#_M1028_g N_X_c_806_n 0.0113628f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A_110_47#_c_201_n N_X_c_806_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_295 N_A_110_47#_c_205_n N_X_c_806_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_110_47#_M1032_g N_X_c_732_n 0.00122723f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_110_47#_M1033_g N_X_c_732_n 0.00118774f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_110_47#_M1033_g N_X_c_733_n 0.0141891f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_299 N_A_110_47#_c_205_n N_X_c_733_n 3.30399e-19 $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_110_47#_M1036_g N_X_c_734_n 0.00121196f $X=8.21 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_110_47#_M1037_g N_X_c_734_n 0.00221636f $X=8.64 $Y=0.445 $X2=0 $Y2=0
cc_302 N_A_110_47#_M1000_g N_X_c_816_n 0.00130422f $X=2.195 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A_110_47#_M1001_g N_X_c_816_n 0.00140908f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A_110_47#_c_201_n N_X_c_816_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_305 N_A_110_47#_c_205_n N_X_c_816_n 0.0155795f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_110_47#_c_201_n N_X_c_735_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_307 N_A_110_47#_c_205_n N_X_c_735_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A_110_47#_M1005_g N_X_c_822_n 0.00141407f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_110_47#_M1006_g N_X_c_822_n 0.00141558f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_310 N_A_110_47#_c_201_n N_X_c_822_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_311 N_A_110_47#_c_205_n N_X_c_822_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_110_47#_c_201_n N_X_c_736_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_313 N_A_110_47#_c_205_n N_X_c_736_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_110_47#_M1010_g N_X_c_828_n 0.00141558f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A_110_47#_M1011_g N_X_c_828_n 0.00141558f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_110_47#_c_201_n N_X_c_828_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_317 N_A_110_47#_c_205_n N_X_c_828_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_110_47#_M1017_g N_X_c_737_n 0.00211052f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_319 N_A_110_47#_c_201_n N_X_c_737_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_320 N_A_110_47#_c_205_n N_X_c_737_n 0.0225791f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_110_47#_M1013_g N_X_c_835_n 0.00141558f $X=4.775 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_110_47#_M1014_g N_X_c_835_n 0.00141558f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_110_47#_c_201_n N_X_c_835_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_324 N_A_110_47#_c_205_n N_X_c_835_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_110_47#_M1020_g N_X_c_738_n 0.00203048f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_326 N_A_110_47#_c_201_n N_X_c_738_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_327 N_A_110_47#_c_205_n N_X_c_738_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_110_47#_M1024_g N_X_c_842_n 0.00140594f $X=6.06 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_110_47#_c_201_n N_X_c_842_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_330 N_A_110_47#_c_205_n N_X_c_842_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_110_47#_M1029_g N_X_c_739_n 0.00203048f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_332 N_A_110_47#_c_201_n N_X_c_739_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_333 N_A_110_47#_c_205_n N_X_c_739_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_110_47#_M1027_g N_X_c_848_n 0.00140594f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_110_47#_c_201_n N_X_c_848_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_336 N_A_110_47#_c_205_n N_X_c_848_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_110_47#_M1032_g N_X_c_740_n 0.00203048f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_110_47#_c_201_n N_X_c_740_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_339 N_A_110_47#_c_205_n N_X_c_740_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_110_47#_M1033_g X 0.00147955f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_341 N_A_110_47#_M1030_g X 0.00539328f $X=7.78 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_110_47#_M1036_g X 0.011848f $X=8.21 $Y=0.445 $X2=0 $Y2=0
cc_343 N_A_110_47#_M1034_g X 0.00593452f $X=8.21 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_110_47#_c_201_n X 0.0567372f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_345 N_A_110_47#_M1037_g X 0.0136957f $X=8.64 $Y=0.445 $X2=0 $Y2=0
cc_346 N_A_110_47#_M1035_g X 0.00761986f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A_110_47#_c_205_n X 0.0208936f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A_110_47#_M1030_g N_X_c_743_n 0.0143099f $X=7.78 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A_110_47#_M1034_g N_X_c_743_n 0.0108311f $X=8.21 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A_110_47#_c_201_n N_X_c_743_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_351 N_A_110_47#_M1035_g N_X_c_743_n 0.0256934f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A_110_47#_c_205_n N_X_c_743_n 0.0170247f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A_110_47#_c_236_n N_VGND_c_1021_n 0.00764914f $X=1.43 $Y=1.2 $X2=0
+ $Y2=0
cc_354 N_A_110_47#_M1002_g N_VGND_c_1022_n 0.00170359f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_355 N_A_110_47#_c_205_n N_VGND_c_1022_n 0.0091835f $X=7.505 $Y=1.16 $X2=0
+ $Y2=0
cc_356 N_A_110_47#_M1003_g N_VGND_c_1023_n 0.00161372f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_357 N_A_110_47#_M1004_g N_VGND_c_1023_n 0.00161372f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_110_47#_M1007_g N_VGND_c_1024_n 0.00161372f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_A_110_47#_M1008_g N_VGND_c_1024_n 0.00161372f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_A_110_47#_M1015_g N_VGND_c_1025_n 0.00160579f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_A_110_47#_M1017_g N_VGND_c_1025_n 0.0015619f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_A_110_47#_M1017_g N_VGND_c_1026_n 0.00438144f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_110_47#_M1018_g N_VGND_c_1026_n 0.00439206f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_A_110_47#_M1018_g N_VGND_c_1027_n 0.00161724f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_365 N_A_110_47#_M1020_g N_VGND_c_1027_n 0.00156827f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_110_47#_M1020_g N_VGND_c_1028_n 0.00439206f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_367 N_A_110_47#_M1023_g N_VGND_c_1028_n 0.00439206f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_368 N_A_110_47#_M1023_g N_VGND_c_1029_n 0.00162174f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_369 N_A_110_47#_M1029_g N_VGND_c_1029_n 0.00157905f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_370 N_A_110_47#_M1031_g N_VGND_c_1030_n 0.00162174f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_110_47#_M1032_g N_VGND_c_1030_n 0.00157905f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_110_47#_M1033_g N_VGND_c_1031_n 0.00162705f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_373 N_A_110_47#_M1036_g N_VGND_c_1031_n 0.00161372f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_110_47#_c_201_n N_VGND_c_1031_n 4.7914e-19 $X=8.64 $Y=0.95 $X2=0
+ $Y2=0
cc_375 N_A_110_47#_M1037_g N_VGND_c_1033_n 0.00341923f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_110_47#_c_204_n N_VGND_c_1034_n 0.0137163f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_110_47#_M1002_g N_VGND_c_1036_n 0.00585385f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_110_47#_M1003_g N_VGND_c_1036_n 0.00439206f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_110_47#_M1004_g N_VGND_c_1038_n 0.00439206f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_380 N_A_110_47#_M1007_g N_VGND_c_1038_n 0.00439206f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_381 N_A_110_47#_M1008_g N_VGND_c_1040_n 0.00439206f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_A_110_47#_M1015_g N_VGND_c_1040_n 0.00439206f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_110_47#_M1032_g N_VGND_c_1042_n 0.00439206f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_384 N_A_110_47#_M1033_g N_VGND_c_1042_n 0.00439206f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_110_47#_c_203_n N_VGND_c_1044_n 0.0128787f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_110_47#_M1029_g N_VGND_c_1045_n 0.00439206f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_110_47#_M1031_g N_VGND_c_1045_n 0.00439206f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_110_47#_M1036_g N_VGND_c_1046_n 0.00439071f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_389 N_A_110_47#_M1037_g N_VGND_c_1046_n 0.00439071f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_110_47#_M1012_d N_VGND_c_1051_n 0.00422994f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_391 N_A_110_47#_M1026_d N_VGND_c_1051_n 0.00336236f $X=1.41 $Y=0.235 $X2=0
+ $Y2=0
cc_392 N_A_110_47#_M1002_g N_VGND_c_1051_n 0.0106694f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_393 N_A_110_47#_M1003_g N_VGND_c_1051_n 0.00590932f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_394 N_A_110_47#_M1004_g N_VGND_c_1051_n 0.00590932f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_110_47#_M1007_g N_VGND_c_1051_n 0.00590932f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_A_110_47#_M1008_g N_VGND_c_1051_n 0.00590932f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_A_110_47#_M1015_g N_VGND_c_1051_n 0.00590932f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_110_47#_M1017_g N_VGND_c_1051_n 0.00587292f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_399 N_A_110_47#_M1018_g N_VGND_c_1051_n 0.00589619f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_400 N_A_110_47#_M1020_g N_VGND_c_1051_n 0.00592128f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_110_47#_M1023_g N_VGND_c_1051_n 0.00590932f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_402 N_A_110_47#_M1029_g N_VGND_c_1051_n 0.00593441f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_403 N_A_110_47#_M1031_g N_VGND_c_1051_n 0.00590932f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_110_47#_M1032_g N_VGND_c_1051_n 0.00593441f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_405 N_A_110_47#_M1033_g N_VGND_c_1051_n 0.00590932f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_406 N_A_110_47#_M1036_g N_VGND_c_1051_n 0.00590684f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_407 N_A_110_47#_M1037_g N_VGND_c_1051_n 0.00691049f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_408 N_A_110_47#_c_203_n N_VGND_c_1051_n 0.00854752f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_409 N_A_110_47#_c_204_n N_VGND_c_1051_n 0.00950576f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_110_47#_M1000_g N_VPWR_c_1180_n 0.0054895f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_411 N_A_110_47#_M1001_g N_VPWR_c_1180_n 0.00585385f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_110_47#_M1005_g N_VPWR_c_1180_n 0.00585385f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_413 N_A_110_47#_M1006_g N_VPWR_c_1180_n 0.00585385f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_414 N_A_110_47#_M1010_g N_VPWR_c_1180_n 0.00585385f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_415 N_A_110_47#_M1011_g N_VPWR_c_1180_n 0.00585385f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_416 N_A_110_47#_M1013_g N_VPWR_c_1180_n 0.00585385f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_417 N_A_110_47#_M1014_g N_VPWR_c_1180_n 0.00585385f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_110_47#_M1016_g N_VPWR_c_1180_n 0.00585385f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_419 N_A_110_47#_M1024_g N_VPWR_c_1180_n 0.00585385f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_420 N_A_110_47#_M1025_g N_VPWR_c_1180_n 0.00585385f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_421 N_A_110_47#_M1027_g N_VPWR_c_1180_n 0.00585385f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_422 N_A_110_47#_M1028_g N_VPWR_c_1180_n 0.00585385f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_423 N_A_110_47#_M1030_g N_VPWR_c_1180_n 0.00585385f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_424 N_A_110_47#_M1034_g N_VPWR_c_1180_n 0.00585385f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_425 N_A_110_47#_M1035_g N_VPWR_c_1180_n 0.00556673f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_426 N_A_110_47#_c_223_n N_VPWR_c_1180_n 0.0124538f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_427 N_A_110_47#_c_224_n N_VPWR_c_1180_n 0.0120686f $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_428 N_A_110_47#_M1009_s N_VPWR_c_1179_n 0.00149727f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_429 N_A_110_47#_M1021_s N_VPWR_c_1179_n 0.00149767f $X=1.41 $Y=1.485 $X2=0
+ $Y2=0
cc_430 N_A_110_47#_M1000_g N_VPWR_c_1179_n 0.00514998f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_A_110_47#_M1001_g N_VPWR_c_1179_n 0.00525209f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_A_110_47#_M1005_g N_VPWR_c_1179_n 0.00525209f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_A_110_47#_M1006_g N_VPWR_c_1179_n 0.00525209f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_434 N_A_110_47#_M1010_g N_VPWR_c_1179_n 0.00525209f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_435 N_A_110_47#_M1011_g N_VPWR_c_1179_n 0.00525209f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_436 N_A_110_47#_M1013_g N_VPWR_c_1179_n 0.00525209f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_437 N_A_110_47#_M1014_g N_VPWR_c_1179_n 0.00523845f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_438 N_A_110_47#_M1016_g N_VPWR_c_1179_n 0.00523845f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_439 N_A_110_47#_M1024_g N_VPWR_c_1179_n 0.00525209f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_A_110_47#_M1025_g N_VPWR_c_1179_n 0.00525209f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_441 N_A_110_47#_M1027_g N_VPWR_c_1179_n 0.00525209f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_442 N_A_110_47#_M1028_g N_VPWR_c_1179_n 0.00525209f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_443 N_A_110_47#_M1030_g N_VPWR_c_1179_n 0.00525209f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_444 N_A_110_47#_M1034_g N_VPWR_c_1179_n 0.00525209f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_445 N_A_110_47#_M1035_g N_VPWR_c_1179_n 0.00622573f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_446 N_A_110_47#_c_223_n N_VPWR_c_1179_n 0.00174489f $X=0.69 $Y=1.615 $X2=0
+ $Y2=0
cc_447 N_A_110_47#_c_224_n N_VPWR_c_1179_n 0.00175268f $X=1.55 $Y=1.615 $X2=0
+ $Y2=0
cc_448 N_KAPWR_c_548_n N_X_M1000_d 0.00202712f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_449 N_KAPWR_c_553_n N_X_M1005_d 2.52013e-19 $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_450 N_KAPWR_c_558_n N_X_M1010_d 2.52013e-19 $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_451 N_KAPWR_c_563_n N_X_M1013_d 2.52013e-19 $X=5.275 $Y=2.21 $X2=0 $Y2=0
cc_452 N_KAPWR_c_569_n N_X_M1016_d 2.83515e-19 $X=6.135 $Y=2.21 $X2=0 $Y2=0
cc_453 N_KAPWR_c_574_n N_X_M1025_d 2.83515e-19 $X=6.99 $Y=2.21 $X2=0 $Y2=0
cc_454 N_KAPWR_c_581_n N_X_M1028_d 2.86889e-19 $X=7.84 $Y=2.21 $X2=0 $Y2=0
cc_455 N_KAPWR_M1001_s N_X_c_755_n 0.00325883f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_456 N_KAPWR_c_546_n N_X_c_755_n 0.0127908f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_457 N_KAPWR_c_548_n N_X_c_755_n 0.00434646f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_458 N_KAPWR_c_550_n N_X_c_755_n 0.0023936f $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_459 N_KAPWR_c_553_n N_X_c_755_n 0.00532372f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_460 N_KAPWR_M1006_s N_X_c_765_n 0.00325489f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_461 N_KAPWR_c_551_n N_X_c_765_n 0.0128604f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_462 N_KAPWR_c_553_n N_X_c_765_n 0.00497471f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_463 N_KAPWR_c_555_n N_X_c_765_n 0.00245411f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_464 N_KAPWR_c_558_n N_X_c_765_n 0.00466059f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_465 N_KAPWR_M1011_s N_X_c_775_n 0.00325489f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_466 N_KAPWR_c_556_n N_X_c_775_n 0.0128604f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_467 N_KAPWR_c_558_n N_X_c_775_n 0.00497471f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_468 N_KAPWR_c_560_n N_X_c_775_n 0.00245411f $X=4.71 $Y=2.21 $X2=0 $Y2=0
cc_469 N_KAPWR_c_563_n N_X_c_775_n 0.00466059f $X=5.275 $Y=2.21 $X2=0 $Y2=0
cc_470 N_KAPWR_M1014_s N_X_c_786_n 0.00316145f $X=5.28 $Y=1.485 $X2=0 $Y2=0
cc_471 N_KAPWR_c_561_n N_X_c_786_n 0.012473f $X=5.42 $Y=2.21 $X2=0 $Y2=0
cc_472 N_KAPWR_c_563_n N_X_c_786_n 0.00481765f $X=5.275 $Y=2.21 $X2=0 $Y2=0
cc_473 N_KAPWR_c_565_n N_X_c_786_n 0.00295229f $X=5.565 $Y=2.21 $X2=0 $Y2=0
cc_474 N_KAPWR_c_569_n N_X_c_786_n 0.00435093f $X=6.135 $Y=2.21 $X2=0 $Y2=0
cc_475 N_KAPWR_M1024_s N_X_c_796_n 0.00325489f $X=6.135 $Y=1.485 $X2=0 $Y2=0
cc_476 N_KAPWR_c_567_n N_X_c_796_n 0.0128604f $X=6.28 $Y=2.21 $X2=0 $Y2=0
cc_477 N_KAPWR_c_569_n N_X_c_796_n 0.00536178f $X=6.135 $Y=2.21 $X2=0 $Y2=0
cc_478 N_KAPWR_c_571_n N_X_c_796_n 0.00300711f $X=6.425 $Y=2.21 $X2=0 $Y2=0
cc_479 N_KAPWR_c_574_n N_X_c_796_n 0.00435093f $X=6.99 $Y=2.21 $X2=0 $Y2=0
cc_480 N_KAPWR_M1027_s N_X_c_806_n 0.00325489f $X=6.995 $Y=1.485 $X2=0 $Y2=0
cc_481 N_KAPWR_c_572_n N_X_c_806_n 0.0128604f $X=7.135 $Y=2.21 $X2=0 $Y2=0
cc_482 N_KAPWR_c_574_n N_X_c_806_n 0.00520471f $X=6.99 $Y=2.21 $X2=0 $Y2=0
cc_483 N_KAPWR_c_576_n N_X_c_806_n 0.00298967f $X=7.28 $Y=2.21 $X2=0 $Y2=0
cc_484 N_KAPWR_c_581_n N_X_c_806_n 0.004508f $X=7.84 $Y=2.21 $X2=0 $Y2=0
cc_485 N_KAPWR_c_545_n N_X_c_816_n 2.66244e-19 $X=2.12 $Y=2.21 $X2=0 $Y2=0
cc_486 N_KAPWR_c_546_n N_X_c_816_n 0.00825548f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_487 N_KAPWR_c_548_n N_X_c_816_n 0.0230251f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_488 N_KAPWR_c_550_n N_X_c_816_n 6.89844e-19 $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_489 N_KAPWR_c_535_n N_X_c_816_n 0.0296427f $X=1.98 $Y=1.66 $X2=0 $Y2=0
cc_490 N_KAPWR_c_546_n N_X_c_822_n 0.0082718f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_491 N_KAPWR_c_550_n N_X_c_822_n 4.70067e-19 $X=2.97 $Y=2.21 $X2=0 $Y2=0
cc_492 N_KAPWR_c_551_n N_X_c_822_n 0.00822181f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_493 N_KAPWR_c_553_n N_X_c_822_n 0.0260214f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_494 N_KAPWR_c_555_n N_X_c_822_n 0.00175189f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_495 N_KAPWR_c_551_n N_X_c_828_n 0.00822181f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_496 N_KAPWR_c_555_n N_X_c_828_n 0.00153797f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_497 N_KAPWR_c_556_n N_X_c_828_n 0.00822181f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_498 N_KAPWR_c_558_n N_X_c_828_n 0.0260313f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_499 N_KAPWR_c_560_n N_X_c_828_n 0.00175189f $X=4.71 $Y=2.21 $X2=0 $Y2=0
cc_500 N_KAPWR_c_556_n N_X_c_835_n 0.00822181f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_501 N_KAPWR_c_560_n N_X_c_835_n 0.00153797f $X=4.71 $Y=2.21 $X2=0 $Y2=0
cc_502 N_KAPWR_c_561_n N_X_c_835_n 0.00821313f $X=5.42 $Y=2.21 $X2=0 $Y2=0
cc_503 N_KAPWR_c_563_n N_X_c_835_n 0.0260313f $X=5.275 $Y=2.21 $X2=0 $Y2=0
cc_504 N_KAPWR_c_565_n N_X_c_835_n 0.00152822f $X=5.565 $Y=2.21 $X2=0 $Y2=0
cc_505 N_KAPWR_c_561_n N_X_c_842_n 0.0178876f $X=5.42 $Y=2.21 $X2=0 $Y2=0
cc_506 N_KAPWR_c_565_n N_X_c_842_n 0.00155772f $X=5.565 $Y=2.21 $X2=0 $Y2=0
cc_507 N_KAPWR_c_567_n N_X_c_842_n 0.00755072f $X=6.28 $Y=2.21 $X2=0 $Y2=0
cc_508 N_KAPWR_c_569_n N_X_c_842_n 0.0261776f $X=6.135 $Y=2.21 $X2=0 $Y2=0
cc_509 N_KAPWR_c_571_n N_X_c_842_n 0.00174799f $X=6.425 $Y=2.21 $X2=0 $Y2=0
cc_510 N_KAPWR_c_567_n N_X_c_848_n 0.0178876f $X=6.28 $Y=2.21 $X2=0 $Y2=0
cc_511 N_KAPWR_c_571_n N_X_c_848_n 0.00155772f $X=6.425 $Y=2.21 $X2=0 $Y2=0
cc_512 N_KAPWR_c_572_n N_X_c_848_n 0.00755072f $X=7.135 $Y=2.21 $X2=0 $Y2=0
cc_513 N_KAPWR_c_574_n N_X_c_848_n 0.0261776f $X=6.99 $Y=2.21 $X2=0 $Y2=0
cc_514 N_KAPWR_c_576_n N_X_c_848_n 0.00152454f $X=7.28 $Y=2.21 $X2=0 $Y2=0
cc_515 N_KAPWR_M1030_s N_X_c_743_n 0.00181589f $X=7.855 $Y=1.485 $X2=0 $Y2=0
cc_516 N_KAPWR_M1035_s N_X_c_743_n 0.00325733f $X=8.715 $Y=1.485 $X2=0 $Y2=0
cc_517 N_KAPWR_c_522_n N_X_c_743_n 0.043721f $X=8.72 $Y=2.24 $X2=0 $Y2=0
cc_518 N_KAPWR_c_572_n N_X_c_743_n 0.0178903f $X=7.135 $Y=2.21 $X2=0 $Y2=0
cc_519 N_KAPWR_c_576_n N_X_c_743_n 6.89749e-19 $X=7.28 $Y=2.21 $X2=0 $Y2=0
cc_520 N_KAPWR_c_578_n N_X_c_743_n 0.0286954f $X=7.985 $Y=2.21 $X2=0 $Y2=0
cc_521 N_KAPWR_c_581_n N_X_c_743_n 0.0309849f $X=7.84 $Y=2.21 $X2=0 $Y2=0
cc_522 N_KAPWR_c_583_n N_X_c_743_n 0.00521589f $X=8.13 $Y=2.21 $X2=0 $Y2=0
cc_523 N_KAPWR_c_523_n N_X_c_743_n 0.0456665f $X=8.865 $Y=2.21 $X2=0 $Y2=0
cc_524 N_KAPWR_c_521_n N_VPWR_c_1180_n 3.60958e-19 $X=0.405 $Y=2.24 $X2=0 $Y2=0
cc_525 N_KAPWR_c_522_n N_VPWR_c_1180_n 0.00180822f $X=8.72 $Y=2.24 $X2=0 $Y2=0
cc_526 N_KAPWR_c_525_n N_VPWR_c_1180_n 0.00207669f $X=0.975 $Y=2.21 $X2=0 $Y2=0
cc_527 N_KAPWR_c_527_n N_VPWR_c_1180_n 0.00207863f $X=1.83 $Y=2.21 $X2=0 $Y2=0
cc_528 N_KAPWR_c_546_n N_VPWR_c_1180_n 0.0147484f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_529 N_KAPWR_c_548_n N_VPWR_c_1180_n 0.00186229f $X=2.68 $Y=2.21 $X2=0 $Y2=0
cc_530 N_KAPWR_c_551_n N_VPWR_c_1180_n 0.0147733f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_531 N_KAPWR_c_553_n N_VPWR_c_1180_n 0.00187059f $X=3.56 $Y=2.21 $X2=0 $Y2=0
cc_532 N_KAPWR_c_555_n N_VPWR_c_1180_n 0.00102221f $X=3.85 $Y=2.21 $X2=0 $Y2=0
cc_533 N_KAPWR_c_556_n N_VPWR_c_1180_n 0.0147733f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_534 N_KAPWR_c_558_n N_VPWR_c_1180_n 0.00102711f $X=4.42 $Y=2.21 $X2=0 $Y2=0
cc_535 N_KAPWR_c_560_n N_VPWR_c_1180_n 0.00102221f $X=4.71 $Y=2.21 $X2=0 $Y2=0
cc_536 N_KAPWR_c_561_n N_VPWR_c_1180_n 0.0140719f $X=5.42 $Y=2.21 $X2=0 $Y2=0
cc_537 N_KAPWR_c_563_n N_VPWR_c_1180_n 0.00102587f $X=5.275 $Y=2.21 $X2=0 $Y2=0
cc_538 N_KAPWR_c_565_n N_VPWR_c_1180_n 0.001017f $X=5.565 $Y=2.21 $X2=0 $Y2=0
cc_539 N_KAPWR_c_567_n N_VPWR_c_1180_n 0.0142411f $X=6.28 $Y=2.21 $X2=0 $Y2=0
cc_540 N_KAPWR_c_569_n N_VPWR_c_1180_n 0.00110732f $X=6.135 $Y=2.21 $X2=0 $Y2=0
cc_541 N_KAPWR_c_571_n N_VPWR_c_1180_n 0.001017f $X=6.425 $Y=2.21 $X2=0 $Y2=0
cc_542 N_KAPWR_c_572_n N_VPWR_c_1180_n 0.0142411f $X=7.135 $Y=2.21 $X2=0 $Y2=0
cc_543 N_KAPWR_c_574_n N_VPWR_c_1180_n 0.00110608f $X=6.99 $Y=2.21 $X2=0 $Y2=0
cc_544 N_KAPWR_c_576_n N_VPWR_c_1180_n 0.00101652f $X=7.28 $Y=2.21 $X2=0 $Y2=0
cc_545 N_KAPWR_c_578_n N_VPWR_c_1180_n 0.0145959f $X=7.985 $Y=2.21 $X2=0 $Y2=0
cc_546 N_KAPWR_c_581_n N_VPWR_c_1180_n 0.00110703f $X=7.84 $Y=2.21 $X2=0 $Y2=0
cc_547 N_KAPWR_c_583_n N_VPWR_c_1180_n 0.00101719f $X=8.13 $Y=2.21 $X2=0 $Y2=0
cc_548 N_KAPWR_c_523_n N_VPWR_c_1180_n 0.0181313f $X=8.865 $Y=2.21 $X2=0 $Y2=0
cc_549 N_KAPWR_c_524_n N_VPWR_c_1180_n 0.0210489f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_550 N_KAPWR_c_532_n N_VPWR_c_1180_n 0.0189253f $X=1.12 $Y=1.66 $X2=0 $Y2=0
cc_551 N_KAPWR_c_535_n N_VPWR_c_1180_n 0.0189253f $X=1.98 $Y=1.66 $X2=0 $Y2=0
cc_552 N_KAPWR_M1009_d N_VPWR_c_1179_n 0.00109164f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_553 N_KAPWR_M1019_d N_VPWR_c_1179_n 0.00113449f $X=0.98 $Y=1.485 $X2=0 $Y2=0
cc_554 N_KAPWR_M1038_d N_VPWR_c_1179_n 0.00113449f $X=1.84 $Y=1.485 $X2=0 $Y2=0
cc_555 N_KAPWR_M1001_s N_VPWR_c_1179_n 0.00122337f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_556 N_KAPWR_M1006_s N_VPWR_c_1179_n 0.00123133f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_557 N_KAPWR_M1011_s N_VPWR_c_1179_n 0.00123133f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_558 N_KAPWR_M1014_s N_VPWR_c_1179_n 0.00125123f $X=5.28 $Y=1.485 $X2=0 $Y2=0
cc_559 N_KAPWR_M1024_s N_VPWR_c_1179_n 0.00129179f $X=6.135 $Y=1.485 $X2=0 $Y2=0
cc_560 N_KAPWR_M1027_s N_VPWR_c_1179_n 0.00129179f $X=6.995 $Y=1.485 $X2=0 $Y2=0
cc_561 N_KAPWR_M1030_s N_VPWR_c_1179_n 0.00125148f $X=7.855 $Y=1.485 $X2=0 $Y2=0
cc_562 N_KAPWR_M1035_s N_VPWR_c_1179_n 0.00126099f $X=8.715 $Y=1.485 $X2=0 $Y2=0
cc_563 N_KAPWR_c_521_n N_VPWR_c_1179_n 0.928394f $X=0.405 $Y=2.24 $X2=0 $Y2=0
cc_564 N_KAPWR_c_546_n N_VPWR_c_1179_n 0.00236391f $X=2.825 $Y=2.21 $X2=0 $Y2=0
cc_565 N_KAPWR_c_551_n N_VPWR_c_1179_n 0.00234462f $X=3.705 $Y=2.21 $X2=0 $Y2=0
cc_566 N_KAPWR_c_556_n N_VPWR_c_1179_n 0.00234462f $X=4.565 $Y=2.21 $X2=0 $Y2=0
cc_567 N_KAPWR_c_561_n N_VPWR_c_1179_n 0.0022083f $X=5.42 $Y=2.21 $X2=0 $Y2=0
cc_568 N_KAPWR_c_567_n N_VPWR_c_1179_n 0.0022083f $X=6.28 $Y=2.21 $X2=0 $Y2=0
cc_569 N_KAPWR_c_572_n N_VPWR_c_1179_n 0.0022083f $X=7.135 $Y=2.21 $X2=0 $Y2=0
cc_570 N_KAPWR_c_578_n N_VPWR_c_1179_n 0.00229918f $X=7.985 $Y=2.21 $X2=0 $Y2=0
cc_571 N_KAPWR_c_523_n N_VPWR_c_1179_n 0.00244244f $X=8.865 $Y=2.21 $X2=0 $Y2=0
cc_572 N_KAPWR_c_524_n N_VPWR_c_1179_n 0.00300101f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_573 N_KAPWR_c_532_n N_VPWR_c_1179_n 0.00295774f $X=1.12 $Y=1.66 $X2=0 $Y2=0
cc_574 N_KAPWR_c_535_n N_VPWR_c_1179_n 0.00295774f $X=1.98 $Y=1.66 $X2=0 $Y2=0
cc_575 N_X_c_720_n N_VGND_c_1023_n 0.0164628f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_576 N_X_c_723_n N_VGND_c_1024_n 0.0164628f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_577 N_X_c_725_n N_VGND_c_1025_n 0.015936f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_578 N_X_c_725_n N_VGND_c_1026_n 0.00226107f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_579 N_X_c_726_n N_VGND_c_1026_n 0.0133875f $X=4.99 $Y=0.445 $X2=0 $Y2=0
cc_580 N_X_c_727_n N_VGND_c_1026_n 0.00224999f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_581 N_X_c_727_n N_VGND_c_1027_n 0.015713f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_582 N_X_c_727_n N_VGND_c_1028_n 0.00225184f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_583 N_X_c_728_n N_VGND_c_1028_n 0.0128416f $X=5.845 $Y=0.445 $X2=0 $Y2=0
cc_584 N_X_c_729_n N_VGND_c_1028_n 0.00239951f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_585 N_X_c_729_n N_VGND_c_1029_n 0.0161116f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_586 N_X_c_731_n N_VGND_c_1030_n 0.0161116f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_587 X N_VGND_c_1031_n 0.0186728f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_588 X N_VGND_c_1033_n 0.0243436f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_589 N_X_c_719_n N_VGND_c_1036_n 0.0128416f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_590 N_X_c_720_n N_VGND_c_1036_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_591 N_X_c_720_n N_VGND_c_1038_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_592 N_X_c_722_n N_VGND_c_1038_n 0.0128416f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_593 N_X_c_723_n N_VGND_c_1038_n 0.00224999f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_594 N_X_c_723_n N_VGND_c_1040_n 0.00224999f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_595 N_X_c_724_n N_VGND_c_1040_n 0.0128416f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_596 N_X_c_725_n N_VGND_c_1040_n 0.00224999f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_597 N_X_c_731_n N_VGND_c_1042_n 0.00225184f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_598 N_X_c_732_n N_VGND_c_1042_n 0.0128416f $X=7.565 $Y=0.445 $X2=0 $Y2=0
cc_599 N_X_c_733_n N_VGND_c_1042_n 0.00232492f $X=7.86 $Y=0.82 $X2=0 $Y2=0
cc_600 N_X_c_729_n N_VGND_c_1045_n 0.00225184f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_601 N_X_c_730_n N_VGND_c_1045_n 0.0128416f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_602 N_X_c_731_n N_VGND_c_1045_n 0.00239951f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_603 N_X_c_734_n N_VGND_c_1046_n 0.0129027f $X=8.425 $Y=0.445 $X2=0 $Y2=0
cc_604 X N_VGND_c_1046_n 0.00498855f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_605 N_X_M1002_s N_VGND_c_1051_n 0.00268444f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_606 N_X_M1004_s N_VGND_c_1051_n 0.00234574f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_607 N_X_M1008_s N_VGND_c_1051_n 0.00234574f $X=3.99 $Y=0.235 $X2=0 $Y2=0
cc_608 N_X_M1017_s N_VGND_c_1051_n 0.00230304f $X=4.85 $Y=0.235 $X2=0 $Y2=0
cc_609 N_X_M1020_s N_VGND_c_1051_n 0.00234574f $X=5.705 $Y=0.235 $X2=0 $Y2=0
cc_610 N_X_M1029_s N_VGND_c_1051_n 0.00234574f $X=6.565 $Y=0.235 $X2=0 $Y2=0
cc_611 N_X_M1032_s N_VGND_c_1051_n 0.00234574f $X=7.425 $Y=0.235 $X2=0 $Y2=0
cc_612 N_X_M1036_s N_VGND_c_1051_n 0.00234544f $X=8.285 $Y=0.235 $X2=0 $Y2=0
cc_613 N_X_c_719_n N_VGND_c_1051_n 0.00979224f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_614 N_X_c_720_n N_VGND_c_1051_n 0.00829353f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_615 N_X_c_722_n N_VGND_c_1051_n 0.00979224f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_616 N_X_c_723_n N_VGND_c_1051_n 0.00829353f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_617 N_X_c_724_n N_VGND_c_1051_n 0.00979224f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_618 N_X_c_725_n N_VGND_c_1051_n 0.0082634f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_619 N_X_c_726_n N_VGND_c_1051_n 0.0103326f $X=4.99 $Y=0.445 $X2=0 $Y2=0
cc_620 N_X_c_727_n N_VGND_c_1051_n 0.00823851f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_621 N_X_c_728_n N_VGND_c_1051_n 0.00979224f $X=5.845 $Y=0.445 $X2=0 $Y2=0
cc_622 N_X_c_729_n N_VGND_c_1051_n 0.00851943f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_623 N_X_c_730_n N_VGND_c_1051_n 0.00979224f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_624 N_X_c_731_n N_VGND_c_1051_n 0.00851943f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_625 N_X_c_732_n N_VGND_c_1051_n 0.00979224f $X=7.565 $Y=0.445 $X2=0 $Y2=0
cc_626 N_X_c_733_n N_VGND_c_1051_n 0.00379347f $X=7.86 $Y=0.82 $X2=0 $Y2=0
cc_627 N_X_c_734_n N_VGND_c_1051_n 0.00981584f $X=8.425 $Y=0.445 $X2=0 $Y2=0
cc_628 X N_VGND_c_1051_n 0.0103915f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_629 N_X_c_816_n N_VPWR_c_1180_n 0.0132747f $X=2.41 $Y=1.66 $X2=0 $Y2=0
cc_630 N_X_c_822_n N_VPWR_c_1180_n 0.0144808f $X=3.27 $Y=1.66 $X2=0 $Y2=0
cc_631 N_X_c_828_n N_VPWR_c_1180_n 0.0144808f $X=4.13 $Y=1.66 $X2=0 $Y2=0
cc_632 N_X_c_835_n N_VPWR_c_1180_n 0.0144808f $X=4.99 $Y=1.66 $X2=0 $Y2=0
cc_633 N_X_c_842_n N_VPWR_c_1180_n 0.0144808f $X=5.845 $Y=1.66 $X2=0 $Y2=0
cc_634 N_X_c_848_n N_VPWR_c_1180_n 0.0144808f $X=6.705 $Y=1.66 $X2=0 $Y2=0
cc_635 N_X_c_743_n N_VPWR_c_1180_n 0.0305634f $X=7.565 $Y=1.66 $X2=0 $Y2=0
cc_636 N_X_M1000_d N_VPWR_c_1179_n 0.00135666f $X=2.27 $Y=1.485 $X2=0 $Y2=0
cc_637 N_X_M1005_d N_VPWR_c_1179_n 0.00121566f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_638 N_X_M1010_d N_VPWR_c_1179_n 0.00121566f $X=3.99 $Y=1.485 $X2=0 $Y2=0
cc_639 N_X_M1013_d N_VPWR_c_1179_n 0.00121566f $X=4.85 $Y=1.485 $X2=0 $Y2=0
cc_640 N_X_M1016_d N_VPWR_c_1179_n 0.00121566f $X=5.705 $Y=1.485 $X2=0 $Y2=0
cc_641 N_X_M1025_d N_VPWR_c_1179_n 0.00121566f $X=6.565 $Y=1.485 $X2=0 $Y2=0
cc_642 N_X_M1028_d N_VPWR_c_1179_n 0.00121566f $X=7.425 $Y=1.485 $X2=0 $Y2=0
cc_643 N_X_M1034_d N_VPWR_c_1179_n 0.00117537f $X=8.285 $Y=1.485 $X2=0 $Y2=0
cc_644 N_X_c_816_n N_VPWR_c_1179_n 0.00207897f $X=2.41 $Y=1.66 $X2=0 $Y2=0
cc_645 N_X_c_822_n N_VPWR_c_1179_n 0.00240527f $X=3.27 $Y=1.66 $X2=0 $Y2=0
cc_646 N_X_c_828_n N_VPWR_c_1179_n 0.00240527f $X=4.13 $Y=1.66 $X2=0 $Y2=0
cc_647 N_X_c_835_n N_VPWR_c_1179_n 0.00240527f $X=4.99 $Y=1.66 $X2=0 $Y2=0
cc_648 N_X_c_842_n N_VPWR_c_1179_n 0.00240527f $X=5.845 $Y=1.66 $X2=0 $Y2=0
cc_649 N_X_c_848_n N_VPWR_c_1179_n 0.00240527f $X=6.705 $Y=1.66 $X2=0 $Y2=0
cc_650 N_X_c_743_n N_VPWR_c_1179_n 0.00505204f $X=7.565 $Y=1.66 $X2=0 $Y2=0

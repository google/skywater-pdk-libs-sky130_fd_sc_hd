* File: sky130_fd_sc_hd__and3_1.spice
* Created: Thu Aug 27 14:07:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and3_1.pex.spice"
.subckt sky130_fd_sc_hd__and3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 A_109_47# N_A_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 A_181_47# N_B_M1002_g A_109_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g A_181_47# VNB NSHORT L=0.15 W=0.42 AD=0.103351
+ AS=0.0441 PD=0.894953 PS=0.63 NRD=61.428 NRS=14.28 M=1 R=2.8 SA=75000.9
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.159949 PD=1.82 PS=1.38505 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_A_27_47#_M1000_d N_B_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06615 AS=0.0567 PD=0.735 PS=0.69 NRD=18.7544 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_C_M1007_g N_A_27_47#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0841331 AS=0.06615 PD=0.789718 PS=0.735 NRD=68.1423 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.200317 PD=2.52 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__and3_1.pxi.spice"
*
.ends
*
*

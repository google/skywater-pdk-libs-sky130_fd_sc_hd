* File: sky130_fd_sc_hd__nor4b_1.spice
* Created: Tue Sep  1 19:19:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor4b_1.pex.spice"
.subckt sky130_fd_sc_hd__nor4b_1  VNB VPB C B A D_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* D_N	D_N
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_A_91_199#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=4.608 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=4.608 M=1 R=4.33333 SA=75001.1
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1007 N_A_91_199#_M1007_d N_D_N_M1007_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0787009 PD=1.36 PS=0.773271 NRD=0 NRS=17.856 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_161_297# N_A_91_199#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.52 PD=1.27 PS=3.04 NRD=15.7403 NRS=50.2153 M=1 R=6.66667
+ SA=75000.4 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1003 A_245_297# N_C_M1003_g A_161_297# VPB PHIGHVT L=0.15 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=15.7403 M=1 R=6.66667 SA=75000.9
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1008 A_341_297# N_B_M1008_g A_245_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.165 PD=1.27 PS=1.33 NRD=15.7403 NRS=21.6503 M=1 R=6.66667 SA=75001.3
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_341_297# VPB PHIGHVT L=0.15 W=1 AD=0.205282
+ AS=0.135 PD=1.88028 PS=1.27 NRD=0 NRS=15.7403 M=1 R=6.66667 SA=75001.8
+ SB=75000.4 A=0.15 P=2.3 MULT=1
MM1009 N_A_91_199#_M1009_d N_D_N_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1092 AS=0.0862183 PD=1.36 PS=0.789718 NRD=0 NRS=70.4866 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__nor4b_1.pxi.spice"
*
.ends
*
*

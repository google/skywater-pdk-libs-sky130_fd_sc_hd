* File: sky130_fd_sc_hd__a2bb2oi_4.spice
* Created: Thu Aug 27 14:03:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2bb2oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a2bb2oi_4  VNB VPB B1 B2 A1_N A2_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_B1_M1014_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75008.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_B1_M1023_g N_A_109_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75008.3 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1023_d N_B1_M1034_g N_A_109_47#_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75007.8 A=0.0975 P=1.6 MULT=1
MM1018 N_Y_M1018_d N_B2_M1018_g N_A_109_47#_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1018_d N_B2_M1019_g N_A_109_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75007 A=0.0975 P=1.6 MULT=1
MM1025 N_Y_M1025_d N_B2_M1025_g N_A_109_47#_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.3
+ SB=75006.6 A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1025_d N_B2_M1033_g N_A_109_47#_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.7
+ SB=75006.2 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1038_d N_B1_M1038_g N_A_109_47#_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75005.7 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1038_d N_A_751_21#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_751_21#_M1006_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1030 N_VGND_M1006_d N_A_751_21#_M1030_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1039 N_VGND_M1039_d N_A_751_21#_M1039_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.8
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1010 N_A_751_21#_M1010_d N_A1_N_M1010_g N_VGND_M1039_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75005.7 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1013 N_A_751_21#_M1010_d N_A1_N_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75006.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1016 N_A_751_21#_M1016_d N_A1_N_M1016_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75006.6 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1020 N_A_751_21#_M1016_d N_A1_N_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75007 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1017 N_A_751_21#_M1017_d N_A2_N_M1017_g N_VGND_M1020_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75007.4 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1026 N_A_751_21#_M1017_d N_A2_N_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75007.8 SB=75001 A=0.0975 P=1.6 MULT=1
MM1031 N_A_751_21#_M1031_d N_A2_N_M1031_g N_VGND_M1026_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75008.3 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1032 N_A_751_21#_M1031_d N_A2_N_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75008.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_A_27_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.8 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1004_d N_B1_M1007_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.4 A=0.15 P=2.3 MULT=1
MM1024 N_VPWR_M1024_d N_B1_M1024_g N_A_27_297#_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75004
+ A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1024_d N_B2_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1008 N_VPWR_M1008_d N_B2_M1008_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1027 N_VPWR_M1008_d N_B2_M1027_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1035 N_VPWR_M1035_d N_B2_M1035_g N_A_27_297#_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1036 N_VPWR_M1035_d N_B1_M1036_g N_A_27_297#_M1036_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1003 N_A_27_297#_M1036_s N_A_751_21#_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1011 N_A_27_297#_M1011_d N_A_751_21#_M1011_g N_Y_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1015 N_A_27_297#_M1011_d N_A_751_21#_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.4
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1021 N_A_27_297#_M1021_d N_A_751_21#_M1021_g N_Y_M1015_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_N_M1002_g N_A_1139_297#_M1002_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1002_d N_A1_N_M1005_g N_A_1139_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1009_d N_A1_N_M1009_g N_A_1139_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1009_d N_A1_N_M1028_g N_A_1139_297#_M1028_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1012 N_A_1139_297#_M1028_s N_A2_N_M1012_g N_A_751_21#_M1012_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75001.9 SB=75001.5 A=0.15 P=2.3 MULT=1
MM1022 N_A_1139_297#_M1022_d N_A2_N_M1022_g N_A_751_21#_M1012_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.3 SB=75001 A=0.15 P=2.3 MULT=1
MM1029 N_A_1139_297#_M1022_d N_A2_N_M1029_g N_A_751_21#_M1029_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75002.7 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1037 N_A_1139_297#_M1037_d N_A2_N_M1037_g N_A_751_21#_M1029_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75003.1 SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_153 VPB 0 6.77964e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__a2bb2oi_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__sdlclkp_1.spice
* Created: Tue Sep  1 19:31:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_hd__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_SCE_M1020_g N_A_27_47#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_27_47#_M1008_d N_GATE_M1008_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0722077 AS=0.0567 PD=0.807692 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1019 N_A_286_413#_M1019_d N_A_256_147#_M1019_g N_A_27_47#_M1008_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0675 AS=0.0618923 PD=0.735 PS=0.692308 NRD=14.988
+ NRS=18.324 M=1 R=2.4 SA=75001.1 SB=75001.9 A=0.054 P=1.02 MULT=1
MM1000 A_394_47# N_A_256_243#_M1000_g N_A_286_413#_M1019_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0833538 AS=0.0675 PD=0.812308 PS=0.735 NRD=58.836 NRS=16.656 M=1
+ R=2.4 SA=75001.6 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1018 N_VGND_M1018_d N_A_464_315#_M1018_g A_394_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.105491 AS=0.0972462 PD=0.855701 PS=0.947692 NRD=25.704 NRS=50.436 M=1
+ R=2.8 SA=75001.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_464_315#_M1003_d N_A_286_413#_M1003_g N_VGND_M1018_d VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.163259 PD=1.82 PS=1.3243 NRD=0 NRS=12.912 M=1
+ R=4.33333 SA=75001.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_A_256_147#_M1011_g N_A_256_243#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_256_147#_M1014_d N_CLK_M1014_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1094_47# N_A_464_315#_M1002_g N_A_1012_47#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0861 AS=0.1092 PD=0.83 PS=1.36 NRD=42.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_CLK_M1004_g A_1094_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.0861 PD=0.765421 PS=0.83 NRD=0 NRS=42.852 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_GCLK_M1013_d N_A_1012_47#_M1013_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 A_109_369# N_SCE_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_27_47#_M1005_d N_GATE_M1005_g A_109_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.134943 AS=0.0672 PD=1.22566 PS=0.85 NRD=13.8491 NRS=15.3857 M=1 R=4.26667
+ SA=75000.5 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1021 N_A_286_413#_M1021_d N_A_256_243#_M1021_g N_A_27_47#_M1005_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0693 AS=0.0885566 PD=0.75 PS=0.80434 NRD=11.7215 NRS=23.443
+ M=1 R=2.8 SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 A_382_413# N_A_256_147#_M1007_g N_A_286_413#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0693 PD=0.86 PS=0.75 NRD=77.3816 NRS=11.7215 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_464_315#_M1017_g A_382_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.108727 AS=0.0924 PD=0.90507 PS=0.86 NRD=70.3487 NRS=77.3816 M=1 R=2.8
+ SA=75002.1 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_A_464_315#_M1001_d N_A_286_413#_M1001_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.2533 AS=0.258873 PD=2.52 PS=2.15493 NRD=0 NRS=19.7 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_256_147#_M1015_g N_A_256_243#_M1015_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.16925 AS=0.1629 PD=1.37 PS=1.8 NRD=64.4584 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1006 N_A_256_147#_M1006_d N_CLK_M1006_g N_VPWR_M1015_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.16925 PD=1.8 PS=1.37 NRD=0 NRS=64.4584 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_A_1012_47#_M1016_d N_A_464_315#_M1016_g N_VPWR_M1016_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_1012_47#_M1016_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.116293 AS=0.0864 PD=1.03415 PS=0.91 NRD=7.683 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_GCLK_M1009_d N_A_1012_47#_M1009_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=3.9203 M=1 R=6.66667
+ SA=75000.8 SB=75000.2 A=0.15 P=2.3 MULT=1
DX22_noxref VNB VPB NWDIODE A=11.6844 P=17.77
*
.include "sky130_fd_sc_hd__sdlclkp_1.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_hd__a2bb2o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VGND A2_N a_313_47# VNB nshort w=420000u l=150000u
+  ad=8.0515e+11p pd=7.55e+06u as=1.134e+11p ps=1.38e+06u
M1001 a_82_21# a_313_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1002 X a_82_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.7e+11p pd=2.54e+06u as=8.098e+11p ps=7.22e+06u
M1003 VGND B1 a_646_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1004 a_646_47# B2 a_82_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_313_297# A1_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1006 a_313_47# A2_N a_313_297# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1007 VGND a_82_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1008 X a_82_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_574_369# a_313_47# a_82_21# VPB phighvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.664e+11p ps=1.8e+06u
M1010 a_574_369# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_313_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_82_21# X VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B2 a_574_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__a211o_1.spice.pex
* Created: Thu Aug 27 13:59:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A211O_1%A_80_21# 1 2 3 10 12 15 20 21 22 23 24 25 28
+ 30 34 38 40
c94 25 0 1.60767e-19 $X=0.825 $Y=1.595
r95 36 38 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.972 $Y=0.625
+ $X2=2.972 $Y2=0.53
r96 32 34 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.685
+ $X2=2.95 $Y2=1.85
r97 31 40 6.55019 $w=1.9e-07 $l=1.28e-07 $layer=LI1_cond $X=2.17 $Y=0.72
+ $X2=2.042 $Y2=0.72
r98 30 36 6.87974 $w=1.9e-07 $l=1.52263e-07 $layer=LI1_cond $X=2.86 $Y=0.72
+ $X2=2.972 $Y2=0.625
r99 30 31 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=2.86 $Y=0.72
+ $X2=2.17 $Y2=0.72
r100 26 40 0.307787 $w=2.55e-07 $l=9.5e-08 $layer=LI1_cond $X=2.042 $Y=0.625
+ $X2=2.042 $Y2=0.72
r101 26 28 4.29342 $w=2.53e-07 $l=9.5e-08 $layer=LI1_cond $X=2.042 $Y=0.625
+ $X2=2.042 $Y2=0.53
r102 24 32 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=2.805 $Y=1.595
+ $X2=2.95 $Y2=1.685
r103 24 25 122 $w=1.78e-07 $l=1.98e-06 $layer=LI1_cond $X=2.805 $Y=1.595
+ $X2=0.825 $Y2=1.595
r104 22 40 6.55019 $w=1.9e-07 $l=1.27e-07 $layer=LI1_cond $X=1.915 $Y=0.72
+ $X2=2.042 $Y2=0.72
r105 22 23 63.6268 $w=1.88e-07 $l=1.09e-06 $layer=LI1_cond $X=1.915 $Y=0.72
+ $X2=0.825 $Y2=0.72
r106 21 41 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.685 $Y=1.16
+ $X2=0.475 $Y2=1.16
r107 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.685
+ $Y=1.16 $X2=0.685 $Y2=1.16
r108 18 25 6.92652 $w=1.8e-07 $l=1.51456e-07 $layer=LI1_cond $X=0.712 $Y=1.505
+ $X2=0.825 $Y2=1.595
r109 18 20 17.6708 $w=2.23e-07 $l=3.45e-07 $layer=LI1_cond $X=0.712 $Y=1.505
+ $X2=0.712 $Y2=1.16
r110 17 23 6.87974 $w=1.9e-07 $l=1.5331e-07 $layer=LI1_cond $X=0.712 $Y=0.815
+ $X2=0.825 $Y2=0.72
r111 17 20 17.6708 $w=2.23e-07 $l=3.45e-07 $layer=LI1_cond $X=0.712 $Y=0.815
+ $X2=0.712 $Y2=1.16
r112 13 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.16
r113 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.325
+ $X2=0.475 $Y2=1.985
r114 10 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.16
r115 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r116 3 34 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=1.485 $X2=2.96 $Y2=1.85
r117 2 38 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.96 $Y2=0.53
r118 1 28 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.07 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%A2 1 3 6 8 14
r33 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.215 $Y=1.16
+ $X2=1.425 $Y2=1.16
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r35 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.325
+ $X2=1.425 $Y2=1.16
r36 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.425 $Y=1.325
+ $X2=1.425 $Y2=1.985
r37 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%A1 3 6 8 11 12 13
r35 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.16
+ $X2=1.845 $Y2=1.325
r36 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.16
+ $X2=1.845 $Y2=0.995
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.845
+ $Y=1.16 $X2=1.845 $Y2=1.16
r38 8 12 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.62 $Y=1.16
+ $X2=1.845 $Y2=1.16
r39 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.855 $Y=1.985
+ $X2=1.855 $Y2=1.325
r40 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.855 $Y=0.56
+ $X2=1.855 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%B1 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.16
+ $X2=2.325 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.16
+ $X2=2.325 $Y2=0.995
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.325
+ $Y=1.16 $X2=2.325 $Y2=1.16
r36 8 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.54 $Y=1.16
+ $X2=2.325 $Y2=1.16
r37 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=1.985
+ $X2=2.285 $Y2=1.325
r38 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.285 $Y=0.56
+ $X2=2.285 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%C1 1 3 6 8 13
r26 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.745 $Y=1.16
+ $X2=2.955 $Y2=1.16
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.16
r29 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.985
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=0.995
+ $X2=2.745 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.745 $Y=0.995
+ $X2=2.745 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%X 1 2 7 8 9 10 11 12 22 38
r15 20 38 0.412815 $w=3.33e-07 $l=1.2e-08 $layer=LI1_cond $X=0.257 $Y=1.518
+ $X2=0.257 $Y2=1.53
r16 11 12 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=2.21
r17 11 41 8.04536 $w=2.63e-07 $l=1.85e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=1.685
r18 10 41 4.62931 $w=3.33e-07 $l=1.19e-07 $layer=LI1_cond $X=0.257 $Y=1.566
+ $X2=0.257 $Y2=1.685
r19 10 38 1.23845 $w=3.33e-07 $l=3.6e-08 $layer=LI1_cond $X=0.257 $Y=1.566
+ $X2=0.257 $Y2=1.53
r20 10 20 1.27285 $w=3.33e-07 $l=3.7e-08 $layer=LI1_cond $X=0.257 $Y=1.481
+ $X2=0.257 $Y2=1.518
r21 9 10 10.0108 $w=3.33e-07 $l=2.91e-07 $layer=LI1_cond $X=0.257 $Y=1.19
+ $X2=0.257 $Y2=1.481
r22 8 9 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=0.85
+ $X2=0.257 $Y2=1.19
r23 7 8 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.85
r24 7 22 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.4
r25 2 10 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r26 1 22 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%VPWR 1 2 9 13 15 17 22 32 33 36 39 44
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 37 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.64 $Y2=2.72
r58 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.64 $Y2=2.72
r65 22 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 19 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r68 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 15 44 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=2.635
+ $X2=1.64 $Y2=2.72
r71 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.64 $Y=2.635
+ $X2=1.64 $Y2=2.36
r72 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.72
r73 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2
r74 2 13 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.485 $X2=1.64 $Y2=2.36
r75 1 9 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%A_217_297# 1 2 7 9 11 13 15
r28 13 20 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=2.105 $Y=2.095
+ $X2=2.105 $Y2=1.98
r29 13 15 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=2.105 $Y=2.095
+ $X2=2.105 $Y2=2.29
r30 12 18 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.305 $Y=1.98
+ $X2=1.175 $Y2=1.98
r31 11 20 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.975 $Y=1.98
+ $X2=2.105 $Y2=1.98
r32 11 12 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=1.98
+ $X2=1.305 $Y2=1.98
r33 7 18 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=1.175 $Y=2.095
+ $X2=1.175 $Y2=1.98
r34 7 9 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.175 $Y=2.095
+ $X2=1.175 $Y2=2.29
r35 2 20 600 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.485 $X2=2.07 $Y2=1.95
r36 2 15 600 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.485 $X2=2.07 $Y2=2.29
r37 1 18 600 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=1.95
r38 1 9 600 $w=1.7e-07 $l=8.65246e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__A211O_1%VGND 1 2 9 11 18 25 26 31 37 39 44
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r49 35 37 10.5432 $w=5.38e-07 $l=2e-07 $layer=LI1_cond $X=1.15 $Y=0.185 $X2=1.35
+ $Y2=0.185
r50 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r51 33 35 0.442992 $w=5.38e-07 $l=2e-08 $layer=LI1_cond $X=1.13 $Y=0.185
+ $X2=1.15 $Y2=0.185
r52 30 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r53 30 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r54 29 33 9.74582 $w=5.38e-07 $l=4.4e-07 $layer=LI1_cond $X=0.69 $Y=0.185
+ $X2=1.13 $Y2=0.185
r55 29 31 7.99599 $w=5.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.185
+ $X2=0.605 $Y2=0.185
r56 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r58 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r59 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.515
+ $Y2=0
r60 23 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.99
+ $Y2=0
r61 22 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r62 22 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r63 21 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.35
+ $Y2=0
r64 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r65 18 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.515
+ $Y2=0
r66 18 21 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.07
+ $Y2=0
r67 15 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.605
+ $Y2=0
r68 15 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 11 44 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r70 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r71 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.36
r72 2 9 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.235 $X2=2.515 $Y2=0.36
r73 1 33 91 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.13 $Y2=0.36
.ends


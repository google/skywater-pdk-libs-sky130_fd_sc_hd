* File: sky130_fd_sc_hd__buf_12.pex.spice
* Created: Tue Sep  1 18:58:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_12%A 3 7 11 15 19 23 25 27 31 33 34 35 36
c82 36 0 1.28215e-19 $X=1.575 $Y=1.19
r83 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.405
+ $Y=1.16 $X2=1.405 $Y2=1.16
r84 42 44 14.9526 $w=2.74e-07 $l=8.5e-08 $layer=POLY_cond $X=0.385 $Y=1.16
+ $X2=0.47 $Y2=1.16
r85 36 49 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.575 $Y=1.175
+ $X2=1.405 $Y2=1.175
r86 35 49 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=1.115 $Y=1.175
+ $X2=1.405 $Y2=1.175
r87 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.655 $Y=1.175
+ $X2=1.115 $Y2=1.175
r88 33 34 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.315 $Y=1.175
+ $X2=0.655 $Y2=1.175
r89 33 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.16 $X2=0.385 $Y2=1.16
r90 25 48 57.1715 $w=2.74e-07 $l=3.25e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.405 $Y2=1.16
r91 25 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r92 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r93 17 48 16.7117 $w=2.74e-07 $l=9.5e-08 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.405 $Y2=1.16
r94 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r95 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r96 9 17 73.8832 $w=2.74e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r97 9 44 73.8832 $w=2.74e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r98 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r99 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r100 5 44 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r101 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.985
r102 1 44 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r103 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_12%A_109_47# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 117 119 120 121 122 125 131
+ 133 136 138 144 148 150 151 166
c270 166 0 1.28215e-19 $X=6.77 $Y=1.16
c271 144 0 1.80041e-19 $X=4.3 $Y=1.16
r272 165 166 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.35 $Y=1.16
+ $X2=6.77 $Y2=1.16
r273 164 165 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.93 $Y=1.16
+ $X2=6.35 $Y2=1.16
r274 163 164 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.51 $Y=1.16
+ $X2=5.93 $Y2=1.16
r275 162 163 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.09 $Y=1.16
+ $X2=5.51 $Y2=1.16
r276 161 162 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.67 $Y=1.16
+ $X2=5.09 $Y2=1.16
r277 158 159 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.83 $Y=1.16
+ $X2=4.25 $Y2=1.16
r278 157 158 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.41 $Y=1.16
+ $X2=3.83 $Y2=1.16
r279 156 157 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.99 $Y=1.16
+ $X2=3.41 $Y2=1.16
r280 155 156 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.57 $Y=1.16
+ $X2=2.99 $Y2=1.16
r281 145 161 82.2043 $w=2.7e-07 $l=3.7e-07 $layer=POLY_cond $X=4.3 $Y=1.16
+ $X2=4.67 $Y2=1.16
r282 145 159 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=4.3 $Y=1.16
+ $X2=4.25 $Y2=1.16
r283 144 145 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=4.3
+ $Y=1.16 $X2=4.3 $Y2=1.16
r284 142 155 68.8738 $w=2.7e-07 $l=3.1e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.57 $Y2=1.16
r285 142 152 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.15 $Y2=1.16
r286 141 144 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=2.26 $Y=1.16
+ $X2=4.3 $Y2=1.16
r287 141 142 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r288 139 151 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.015 $Y=1.16
+ $X2=1.927 $Y2=1.16
r289 139 141 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.015 $Y=1.16
+ $X2=2.26 $Y2=1.16
r290 138 148 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.927 $Y=1.445
+ $X2=1.927 $Y2=1.53
r291 137 151 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.927 $Y=1.245
+ $X2=1.927 $Y2=1.16
r292 137 138 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.927 $Y=1.245
+ $X2=1.927 $Y2=1.445
r293 136 151 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.927 $Y=1.075
+ $X2=1.927 $Y2=1.16
r294 135 136 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.927 $Y=0.905
+ $X2=1.927 $Y2=1.075
r295 134 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.82
+ $X2=1.52 $Y2=0.82
r296 133 135 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.84 $Y=0.82
+ $X2=1.927 $Y2=0.905
r297 133 134 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.84 $Y=0.82
+ $X2=1.605 $Y2=0.82
r298 129 150 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.735
+ $X2=1.52 $Y2=0.82
r299 129 131 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.52 $Y=0.735
+ $X2=1.52 $Y2=0.56
r300 125 127 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.52 $Y=1.63
+ $X2=1.52 $Y2=2.31
r301 123 148 26.5529 $w=1.68e-07 $l=4.07e-07 $layer=LI1_cond $X=1.52 $Y=1.53
+ $X2=1.927 $Y2=1.53
r302 123 125 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.52 $Y=1.615
+ $X2=1.52 $Y2=1.63
r303 121 123 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=1.53
+ $X2=1.52 $Y2=1.53
r304 121 122 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.355 $Y=1.53
+ $X2=0.845 $Y2=1.53
r305 119 150 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=0.82
+ $X2=1.52 $Y2=0.82
r306 119 120 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.82
+ $X2=0.765 $Y2=0.82
r307 115 120 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.765 $Y2=0.82
r308 115 117 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.68 $Y=0.735
+ $X2=0.68 $Y2=0.56
r309 111 113 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=2.31
r310 109 122 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.68 $Y=1.615
+ $X2=0.845 $Y2=1.53
r311 109 111 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.68 $Y=1.615
+ $X2=0.68 $Y2=1.63
r312 105 166 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.16
r313 105 107 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.77 $Y=1.295
+ $X2=6.77 $Y2=1.985
r314 101 166 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=1.16
r315 101 103 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.77 $Y=1.025
+ $X2=6.77 $Y2=0.56
r316 97 165 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.16
r317 97 99 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.35 $Y=1.295
+ $X2=6.35 $Y2=1.985
r318 93 165 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=1.16
r319 93 95 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.35 $Y=1.025
+ $X2=6.35 $Y2=0.56
r320 89 164 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.16
r321 89 91 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.985
r322 85 164 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=1.16
r323 85 87 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.93 $Y=1.025
+ $X2=5.93 $Y2=0.56
r324 81 163 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.16
r325 81 83 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.51 $Y=1.295
+ $X2=5.51 $Y2=1.985
r326 77 163 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=1.16
r327 77 79 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.51 $Y=1.025
+ $X2=5.51 $Y2=0.56
r328 73 162 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.16
r329 73 75 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.09 $Y=1.295
+ $X2=5.09 $Y2=1.985
r330 69 162 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=1.16
r331 69 71 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.09 $Y=1.025
+ $X2=5.09 $Y2=0.56
r332 65 161 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.16
r333 65 67 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.67 $Y=1.295
+ $X2=4.67 $Y2=1.985
r334 61 161 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=1.16
r335 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.67 $Y=1.025
+ $X2=4.67 $Y2=0.56
r336 57 159 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.16
r337 57 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.25 $Y=1.295
+ $X2=4.25 $Y2=1.985
r338 53 159 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=1.16
r339 53 55 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
r340 49 158 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.16
r341 49 51 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.295
+ $X2=3.83 $Y2=1.985
r342 45 158 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.16
r343 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r344 41 157 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.16
r345 41 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.41 $Y=1.295
+ $X2=3.41 $Y2=1.985
r346 37 157 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=1.16
r347 37 39 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.41 $Y=1.025
+ $X2=3.41 $Y2=0.56
r348 33 156 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.16
r349 33 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.99 $Y=1.295
+ $X2=2.99 $Y2=1.985
r350 29 156 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=1.16
r351 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.99 $Y=1.025
+ $X2=2.99 $Y2=0.56
r352 25 155 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.16
r353 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.57 $Y=1.295
+ $X2=2.57 $Y2=1.985
r354 21 155 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=1.16
r355 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.57 $Y=1.025
+ $X2=2.57 $Y2=0.56
r356 17 152 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.16
r357 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.15 $Y=1.295
+ $X2=2.15 $Y2=1.985
r358 13 152 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=1.16
r359 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.15 $Y=1.025
+ $X2=2.15 $Y2=0.56
r360 4 127 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.31
r361 4 125 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.63
r362 3 113 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.31
r363 3 111 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r364 2 131 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.56
r365 1 117 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_12%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 48
+ 52 56 60 62 64 69 70 72 73 75 76 77 78 79 81 97 102 107 116 119 122 126
c130 38 0 1.80041e-19 $X=1.94 $Y=2
r131 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r132 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r136 111 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r137 111 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r138 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r139 108 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=2.72
+ $X2=6.14 $Y2=2.72
r140 108 110 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.305 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 107 125 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=6.815 $Y=2.72
+ $X2=7.087 $Y2=2.72
r142 107 110 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.815 $Y=2.72
+ $X2=6.67 $Y2=2.72
r143 106 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r144 106 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r145 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 103 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.3 $Y2=2.72
r147 103 105 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.465 $Y=2.72
+ $X2=5.75 $Y2=2.72
r148 102 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=2.72
+ $X2=6.14 $Y2=2.72
r149 102 105 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.975 $Y=2.72
+ $X2=5.75 $Y2=2.72
r150 101 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r151 101 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r152 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r153 98 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.46 $Y2=2.72
r154 98 100 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.83 $Y2=2.72
r155 97 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.3 $Y2=2.72
r156 97 100 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=4.83 $Y2=2.72
r157 96 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r158 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r159 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r161 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r162 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r163 83 113 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r164 81 90 0.271737 $w=4.8e-07 $l=9.55e-07 $layer=MET1_cond $X=0.655 $Y=2.72
+ $X2=1.61 $Y2=2.72
r165 81 114 0.12093 $w=4.8e-07 $l=4.25e-07 $layer=MET1_cond $X=0.655 $Y=2.72
+ $X2=0.23 $Y2=2.72
r166 79 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r167 79 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.655 $Y=2.72
+ $X2=0.345 $Y2=2.72
r168 77 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.45 $Y2=2.72
r169 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.62 $Y2=2.72
r170 75 92 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.53 $Y2=2.72
r171 75 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.72
+ $X2=2.78 $Y2=2.72
r172 74 95 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.45 $Y2=2.72
r173 74 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.78 $Y2=2.72
r174 72 89 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r175 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.94 $Y2=2.72
r176 71 92 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=2.72
+ $X2=1.94 $Y2=2.72
r178 69 79 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.655 $Y2=2.72
r179 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r180 68 89 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r181 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r182 64 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.98 $Y=1.66
+ $X2=6.98 $Y2=2.34
r183 62 125 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.98 $Y=2.635
+ $X2=7.087 $Y2=2.72
r184 62 67 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.98 $Y=2.635
+ $X2=6.98 $Y2=2.34
r185 58 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2.72
r186 58 60 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.14 $Y=2.635
+ $X2=6.14 $Y2=2
r187 54 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2.72
r188 54 56 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.3 $Y=2.635
+ $X2=5.3 $Y2=2
r189 50 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2.72
r190 50 52 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.46 $Y=2.635
+ $X2=4.46 $Y2=2
r191 49 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=2.72
+ $X2=3.62 $Y2=2.72
r192 48 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.46 $Y2=2.72
r193 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=3.785 $Y2=2.72
r194 44 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r195 44 46 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2
r196 40 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2.72
r197 40 42 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.78 $Y=2.635
+ $X2=2.78 $Y2=2
r198 36 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2.72
r199 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=2.635
+ $X2=1.94 $Y2=2
r200 32 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r201 32 34 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r202 28 113 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r203 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r204 9 67 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.98 $Y2=2.34
r205 9 64 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.98 $Y2=1.66
r206 8 60 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.005
+ $Y=1.485 $X2=6.14 $Y2=2
r207 7 56 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.485 $X2=5.3 $Y2=2
r208 6 52 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.325
+ $Y=1.485 $X2=4.46 $Y2=2
r209 5 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.485 $X2=3.62 $Y2=2
r210 4 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2
r211 3 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r212 2 34 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r213 1 30 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_12%X 1 2 3 4 5 6 7 8 9 10 11 12 39 43 45 46 47
+ 48 51 55 57 59 63 67 71 75 79 83 87 89 90 92 94 95 109 118
r143 117 118 11.6455 $w=8.78e-07 $l=8.4e-07 $layer=LI1_cond $X=5.72 $Y=1.175
+ $X2=6.56 $Y2=1.175
r144 116 117 11.6455 $w=8.78e-07 $l=8.4e-07 $layer=LI1_cond $X=4.88 $Y=1.175
+ $X2=5.72 $Y2=1.175
r145 95 116 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=4.88 $Y=1.615
+ $X2=4.88 $Y2=1.175
r146 95 116 1.17841 $w=8.78e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=1.175
+ $X2=4.88 $Y2=1.175
r147 95 109 7.61063 $w=2.53e-07 $l=1.4e-07 $layer=LI1_cond $X=4.88 $Y=1.615
+ $X2=4.88 $Y2=1.755
r148 93 95 21.2684 $w=3.38e-07 $l=5.85e-07 $layer=LI1_cond $X=4.125 $Y=1.53
+ $X2=4.71 $Y2=1.53
r149 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=1.53
+ $X2=4.04 $Y2=1.53
r150 91 95 23.0544 $w=3.08e-07 $l=5.85e-07 $layer=LI1_cond $X=4.125 $Y=0.82
+ $X2=4.71 $Y2=0.82
r151 91 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=0.82
+ $X2=4.04 $Y2=0.82
r152 85 118 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=6.56 $Y=1.615
+ $X2=6.56 $Y2=1.175
r153 85 87 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.56 $Y=1.615
+ $X2=6.56 $Y2=1.755
r154 81 118 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=6.56 $Y=0.735
+ $X2=6.56 $Y2=1.175
r155 81 83 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.56 $Y=0.735
+ $X2=6.56 $Y2=0.56
r156 77 117 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=5.72 $Y=1.615
+ $X2=5.72 $Y2=1.175
r157 77 79 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.72 $Y=1.615
+ $X2=5.72 $Y2=1.755
r158 73 117 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=5.72 $Y=0.735
+ $X2=5.72 $Y2=1.175
r159 73 75 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.72 $Y=0.735
+ $X2=5.72 $Y2=0.56
r160 69 116 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=4.88 $Y=0.735
+ $X2=4.88 $Y2=1.175
r161 69 71 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.88 $Y=0.735
+ $X2=4.88 $Y2=0.56
r162 65 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=1.615
+ $X2=4.04 $Y2=1.53
r163 65 67 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.04 $Y=1.615
+ $X2=4.04 $Y2=1.755
r164 61 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.735
+ $X2=4.04 $Y2=0.82
r165 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.04 $Y=0.735
+ $X2=4.04 $Y2=0.56
r166 60 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=1.53
+ $X2=3.2 $Y2=1.53
r167 59 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=1.53
+ $X2=4.04 $Y2=1.53
r168 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.955 $Y=1.53
+ $X2=3.285 $Y2=1.53
r169 58 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=0.82
+ $X2=3.2 $Y2=0.82
r170 57 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0.82
+ $X2=4.04 $Y2=0.82
r171 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.955 $Y=0.82
+ $X2=3.285 $Y2=0.82
r172 53 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.615 $X2=3.2
+ $Y2=1.53
r173 53 55 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.2 $Y=1.615
+ $X2=3.2 $Y2=1.755
r174 49 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.735 $X2=3.2
+ $Y2=0.82
r175 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.2 $Y=0.735
+ $X2=3.2 $Y2=0.56
r176 47 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.53
+ $X2=3.2 $Y2=1.53
r177 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=1.53
+ $X2=2.445 $Y2=1.53
r178 45 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.82
+ $X2=3.2 $Y2=0.82
r179 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.115 $Y=0.82
+ $X2=2.445 $Y2=0.82
r180 41 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=1.615
+ $X2=2.445 $Y2=1.53
r181 41 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.36 $Y=1.615
+ $X2=2.36 $Y2=1.755
r182 37 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.445 $Y2=0.82
r183 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.36 $Y2=0.56
r184 12 87 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=6.425
+ $Y=1.485 $X2=6.56 $Y2=1.755
r185 11 79 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=5.585
+ $Y=1.485 $X2=5.72 $Y2=1.755
r186 10 109 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=4.745
+ $Y=1.485 $X2=4.88 $Y2=1.755
r187 9 67 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.485 $X2=4.04 $Y2=1.755
r188 8 55 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.2 $Y2=1.755
r189 7 43 300 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.755
r190 6 83 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=6.425
+ $Y=0.235 $X2=6.56 $Y2=0.56
r191 5 75 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.56
r192 4 71 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.88 $Y2=0.56
r193 3 63 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.56
r194 2 51 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.2 $Y2=0.56
r195 1 39 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_12%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 48
+ 52 56 60 62 64 67 68 70 71 72 73 74 76 78 81 95 100 105 114 117 120 123 127
+ 131
r153 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r154 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r155 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r156 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r158 112 131 0.119507 $w=4.8e-07 $l=4.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.65 $Y2=0
r159 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r160 109 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r161 109 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r162 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r163 106 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0
+ $X2=6.14 $Y2=0
r164 106 108 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.305 $Y=0
+ $X2=6.67 $Y2=0
r165 105 126 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=7.087 $Y2=0
r166 105 108 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.67 $Y2=0
r167 104 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r168 104 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r169 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r170 101 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.3 $Y2=0
r171 101 103 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.75 $Y2=0
r172 100 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=6.14 $Y2=0
r173 100 103 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.975 $Y=0
+ $X2=5.75 $Y2=0
r174 99 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r175 99 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=4.37 $Y2=0
r176 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r177 96 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=4.46 $Y2=0
r178 96 98 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=4.83 $Y2=0
r179 95 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.3
+ $Y2=0
r180 95 98 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=0
+ $X2=4.83 $Y2=0
r181 94 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r182 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r183 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r184 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r185 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r186 88 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r187 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r188 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r189 85 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r190 79 111 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r191 79 81 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.65 $Y2=0
r192 78 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r193 76 115 0.140848 $w=4.8e-07 $l=4.95e-07 $layer=MET1_cond $X=0.655 $Y=0
+ $X2=1.15 $Y2=0
r194 76 131 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.655 $Y=0
+ $X2=0.65 $Y2=0
r195 74 78 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.655 $Y=0
+ $X2=0.935 $Y2=0
r196 74 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r197 74 81 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.655 $Y=0 $X2=0.65
+ $Y2=0
r198 72 93 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.45
+ $Y2=0
r199 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=0 $X2=3.62
+ $Y2=0
r200 70 90 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.53
+ $Y2=0
r201 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.78
+ $Y2=0
r202 69 93 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=3.45 $Y2=0
r203 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.78
+ $Y2=0
r204 67 87 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r205 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.94
+ $Y2=0
r206 66 90 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.105 $Y=0
+ $X2=2.53 $Y2=0
r207 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.94
+ $Y2=0
r208 62 126 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.98 $Y=0.085
+ $X2=7.087 $Y2=0
r209 62 64 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.98 $Y=0.085
+ $X2=6.98 $Y2=0.38
r210 58 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0
r211 58 60 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.14 $Y=0.085
+ $X2=6.14 $Y2=0.4
r212 54 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0
r213 54 56 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0.4
r214 50 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0
r215 50 52 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.46 $Y=0.085
+ $X2=4.46 $Y2=0.4
r216 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.785 $Y=0 $X2=3.62
+ $Y2=0
r217 48 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.46 $Y2=0
r218 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=3.785 $Y2=0
r219 44 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0
r220 44 46 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.62 $Y=0.085
+ $X2=3.62 $Y2=0.4
r221 40 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0
r222 40 42 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.78 $Y=0.085
+ $X2=2.78 $Y2=0.4
r223 36 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r224 36 38 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.4
r225 32 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r226 32 34 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.4
r227 28 111 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r228 28 30 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r229 9 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.845
+ $Y=0.235 $X2=6.98 $Y2=0.38
r230 8 60 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.005
+ $Y=0.235 $X2=6.14 $Y2=0.4
r231 7 56 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.3 $Y2=0.4
r232 6 52 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=4.325
+ $Y=0.235 $X2=4.46 $Y2=0.4
r233 5 46 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.4
r234 4 42 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.4
r235 3 38 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.4
r236 2 34 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.4
r237 1 30 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


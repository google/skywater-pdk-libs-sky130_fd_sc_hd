* File: sky130_fd_sc_hd__clkdlybuf4s18_2.spice
* Created: Tue Sep  1 19:00:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__clkdlybuf4s18_2.pex.spice"
.subckt sky130_fd_sc_hd__clkdlybuf4s18_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0921252 AS=0.1134 PD=0.824299 PS=1.38 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_227_47#_M1003_d N_A_27_47#_M1003_g N_VGND_M1000_d VNB NSHORT L=0.18
+ W=0.65 AD=0.17225 AS=0.142575 PD=1.83 PS=1.2757 NRD=0 NRS=11.988 M=1 R=3.61111
+ SA=90000.5 SB=90000.2 A=0.117 P=1.66 MULT=1
MM1005 N_VGND_M1005_d N_A_227_47#_M1005_g N_A_334_47#_M1005_s VNB NSHORT L=0.18
+ W=0.65 AD=0.175682 AS=0.17225 PD=1.36682 PS=1.83 NRD=15.684 NRS=0 M=1
+ R=3.61111 SA=90000.2 SB=90001 A=0.117 P=1.66 MULT=1
MM1001 N_VGND_M1005_d N_A_334_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.113518 AS=0.0588 PD=0.883178 PS=0.7 NRD=31.428 NRS=0 M=1 R=2.8 SA=75000.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_334_47#_M1008_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1575 AS=0.0588 PD=1.59 PS=0.7 NRD=27.132 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.204945 AS=0.27 PD=1.53846 PS=2.54 NRD=13.7703 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1009 N_A_227_47#_M1009_d N_A_27_47#_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2173 AS=0.168055 PD=2.17 PS=1.26154 NRD=0 NRS=11.9973 M=1
+ R=4.55556 SA=90000.7 SB=90000.2 A=0.1476 P=2 MULT=1
MM1007 N_VPWR_M1007_d N_A_227_47#_M1007_g N_A_334_47#_M1007_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.195764 AS=0.2173 PD=1.32912 PS=2.17 NRD=22.8126 NRS=0 M=1
+ R=4.55556 SA=90000.2 SB=90001.3 A=0.1476 P=2 MULT=1
MM1002 N_VPWR_M1007_d N_A_334_47#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.238736 AS=0.14 PD=1.62088 PS=1.28 NRD=19.7 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_334_47#_M1006_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.375 AS=0.14 PD=2.75 PS=1.28 NRD=18.715 NRS=0 M=1 R=6.66667 SA=75001.2
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__clkdlybuf4s18_2.pxi.spice"
*
.ends
*
*

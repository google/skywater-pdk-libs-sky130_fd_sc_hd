* File: sky130_fd_sc_hd__nor4bb_4.pxi.spice
* Created: Thu Aug 27 14:33:38 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4BB_4%C_N N_C_N_c_151_n N_C_N_M1018_g N_C_N_M1005_g C_N
+ N_C_N_c_153_n C_N PM_SKY130_FD_SC_HD__NOR4BB_4%C_N
x_PM_SKY130_FD_SC_HD__NOR4BB_4%D_N N_D_N_c_176_n N_D_N_M1011_g N_D_N_M1035_g D_N
+ N_D_N_c_178_n D_N PM_SKY130_FD_SC_HD__NOR4BB_4%D_N
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A_197_47# N_A_197_47#_M1011_d N_A_197_47#_M1035_d
+ N_A_197_47#_c_215_n N_A_197_47#_M1012_g N_A_197_47#_M1003_g
+ N_A_197_47#_c_216_n N_A_197_47#_M1019_g N_A_197_47#_M1008_g
+ N_A_197_47#_c_217_n N_A_197_47#_M1025_g N_A_197_47#_M1023_g
+ N_A_197_47#_c_218_n N_A_197_47#_M1033_g N_A_197_47#_M1029_g
+ N_A_197_47#_c_219_n N_A_197_47#_c_231_n N_A_197_47#_c_220_n
+ N_A_197_47#_c_221_n N_A_197_47#_c_222_n N_A_197_47#_c_223_n
+ N_A_197_47#_c_224_n N_A_197_47#_c_225_n N_A_197_47#_c_226_n
+ PM_SKY130_FD_SC_HD__NOR4BB_4%A_197_47#
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A_27_297# N_A_27_297#_M1018_s N_A_27_297#_M1005_s
+ N_A_27_297#_c_339_n N_A_27_297#_M1020_g N_A_27_297#_M1000_g
+ N_A_27_297#_c_340_n N_A_27_297#_M1026_g N_A_27_297#_M1009_g
+ N_A_27_297#_c_341_n N_A_27_297#_M1027_g N_A_27_297#_M1014_g
+ N_A_27_297#_c_342_n N_A_27_297#_M1034_g N_A_27_297#_M1030_g
+ N_A_27_297#_c_343_n N_A_27_297#_c_353_n N_A_27_297#_c_344_n
+ N_A_27_297#_c_355_n N_A_27_297#_c_356_n N_A_27_297#_c_345_n
+ N_A_27_297#_c_346_n N_A_27_297#_c_347_n N_A_27_297#_c_357_n
+ N_A_27_297#_c_348_n PM_SKY130_FD_SC_HD__NOR4BB_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_4%B N_B_c_483_n N_B_M1002_g N_B_M1010_g N_B_c_484_n
+ N_B_M1006_g N_B_M1015_g N_B_c_485_n N_B_M1013_g N_B_M1031_g N_B_c_486_n
+ N_B_M1021_g N_B_M1032_g B N_B_c_487_n N_B_c_488_n
+ PM_SKY130_FD_SC_HD__NOR4BB_4%B
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A N_A_c_561_n N_A_M1007_g N_A_M1001_g N_A_c_562_n
+ N_A_M1017_g N_A_M1004_g N_A_c_563_n N_A_M1022_g N_A_M1016_g N_A_c_564_n
+ N_A_M1028_g N_A_M1024_g A N_A_c_565_n N_A_c_566_n
+ PM_SKY130_FD_SC_HD__NOR4BB_4%A
x_PM_SKY130_FD_SC_HD__NOR4BB_4%VPWR N_VPWR_M1005_d N_VPWR_M1001_s N_VPWR_M1016_s
+ N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n VPWR N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_632_n N_VPWR_c_641_n
+ N_VPWR_c_642_n N_VPWR_c_643_n PM_SKY130_FD_SC_HD__NOR4BB_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A_311_297# N_A_311_297#_M1003_d
+ N_A_311_297#_M1008_d N_A_311_297#_M1029_d N_A_311_297#_M1009_d
+ N_A_311_297#_M1030_d N_A_311_297#_c_738_n N_A_311_297#_c_753_n
+ N_A_311_297#_c_778_p N_A_311_297#_c_739_n N_A_311_297#_c_740_n
+ N_A_311_297#_c_757_n N_A_311_297#_c_769_n
+ PM_SKY130_FD_SC_HD__NOR4BB_4%A_311_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_4%Y N_Y_M1012_d N_Y_M1025_d N_Y_M1020_s N_Y_M1027_s
+ N_Y_M1002_s N_Y_M1013_s N_Y_M1007_d N_Y_M1022_d N_Y_M1003_s N_Y_M1023_s
+ N_Y_c_804_n N_Y_c_787_n N_Y_c_788_n N_Y_c_818_n N_Y_c_789_n N_Y_c_790_n
+ N_Y_c_828_n N_Y_c_791_n N_Y_c_859_n N_Y_c_792_n N_Y_c_875_n N_Y_c_793_n
+ N_Y_c_882_n N_Y_c_794_n N_Y_c_887_n N_Y_c_795_n N_Y_c_907_n N_Y_c_796_n
+ N_Y_c_797_n N_Y_c_798_n N_Y_c_799_n N_Y_c_800_n N_Y_c_801_n Y N_Y_c_803_n Y
+ PM_SKY130_FD_SC_HD__NOR4BB_4%Y
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A_729_297# N_A_729_297#_M1000_s
+ N_A_729_297#_M1014_s N_A_729_297#_M1010_d N_A_729_297#_M1031_d
+ N_A_729_297#_c_984_n N_A_729_297#_c_985_n N_A_729_297#_c_986_n
+ N_A_729_297#_c_987_n N_A_729_297#_c_988_n N_A_729_297#_c_989_n
+ N_A_729_297#_c_990_n PM_SKY130_FD_SC_HD__NOR4BB_4%A_729_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_4%A_1087_297# N_A_1087_297#_M1010_s
+ N_A_1087_297#_M1015_s N_A_1087_297#_M1032_s N_A_1087_297#_M1004_d
+ N_A_1087_297#_M1024_d N_A_1087_297#_c_1042_n N_A_1087_297#_c_1050_n
+ N_A_1087_297#_c_1043_n N_A_1087_297#_c_1100_n N_A_1087_297#_c_1052_n
+ N_A_1087_297#_c_1044_n N_A_1087_297#_c_1077_n N_A_1087_297#_c_1045_n
+ N_A_1087_297#_c_1081_n N_A_1087_297#_c_1046_n N_A_1087_297#_c_1047_n
+ N_A_1087_297#_c_1048_n N_A_1087_297#_c_1087_n N_A_1087_297#_c_1049_n
+ PM_SKY130_FD_SC_HD__NOR4BB_4%A_1087_297#
x_PM_SKY130_FD_SC_HD__NOR4BB_4%VGND N_VGND_M1018_d N_VGND_M1012_s N_VGND_M1019_s
+ N_VGND_M1033_s N_VGND_M1026_d N_VGND_M1034_d N_VGND_M1006_d N_VGND_M1021_d
+ N_VGND_M1017_s N_VGND_M1028_s N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n
+ N_VGND_c_1108_n N_VGND_c_1109_n N_VGND_c_1110_n N_VGND_c_1111_n
+ N_VGND_c_1112_n N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n
+ N_VGND_c_1116_n N_VGND_c_1117_n N_VGND_c_1118_n N_VGND_c_1119_n
+ N_VGND_c_1120_n N_VGND_c_1121_n N_VGND_c_1122_n N_VGND_c_1123_n
+ N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n VGND N_VGND_c_1127_n
+ N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n VGND PM_SKY130_FD_SC_HD__NOR4BB_4%VGND
cc_1 VNB N_C_N_c_151_n 0.0218983f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB C_N 0.00888732f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_153_n 0.0368018f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_4 VNB N_D_N_c_176_n 0.0200575f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_5 VNB D_N 0.00175619f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_D_N_c_178_n 0.0346454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_197_47#_c_215_n 0.0191932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_197_47#_c_216_n 0.0157805f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_9 VNB N_A_197_47#_c_217_n 0.0157832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_197_47#_c_218_n 0.0156271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_197_47#_c_219_n 0.00590512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_197_47#_c_220_n 0.0082966f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_197_47#_c_221_n 0.00205232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_197_47#_c_222_n 0.00455221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_197_47#_c_223_n 0.00129226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_197_47#_c_224_n 0.00655567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_197_47#_c_225_n 0.00210943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_197_47#_c_226_n 0.0660655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_339_n 0.0159825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_340_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_21 VNB N_A_27_297#_c_341_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_297#_c_342_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_297#_c_343_n 0.0191875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_297#_c_344_n 0.00785471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_297#_c_345_n 0.00257705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_297#_c_346_n 0.0022324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_297#_c_347_n 0.0109791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_297#_c_348_n 0.0687477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_B_c_483_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_30 VNB N_B_c_484_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_31 VNB N_B_c_485_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_B_c_486_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_B_c_487_n 0.0159176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_B_c_488_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_c_561_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_36 VNB N_A_c_562_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_37 VNB N_A_c_563_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_c_564_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_c_565_n 0.0184554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_c_566_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_632_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_787_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_788_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_789_n 8.79379e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_790_n 0.00578238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_791_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_792_n 0.00904229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_Y_c_793_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Y_c_794_n 0.00429924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_795_n 0.00440603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Y_c_796_n 0.00207163f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_797_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Y_c_798_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_Y_c_799_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_Y_c_800_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_Y_c_801_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1105_n 0.0046277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1106_n 0.0213623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1107_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1108_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1109_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1110_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1111_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1112_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1113_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1114_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1115_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1116_n 0.0329389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1117_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1118_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1119_n 0.0166678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1120_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1121_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1122_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1123_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1124_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1125_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1126_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1127_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1128_n 0.0208123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1129_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1130_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1131_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1132_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1133_n 0.431404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VPB N_C_N_M1005_g 0.0252901f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_87 VPB C_N 0.00503237f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_88 VPB N_C_N_c_153_n 0.00954313f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_89 VPB N_D_N_M1035_g 0.0229305f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_90 VPB D_N 2.38458e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_91 VPB N_D_N_c_178_n 0.00916147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_197_47#_M1003_g 0.0217479f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_93 VPB N_A_197_47#_M1008_g 0.0178669f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.22
cc_94 VPB N_A_197_47#_M1023_g 0.0178525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_197_47#_M1029_g 0.0180891f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_197_47#_c_231_n 0.00716661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_197_47#_c_223_n 0.00554061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_197_47#_c_226_n 0.0101926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_27_297#_M1000_g 0.0178834f $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_100 VPB N_A_27_297#_M1009_g 0.0182122f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.22
cc_101 VPB N_A_27_297#_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_27_297#_M1030_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_27_297#_c_353_n 0.0165958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_297#_c_344_n 0.00341622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_27_297#_c_355_n 0.00813339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_27_297#_c_356_n 0.00105715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_297#_c_357_n 0.0224114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_297#_c_348_n 0.0107446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_B_M1010_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_110 VPB N_B_M1015_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_B_M1031_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_B_M1032_g 0.018818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_B_c_488_n 0.0108798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_M1001_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_115 VPB N_A_M1004_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_M1016_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_M1024_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_c_566_n 0.0108808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_633_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.28 $Y2=1.16
cc_120 VPB N_VPWR_c_634_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.22
cc_121 VPB N_VPWR_c_635_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_636_n 0.0147956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_637_n 0.153718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_638_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_639_n 0.0174963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_632_n 0.0568121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_641_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_642_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_643_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_311_297#_c_738_n 0.00412953f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.22
cc_131 VPB N_A_311_297#_c_739_n 0.00166092f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_311_297#_c_740_n 0.00451061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_Y_c_789_n 8.79379e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_Y_c_803_n 0.00645226f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_729_297#_c_984_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_729_297#_c_985_n 0.0179302f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.22
cc_137 VPB N_A_729_297#_c_986_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_729_297#_c_987_n 0.00184676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_729_297#_c_988_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_729_297#_c_989_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_729_297#_c_990_n 0.00225182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_1087_297#_c_1042_n 0.00516601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_1087_297#_c_1043_n 0.00198437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_1087_297#_c_1044_n 0.00414042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_1087_297#_c_1045_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_1087_297#_c_1046_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_1087_297#_c_1047_n 0.0102662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1087_297#_c_1048_n 0.0327764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_1087_297#_c_1049_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 N_C_N_c_151_n N_D_N_c_176_n 0.0255799f $X=0.49 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_151 N_C_N_M1005_g N_D_N_M1035_g 0.0255799f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_152 N_C_N_c_153_n N_D_N_c_178_n 0.0255799f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_153 N_C_N_c_151_n N_A_197_47#_c_219_n 5.34423e-19 $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_C_N_c_151_n N_A_27_297#_c_343_n 0.0064154f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C_N_c_151_n N_A_27_297#_c_344_n 0.00974094f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_156 C_N N_A_27_297#_c_344_n 0.0217359f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_C_N_c_151_n N_A_27_297#_c_347_n 0.0109681f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_158 C_N N_A_27_297#_c_347_n 0.0239086f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_159 N_C_N_c_153_n N_A_27_297#_c_347_n 0.00661237f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_160 N_C_N_M1005_g N_A_27_297#_c_357_n 0.019012f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_161 C_N N_A_27_297#_c_357_n 0.0253738f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_162 N_C_N_c_153_n N_A_27_297#_c_357_n 0.0017135f $X=0.49 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C_N_M1005_g N_VPWR_c_633_n 0.00875461f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_164 N_C_N_M1005_g N_VPWR_c_636_n 0.00343969f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_165 N_C_N_M1005_g N_VPWR_c_632_n 0.00499499f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_166 N_C_N_c_151_n N_VGND_c_1105_n 0.00268723f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_167 N_C_N_c_151_n N_VGND_c_1128_n 0.0042235f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_168 N_C_N_c_151_n N_VGND_c_1133_n 0.00673103f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_169 N_D_N_c_176_n N_A_197_47#_c_219_n 0.00641302f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_D_N_M1035_g N_A_197_47#_c_231_n 0.00259637f $X=0.91 $Y=1.985 $X2=0
+ $Y2=0
cc_171 D_N N_A_197_47#_c_231_n 0.0190949f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_172 N_D_N_c_178_n N_A_197_47#_c_231_n 0.00641049f $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_173 D_N N_A_197_47#_c_220_n 7.38065e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_174 N_D_N_c_176_n N_A_197_47#_c_221_n 0.00263836f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_175 D_N N_A_197_47#_c_221_n 0.0270711f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_176 N_D_N_c_178_n N_A_197_47#_c_221_n 0.00767804f $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_177 N_D_N_c_176_n N_A_197_47#_c_222_n 0.00220008f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_D_N_c_178_n N_A_197_47#_c_222_n 0.0019362f $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_179 N_D_N_M1035_g N_A_197_47#_c_223_n 0.00455646f $X=0.91 $Y=1.985 $X2=0
+ $Y2=0
cc_180 D_N N_A_197_47#_c_223_n 0.00626859f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_181 N_D_N_c_178_n N_A_197_47#_c_223_n 2.91626e-19 $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_182 D_N N_A_197_47#_c_225_n 0.0150481f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_183 N_D_N_c_178_n N_A_197_47#_c_225_n 7.70091e-19 $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_184 D_N N_A_197_47#_c_226_n 4.3473e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_185 N_D_N_c_178_n N_A_197_47#_c_226_n 0.00574752f $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_186 N_D_N_c_176_n N_A_27_297#_c_343_n 5.2253e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_187 N_D_N_c_176_n N_A_27_297#_c_344_n 0.0102774f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_188 D_N N_A_27_297#_c_344_n 0.0187708f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_189 N_D_N_M1035_g N_A_27_297#_c_355_n 0.017313f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_190 N_D_N_c_176_n N_A_27_297#_c_347_n 7.24136e-19 $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_D_N_M1035_g N_VPWR_c_633_n 0.0115803f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_192 N_D_N_M1035_g N_VPWR_c_637_n 0.00343969f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_193 N_D_N_M1035_g N_VPWR_c_632_n 0.0054428f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_194 N_D_N_M1035_g N_A_311_297#_c_738_n 0.00417809f $X=0.91 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_D_N_c_176_n N_VGND_c_1105_n 0.00268723f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_196 N_D_N_c_176_n N_VGND_c_1106_n 0.00541359f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_197 N_D_N_c_176_n N_VGND_c_1107_n 0.0018189f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_198 N_D_N_c_176_n N_VGND_c_1133_n 0.0108548f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_197_47#_c_218_n N_A_27_297#_c_339_n 0.0276379f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_197_47#_M1029_g N_A_27_297#_M1000_g 0.0276379f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_197_47#_c_219_n N_A_27_297#_c_343_n 0.00523552f $X=1.12 $Y=0.39 $X2=0
+ $Y2=0
cc_202 N_A_197_47#_c_221_n N_A_27_297#_c_344_n 7.99055e-19 $X=1.285 $Y=0.82
+ $X2=0 $Y2=0
cc_203 N_A_197_47#_M1035_d N_A_27_297#_c_355_n 0.0071406f $X=0.985 $Y=1.485
+ $X2=0 $Y2=0
cc_204 N_A_197_47#_M1003_g N_A_27_297#_c_355_n 0.0128101f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_197_47#_M1008_g N_A_27_297#_c_355_n 0.0103496f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_197_47#_M1023_g N_A_27_297#_c_355_n 0.0103496f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_197_47#_M1029_g N_A_27_297#_c_355_n 0.0115089f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_197_47#_c_231_n N_A_27_297#_c_355_n 0.0472379f $X=1.465 $Y=1.62 $X2=0
+ $Y2=0
cc_209 N_A_197_47#_c_224_n N_A_27_297#_c_355_n 0.00494954f $X=2.68 $Y=1.16 $X2=0
+ $Y2=0
cc_210 N_A_197_47#_c_226_n N_A_27_297#_c_356_n 0.00617381f $X=3.15 $Y=1.16 $X2=0
+ $Y2=0
cc_211 N_A_197_47#_c_226_n N_A_27_297#_c_345_n 0.00174654f $X=3.15 $Y=1.16 $X2=0
+ $Y2=0
cc_212 N_A_197_47#_c_221_n N_A_27_297#_c_347_n 0.00710591f $X=1.285 $Y=0.82
+ $X2=0 $Y2=0
cc_213 N_A_197_47#_c_226_n N_A_27_297#_c_348_n 0.0276379f $X=3.15 $Y=1.16 $X2=0
+ $Y2=0
cc_214 N_A_197_47#_M1003_g N_VPWR_c_637_n 0.00357877f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_197_47#_M1008_g N_VPWR_c_637_n 0.00357877f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_197_47#_M1023_g N_VPWR_c_637_n 0.00357877f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_197_47#_M1029_g N_VPWR_c_637_n 0.00357877f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_197_47#_M1035_d N_VPWR_c_632_n 0.00344981f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_219 N_A_197_47#_M1003_g N_VPWR_c_632_n 0.00655123f $X=1.89 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_197_47#_M1008_g N_VPWR_c_632_n 0.00522516f $X=2.31 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_197_47#_M1023_g N_VPWR_c_632_n 0.00522516f $X=2.73 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_197_47#_M1029_g N_VPWR_c_632_n 0.00525237f $X=3.15 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_197_47#_c_231_n N_A_311_297#_M1003_d 0.00320594f $X=1.465 $Y=1.62
+ $X2=-0.19 $Y2=-0.24
cc_224 N_A_197_47#_c_223_n N_A_311_297#_M1003_d 6.5575e-19 $X=1.55 $Y=1.535
+ $X2=-0.19 $Y2=-0.24
cc_225 N_A_197_47#_M1003_g N_A_311_297#_c_738_n 0.00970685f $X=1.89 $Y=1.985
+ $X2=0 $Y2=0
cc_226 N_A_197_47#_M1008_g N_A_311_297#_c_738_n 0.00970685f $X=2.31 $Y=1.985
+ $X2=0 $Y2=0
cc_227 N_A_197_47#_M1023_g N_A_311_297#_c_738_n 0.00970685f $X=2.73 $Y=1.985
+ $X2=0 $Y2=0
cc_228 N_A_197_47#_M1029_g N_A_311_297#_c_738_n 0.00969293f $X=3.15 $Y=1.985
+ $X2=0 $Y2=0
cc_229 N_A_197_47#_c_215_n N_Y_c_804_n 0.00730874f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_197_47#_c_216_n N_Y_c_804_n 0.00630972f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_197_47#_c_217_n N_Y_c_804_n 5.22228e-19 $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_197_47#_c_219_n N_Y_c_804_n 0.00484536f $X=1.12 $Y=0.39 $X2=0 $Y2=0
cc_233 N_A_197_47#_c_216_n N_Y_c_787_n 0.00870364f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_197_47#_c_217_n N_Y_c_787_n 0.00870364f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_197_47#_c_224_n N_Y_c_787_n 0.0356734f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_197_47#_c_226_n N_Y_c_787_n 0.00222133f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_197_47#_c_215_n N_Y_c_788_n 0.00331113f $X=1.89 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_197_47#_c_216_n N_Y_c_788_n 0.00113286f $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A_197_47#_c_219_n N_Y_c_788_n 2.84208e-19 $X=1.12 $Y=0.39 $X2=0 $Y2=0
cc_240 N_A_197_47#_c_220_n N_Y_c_788_n 0.00961296f $X=1.465 $Y=0.82 $X2=0 $Y2=0
cc_241 N_A_197_47#_c_224_n N_Y_c_788_n 0.026256f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_197_47#_c_226_n N_Y_c_788_n 0.00230339f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_197_47#_c_216_n N_Y_c_818_n 5.22228e-19 $X=2.31 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_197_47#_c_217_n N_Y_c_818_n 0.00630972f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_197_47#_c_218_n N_Y_c_818_n 0.00630972f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_197_47#_c_217_n N_Y_c_789_n 0.0017444f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_197_47#_M1023_g N_Y_c_789_n 0.0017444f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_197_47#_c_218_n N_Y_c_789_n 0.00248022f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_197_47#_M1029_g N_Y_c_789_n 0.00874379f $X=3.15 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_197_47#_c_224_n N_Y_c_789_n 0.0127974f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_197_47#_c_226_n N_Y_c_789_n 0.0171266f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_197_47#_c_218_n N_Y_c_790_n 0.0053917f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_197_47#_c_218_n N_Y_c_828_n 5.22228e-19 $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_197_47#_c_217_n N_Y_c_796_n 0.00113286f $X=2.73 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_197_47#_c_218_n N_Y_c_796_n 0.00409494f $X=3.15 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_197_47#_c_224_n N_Y_c_796_n 0.00549243f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_197_47#_c_226_n N_Y_c_796_n 0.00280876f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_197_47#_M1003_g N_Y_c_803_n 0.00949903f $X=1.89 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A_197_47#_M1008_g N_Y_c_803_n 0.0123561f $X=2.31 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_197_47#_M1023_g N_Y_c_803_n 0.0123561f $X=2.73 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A_197_47#_c_231_n N_Y_c_803_n 0.0127689f $X=1.465 $Y=1.62 $X2=0 $Y2=0
cc_262 N_A_197_47#_c_223_n N_Y_c_803_n 0.00815099f $X=1.55 $Y=1.535 $X2=0 $Y2=0
cc_263 N_A_197_47#_c_224_n N_Y_c_803_n 0.0733702f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_197_47#_c_226_n N_Y_c_803_n 0.00716348f $X=3.15 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_197_47#_c_220_n N_VGND_M1012_s 0.00356387f $X=1.465 $Y=0.82 $X2=0
+ $Y2=0
cc_266 N_A_197_47#_c_219_n N_VGND_c_1106_n 0.0209752f $X=1.12 $Y=0.39 $X2=0
+ $Y2=0
cc_267 N_A_197_47#_c_220_n N_VGND_c_1106_n 0.00480319f $X=1.465 $Y=0.82 $X2=0
+ $Y2=0
cc_268 N_A_197_47#_c_215_n N_VGND_c_1107_n 0.00316354f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_197_47#_c_219_n N_VGND_c_1107_n 0.0152424f $X=1.12 $Y=0.39 $X2=0
+ $Y2=0
cc_270 N_A_197_47#_c_220_n N_VGND_c_1107_n 0.00321628f $X=1.465 $Y=0.82 $X2=0
+ $Y2=0
cc_271 N_A_197_47#_c_224_n N_VGND_c_1107_n 0.00460552f $X=2.68 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_197_47#_c_216_n N_VGND_c_1108_n 0.00146448f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_A_197_47#_c_217_n N_VGND_c_1108_n 0.00146448f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_197_47#_c_218_n N_VGND_c_1109_n 0.00146448f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_197_47#_c_215_n N_VGND_c_1117_n 0.00541359f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_197_47#_c_216_n N_VGND_c_1117_n 0.00423334f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_197_47#_c_217_n N_VGND_c_1119_n 0.00423334f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_197_47#_c_218_n N_VGND_c_1119_n 0.00423261f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_197_47#_M1011_d N_VGND_c_1133_n 0.00209319f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_280 N_A_197_47#_c_215_n N_VGND_c_1133_n 0.0108276f $X=1.89 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_197_47#_c_216_n N_VGND_c_1133_n 0.0057163f $X=2.31 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_197_47#_c_217_n N_VGND_c_1133_n 0.0057163f $X=2.73 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_197_47#_c_218_n N_VGND_c_1133_n 0.00574217f $X=3.15 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_197_47#_c_219_n N_VGND_c_1133_n 0.0124119f $X=1.12 $Y=0.39 $X2=0
+ $Y2=0
cc_285 N_A_197_47#_c_220_n N_VGND_c_1133_n 0.00855541f $X=1.465 $Y=0.82 $X2=0
+ $Y2=0
cc_286 N_A_27_297#_c_346_n N_B_c_487_n 0.0140827f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_27_297#_c_348_n N_B_c_487_n 0.00155889f $X=4.83 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_344_n N_VPWR_M1005_d 5.44303e-19 $X=0.7 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_289 N_A_27_297#_c_357_n N_VPWR_M1005_d 0.00238861f $X=0.785 $Y=1.79 $X2=-0.19
+ $Y2=-0.24
cc_290 N_A_27_297#_c_357_n N_VPWR_c_633_n 0.0172472f $X=0.785 $Y=1.79 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_c_353_n N_VPWR_c_636_n 0.0187476f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_292 N_A_27_297#_c_357_n N_VPWR_c_636_n 0.00237903f $X=0.785 $Y=1.79 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_M1000_g N_VPWR_c_637_n 0.00357877f $X=3.57 $Y=1.985 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_M1009_g N_VPWR_c_637_n 0.00357877f $X=3.99 $Y=1.985 $X2=0
+ $Y2=0
cc_295 N_A_27_297#_M1014_g N_VPWR_c_637_n 0.00357877f $X=4.41 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_27_297#_M1030_g N_VPWR_c_637_n 0.00357877f $X=4.83 $Y=1.985 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_c_355_n N_VPWR_c_637_n 0.0100714f $X=3.355 $Y=1.96 $X2=0
+ $Y2=0
cc_298 N_A_27_297#_M1005_s N_VPWR_c_632_n 0.00246869f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_299 N_A_27_297#_M1000_g N_VPWR_c_632_n 0.00525237f $X=3.57 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A_27_297#_M1009_g N_VPWR_c_632_n 0.00522516f $X=3.99 $Y=1.985 $X2=0
+ $Y2=0
cc_301 N_A_27_297#_M1014_g N_VPWR_c_632_n 0.00522516f $X=4.41 $Y=1.985 $X2=0
+ $Y2=0
cc_302 N_A_27_297#_M1030_g N_VPWR_c_632_n 0.00655123f $X=4.83 $Y=1.985 $X2=0
+ $Y2=0
cc_303 N_A_27_297#_c_353_n N_VPWR_c_632_n 0.0105763f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_355_n N_VPWR_c_632_n 0.0204215f $X=3.355 $Y=1.96 $X2=0
+ $Y2=0
cc_305 N_A_27_297#_c_357_n N_VPWR_c_632_n 0.00576627f $X=0.785 $Y=1.79 $X2=0
+ $Y2=0
cc_306 N_A_27_297#_c_355_n N_A_311_297#_M1003_d 0.00619198f $X=3.355 $Y=1.96
+ $X2=-0.19 $Y2=-0.24
cc_307 N_A_27_297#_c_355_n N_A_311_297#_M1008_d 0.00317879f $X=3.355 $Y=1.96
+ $X2=0 $Y2=0
cc_308 N_A_27_297#_c_355_n N_A_311_297#_M1029_d 0.00437149f $X=3.355 $Y=1.96
+ $X2=0 $Y2=0
cc_309 N_A_27_297#_c_356_n N_A_311_297#_M1029_d 0.00371963f $X=3.44 $Y=1.875
+ $X2=0 $Y2=0
cc_310 N_A_27_297#_c_355_n N_A_311_297#_c_738_n 0.10478f $X=3.355 $Y=1.96 $X2=0
+ $Y2=0
cc_311 N_A_27_297#_M1000_g N_A_311_297#_c_753_n 0.0101149f $X=3.57 $Y=1.985
+ $X2=0 $Y2=0
cc_312 N_A_27_297#_M1009_g N_A_311_297#_c_753_n 0.00988743f $X=3.99 $Y=1.985
+ $X2=0 $Y2=0
cc_313 N_A_27_297#_M1014_g N_A_311_297#_c_739_n 0.00984328f $X=4.41 $Y=1.985
+ $X2=0 $Y2=0
cc_314 N_A_27_297#_M1030_g N_A_311_297#_c_739_n 0.00988743f $X=4.83 $Y=1.985
+ $X2=0 $Y2=0
cc_315 N_A_27_297#_M1000_g N_A_311_297#_c_757_n 0.00252196f $X=3.57 $Y=1.985
+ $X2=0 $Y2=0
cc_316 N_A_27_297#_M1009_g N_A_311_297#_c_757_n 2.35016e-19 $X=3.99 $Y=1.985
+ $X2=0 $Y2=0
cc_317 N_A_27_297#_c_355_n N_Y_M1003_s 0.00317879f $X=3.355 $Y=1.96 $X2=0 $Y2=0
cc_318 N_A_27_297#_c_355_n N_Y_M1023_s 0.00314682f $X=3.355 $Y=1.96 $X2=0 $Y2=0
cc_319 N_A_27_297#_c_339_n N_Y_c_818_n 5.22228e-19 $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_27_297#_c_339_n N_Y_c_789_n 0.00107087f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_27_297#_M1000_g N_Y_c_789_n 2.73143e-19 $X=3.57 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_27_297#_c_355_n N_Y_c_789_n 0.00853911f $X=3.355 $Y=1.96 $X2=0 $Y2=0
cc_323 N_A_27_297#_c_356_n N_Y_c_789_n 0.0320778f $X=3.44 $Y=1.875 $X2=0 $Y2=0
cc_324 N_A_27_297#_c_345_n N_Y_c_789_n 0.0169426f $X=3.525 $Y=1.18 $X2=0 $Y2=0
cc_325 N_A_27_297#_c_348_n N_Y_c_789_n 3.20211e-19 $X=4.83 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_27_297#_c_339_n N_Y_c_790_n 0.00865562f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_27_297#_c_345_n N_Y_c_790_n 0.014165f $X=3.525 $Y=1.18 $X2=0 $Y2=0
cc_328 N_A_27_297#_c_346_n N_Y_c_790_n 0.00615875f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_27_297#_c_339_n N_Y_c_828_n 0.00630972f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_27_297#_c_340_n N_Y_c_828_n 0.00630972f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_27_297#_c_341_n N_Y_c_828_n 5.22228e-19 $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_27_297#_c_340_n N_Y_c_791_n 0.00870364f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_27_297#_c_341_n N_Y_c_791_n 0.00870364f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_27_297#_c_346_n N_Y_c_791_n 0.0362443f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_27_297#_c_348_n N_Y_c_791_n 0.00222133f $X=4.83 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_27_297#_c_340_n N_Y_c_859_n 5.22228e-19 $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A_27_297#_c_341_n N_Y_c_859_n 0.00630972f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_27_297#_c_342_n N_Y_c_859_n 0.0109565f $X=4.83 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_27_297#_c_342_n N_Y_c_792_n 0.0109318f $X=4.83 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_27_297#_c_346_n N_Y_c_792_n 0.00826974f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_27_297#_c_339_n N_Y_c_797_n 0.00113286f $X=3.57 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A_27_297#_c_340_n N_Y_c_797_n 0.00113286f $X=3.99 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A_27_297#_c_346_n N_Y_c_797_n 0.0266272f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_27_297#_c_348_n N_Y_c_797_n 0.00230339f $X=4.83 $Y=1.16 $X2=0 $Y2=0
cc_345 N_A_27_297#_c_341_n N_Y_c_798_n 0.00113286f $X=4.41 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A_27_297#_c_342_n N_Y_c_798_n 0.00113286f $X=4.83 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A_27_297#_c_346_n N_Y_c_798_n 0.0266272f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A_27_297#_c_348_n N_Y_c_798_n 0.00230339f $X=4.83 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A_27_297#_c_355_n N_Y_c_803_n 0.065068f $X=3.355 $Y=1.96 $X2=0 $Y2=0
cc_350 N_A_27_297#_M1009_g N_A_729_297#_c_984_n 0.0109047f $X=3.99 $Y=1.985
+ $X2=0 $Y2=0
cc_351 N_A_27_297#_M1014_g N_A_729_297#_c_984_n 0.01094f $X=4.41 $Y=1.985 $X2=0
+ $Y2=0
cc_352 N_A_27_297#_c_346_n N_A_729_297#_c_984_n 0.0416643f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_353 N_A_27_297#_c_348_n N_A_729_297#_c_984_n 0.00211509f $X=4.83 $Y=1.16
+ $X2=0 $Y2=0
cc_354 N_A_27_297#_M1030_g N_A_729_297#_c_985_n 0.0130871f $X=4.83 $Y=1.985
+ $X2=0 $Y2=0
cc_355 N_A_27_297#_c_346_n N_A_729_297#_c_985_n 0.0110239f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_356 N_A_27_297#_M1000_g N_A_729_297#_c_987_n 2.36936e-19 $X=3.57 $Y=1.985
+ $X2=0 $Y2=0
cc_357 N_A_27_297#_c_356_n N_A_729_297#_c_987_n 0.00714067f $X=3.44 $Y=1.875
+ $X2=0 $Y2=0
cc_358 N_A_27_297#_c_346_n N_A_729_297#_c_987_n 0.0171602f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_359 N_A_27_297#_c_348_n N_A_729_297#_c_987_n 0.00219557f $X=4.83 $Y=1.16
+ $X2=0 $Y2=0
cc_360 N_A_27_297#_c_346_n N_A_729_297#_c_988_n 0.0204292f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_361 N_A_27_297#_c_348_n N_A_729_297#_c_988_n 0.00219557f $X=4.83 $Y=1.16
+ $X2=0 $Y2=0
cc_362 N_A_27_297#_c_347_n N_VGND_M1018_d 0.00188206f $X=0.7 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_363 N_A_27_297#_c_347_n N_VGND_c_1105_n 0.0122105f $X=0.7 $Y=0.81 $X2=0 $Y2=0
cc_364 N_A_27_297#_c_339_n N_VGND_c_1109_n 0.00146448f $X=3.57 $Y=0.995 $X2=0
+ $Y2=0
cc_365 N_A_27_297#_c_340_n N_VGND_c_1110_n 0.00146448f $X=3.99 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_27_297#_c_341_n N_VGND_c_1110_n 0.00146339f $X=4.41 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_339_n N_VGND_c_1121_n 0.00423334f $X=3.57 $Y=0.995 $X2=0
+ $Y2=0
cc_368 N_A_27_297#_c_340_n N_VGND_c_1121_n 0.00423334f $X=3.99 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_343_n N_VGND_c_1128_n 0.0226078f $X=0.28 $Y=0.39 $X2=0
+ $Y2=0
cc_370 N_A_27_297#_c_347_n N_VGND_c_1128_n 0.00201529f $X=0.7 $Y=0.81 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_341_n N_VGND_c_1130_n 0.00423334f $X=4.41 $Y=0.995 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_342_n N_VGND_c_1130_n 0.00423334f $X=4.83 $Y=0.995 $X2=0
+ $Y2=0
cc_373 N_A_27_297#_c_342_n N_VGND_c_1131_n 0.00335921f $X=4.83 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_M1018_s N_VGND_c_1133_n 0.00221616f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_c_339_n N_VGND_c_1133_n 0.0057435f $X=3.57 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_c_340_n N_VGND_c_1133_n 0.0057163f $X=3.99 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_c_341_n N_VGND_c_1133_n 0.0057163f $X=4.41 $Y=0.995 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_342_n N_VGND_c_1133_n 0.0070399f $X=4.83 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_27_297#_c_343_n N_VGND_c_1133_n 0.0134533f $X=0.28 $Y=0.39 $X2=0
+ $Y2=0
cc_380 N_A_27_297#_c_347_n N_VGND_c_1133_n 0.00454306f $X=0.7 $Y=0.81 $X2=0
+ $Y2=0
cc_381 N_B_c_486_n N_A_c_561_n 0.0195974f $X=7.03 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_382 N_B_M1032_g N_A_M1001_g 0.0195974f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_383 N_B_c_487_n N_A_c_565_n 0.0121231f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_384 N_B_c_488_n N_A_c_565_n 2.62535e-19 $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_385 N_B_c_487_n N_A_c_566_n 2.62535e-19 $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_386 N_B_c_488_n N_A_c_566_n 0.0195974f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B_M1010_g N_VPWR_c_637_n 0.00357877f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_388 N_B_M1015_g N_VPWR_c_637_n 0.00357877f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_389 N_B_M1031_g N_VPWR_c_637_n 0.00357877f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_390 N_B_M1032_g N_VPWR_c_637_n 0.00357877f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_391 N_B_M1010_g N_VPWR_c_632_n 0.00655123f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_392 N_B_M1015_g N_VPWR_c_632_n 0.00522516f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_393 N_B_M1031_g N_VPWR_c_632_n 0.00522516f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_394 N_B_M1032_g N_VPWR_c_632_n 0.00525237f $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_395 N_B_c_483_n N_Y_c_792_n 0.0109318f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_396 N_B_c_487_n N_Y_c_792_n 0.0501575f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_397 N_B_c_483_n N_Y_c_875_n 0.0109565f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_398 N_B_c_484_n N_Y_c_875_n 0.00630972f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B_c_485_n N_Y_c_875_n 5.22228e-19 $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_400 N_B_c_484_n N_Y_c_793_n 0.00870364f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_401 N_B_c_485_n N_Y_c_793_n 0.00870364f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_402 N_B_c_487_n N_Y_c_793_n 0.0362443f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_403 N_B_c_488_n N_Y_c_793_n 0.00222133f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_404 N_B_c_484_n N_Y_c_882_n 5.22228e-19 $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_405 N_B_c_485_n N_Y_c_882_n 0.00630972f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_406 N_B_c_486_n N_Y_c_882_n 0.00630972f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B_c_486_n N_Y_c_794_n 0.00865686f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_408 N_B_c_487_n N_Y_c_794_n 0.00826974f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_409 N_B_c_486_n N_Y_c_887_n 5.22228e-19 $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_410 N_B_c_483_n N_Y_c_799_n 0.00113286f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_411 N_B_c_484_n N_Y_c_799_n 0.00113286f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_412 N_B_c_487_n N_Y_c_799_n 0.0266272f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_413 N_B_c_488_n N_Y_c_799_n 0.00230339f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_414 N_B_c_485_n N_Y_c_800_n 0.00113286f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_415 N_B_c_486_n N_Y_c_800_n 0.00113286f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_416 N_B_c_487_n N_Y_c_800_n 0.0266272f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_417 N_B_c_488_n N_Y_c_800_n 0.00230339f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_418 N_B_M1010_g N_A_729_297#_c_985_n 0.0130871f $X=5.77 $Y=1.985 $X2=0 $Y2=0
cc_419 N_B_c_487_n N_A_729_297#_c_985_n 0.0527326f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_420 N_B_M1015_g N_A_729_297#_c_986_n 0.01094f $X=6.19 $Y=1.985 $X2=0 $Y2=0
cc_421 N_B_M1031_g N_A_729_297#_c_986_n 0.0109258f $X=6.61 $Y=1.985 $X2=0 $Y2=0
cc_422 N_B_c_487_n N_A_729_297#_c_986_n 0.0416643f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_423 N_B_c_488_n N_A_729_297#_c_986_n 0.00211509f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_424 N_B_c_487_n N_A_729_297#_c_989_n 0.0204292f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_425 N_B_c_488_n N_A_729_297#_c_989_n 0.00219557f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_426 N_B_M1032_g N_A_729_297#_c_990_n 2.57315e-19 $X=7.03 $Y=1.985 $X2=0 $Y2=0
cc_427 N_B_c_487_n N_A_729_297#_c_990_n 0.0204292f $X=6.94 $Y=1.16 $X2=0 $Y2=0
cc_428 N_B_c_488_n N_A_729_297#_c_990_n 0.00219557f $X=7.03 $Y=1.16 $X2=0 $Y2=0
cc_429 N_B_M1010_g N_A_1087_297#_c_1050_n 0.00988743f $X=5.77 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_B_M1015_g N_A_1087_297#_c_1050_n 0.00988743f $X=6.19 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_B_M1031_g N_A_1087_297#_c_1052_n 0.00984328f $X=6.61 $Y=1.985 $X2=0
+ $Y2=0
cc_432 N_B_M1032_g N_A_1087_297#_c_1052_n 0.0121747f $X=7.03 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_B_M1032_g N_A_1087_297#_c_1044_n 2.57315e-19 $X=7.03 $Y=1.985 $X2=0
+ $Y2=0
cc_434 N_B_c_484_n N_VGND_c_1111_n 0.00146339f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_485_n N_VGND_c_1111_n 0.00146448f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_436 N_B_c_486_n N_VGND_c_1112_n 0.00146448f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_483_n N_VGND_c_1123_n 0.00423334f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_438 N_B_c_484_n N_VGND_c_1123_n 0.00423334f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_485_n N_VGND_c_1125_n 0.00423334f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B_c_486_n N_VGND_c_1125_n 0.00423334f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_483_n N_VGND_c_1131_n 0.00335921f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_483_n N_VGND_c_1133_n 0.0070399f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_484_n N_VGND_c_1133_n 0.0057163f $X=6.19 $Y=0.995 $X2=0 $Y2=0
cc_444 N_B_c_485_n N_VGND_c_1133_n 0.0057163f $X=6.61 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_486_n N_VGND_c_1133_n 0.0057435f $X=7.03 $Y=0.995 $X2=0 $Y2=0
cc_446 N_A_M1001_g N_VPWR_c_634_n 0.00302074f $X=7.45 $Y=1.985 $X2=0 $Y2=0
cc_447 N_A_M1004_g N_VPWR_c_634_n 0.00157837f $X=7.87 $Y=1.985 $X2=0 $Y2=0
cc_448 N_A_M1016_g N_VPWR_c_635_n 0.00157837f $X=8.29 $Y=1.985 $X2=0 $Y2=0
cc_449 N_A_M1024_g N_VPWR_c_635_n 0.00302074f $X=8.71 $Y=1.985 $X2=0 $Y2=0
cc_450 N_A_M1001_g N_VPWR_c_637_n 0.00585385f $X=7.45 $Y=1.985 $X2=0 $Y2=0
cc_451 N_A_M1004_g N_VPWR_c_638_n 0.00585385f $X=7.87 $Y=1.985 $X2=0 $Y2=0
cc_452 N_A_M1016_g N_VPWR_c_638_n 0.00585385f $X=8.29 $Y=1.985 $X2=0 $Y2=0
cc_453 N_A_M1024_g N_VPWR_c_639_n 0.00585385f $X=8.71 $Y=1.985 $X2=0 $Y2=0
cc_454 N_A_M1001_g N_VPWR_c_632_n 0.010464f $X=7.45 $Y=1.985 $X2=0 $Y2=0
cc_455 N_A_M1004_g N_VPWR_c_632_n 0.0104367f $X=7.87 $Y=1.985 $X2=0 $Y2=0
cc_456 N_A_M1016_g N_VPWR_c_632_n 0.0104367f $X=8.29 $Y=1.985 $X2=0 $Y2=0
cc_457 N_A_M1024_g N_VPWR_c_632_n 0.0114096f $X=8.71 $Y=1.985 $X2=0 $Y2=0
cc_458 N_A_c_561_n N_Y_c_882_n 5.22228e-19 $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_459 N_A_c_561_n N_Y_c_794_n 0.00865686f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_460 N_A_c_565_n N_Y_c_794_n 0.00826974f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_461 N_A_c_561_n N_Y_c_887_n 0.00630972f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_462 N_A_c_562_n N_Y_c_887_n 0.00630972f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_463 N_A_c_563_n N_Y_c_887_n 5.22228e-19 $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_464 N_A_c_562_n N_Y_c_795_n 0.00870364f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_465 N_A_c_563_n N_Y_c_795_n 0.0098365f $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_466 N_A_c_564_n N_Y_c_795_n 0.00262807f $X=8.71 $Y=0.995 $X2=0 $Y2=0
cc_467 N_A_c_565_n N_Y_c_795_n 0.0628716f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_468 N_A_c_566_n N_Y_c_795_n 0.00452472f $X=8.71 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_c_562_n N_Y_c_907_n 5.22228e-19 $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_470 N_A_c_563_n N_Y_c_907_n 0.00630972f $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_471 N_A_c_564_n N_Y_c_907_n 0.00539651f $X=8.71 $Y=0.995 $X2=0 $Y2=0
cc_472 N_A_c_561_n N_Y_c_801_n 0.00113286f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_473 N_A_c_562_n N_Y_c_801_n 0.00113286f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_474 N_A_c_565_n N_Y_c_801_n 0.0266272f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_475 N_A_c_566_n N_Y_c_801_n 0.00230339f $X=8.71 $Y=1.16 $X2=0 $Y2=0
cc_476 N_A_M1001_g N_A_1087_297#_c_1045_n 0.0132131f $X=7.45 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_M1004_g N_A_1087_297#_c_1045_n 0.0132273f $X=7.87 $Y=1.985 $X2=0
+ $Y2=0
cc_478 N_A_c_565_n N_A_1087_297#_c_1045_n 0.0409754f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_c_566_n N_A_1087_297#_c_1045_n 0.00211509f $X=8.71 $Y=1.16 $X2=0
+ $Y2=0
cc_480 N_A_M1016_g N_A_1087_297#_c_1046_n 0.0132714f $X=8.29 $Y=1.985 $X2=0
+ $Y2=0
cc_481 N_A_M1024_g N_A_1087_297#_c_1046_n 0.0135215f $X=8.71 $Y=1.985 $X2=0
+ $Y2=0
cc_482 N_A_c_565_n N_A_1087_297#_c_1046_n 0.041703f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_483 N_A_c_566_n N_A_1087_297#_c_1046_n 0.00211509f $X=8.71 $Y=1.16 $X2=0
+ $Y2=0
cc_484 N_A_c_565_n N_A_1087_297#_c_1047_n 0.0269937f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_485 N_A_c_565_n N_A_1087_297#_c_1049_n 0.0204549f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_486 N_A_c_566_n N_A_1087_297#_c_1049_n 0.00220041f $X=8.71 $Y=1.16 $X2=0
+ $Y2=0
cc_487 N_A_c_561_n N_VGND_c_1112_n 0.00146448f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_488 N_A_c_561_n N_VGND_c_1113_n 0.00423334f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_489 N_A_c_562_n N_VGND_c_1113_n 0.00423334f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_490 N_A_c_562_n N_VGND_c_1114_n 0.00146448f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_491 N_A_c_563_n N_VGND_c_1114_n 0.00146448f $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_492 N_A_c_564_n N_VGND_c_1116_n 0.00366968f $X=8.71 $Y=0.995 $X2=0 $Y2=0
cc_493 N_A_c_565_n N_VGND_c_1116_n 0.0233945f $X=8.62 $Y=1.16 $X2=0 $Y2=0
cc_494 N_A_c_563_n N_VGND_c_1127_n 0.00423334f $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_495 N_A_c_564_n N_VGND_c_1127_n 0.00541359f $X=8.71 $Y=0.995 $X2=0 $Y2=0
cc_496 N_A_c_561_n N_VGND_c_1133_n 0.0057435f $X=7.45 $Y=0.995 $X2=0 $Y2=0
cc_497 N_A_c_562_n N_VGND_c_1133_n 0.0057163f $X=7.87 $Y=0.995 $X2=0 $Y2=0
cc_498 N_A_c_563_n N_VGND_c_1133_n 0.0057163f $X=8.29 $Y=0.995 $X2=0 $Y2=0
cc_499 N_A_c_564_n N_VGND_c_1133_n 0.0104744f $X=8.71 $Y=0.995 $X2=0 $Y2=0
cc_500 N_VPWR_c_632_n N_A_311_297#_M1003_d 0.00209344f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_501 N_VPWR_c_632_n N_A_311_297#_M1008_d 0.00215227f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_632_n N_A_311_297#_M1029_d 0.00215227f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_632_n N_A_311_297#_M1009_d 0.00215203f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_632_n N_A_311_297#_M1030_d 0.0020932f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_633_n N_A_311_297#_c_738_n 0.0075644f $X=0.7 $Y=2.3 $X2=0 $Y2=0
cc_506 N_VPWR_c_637_n N_A_311_297#_c_738_n 0.144936f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_632_n N_A_311_297#_c_738_n 0.0914424f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_637_n N_A_311_297#_c_739_n 0.0510931f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_632_n N_A_311_297#_c_739_n 0.0312418f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_637_n N_A_311_297#_c_769_n 0.0142933f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_632_n N_A_311_297#_c_769_n 0.00962421f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_632_n N_Y_M1003_s 0.00216833f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_c_632_n N_Y_M1023_s 0.00216833f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_514 N_VPWR_c_632_n N_A_729_297#_M1000_s 0.00216833f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_515 N_VPWR_c_632_n N_A_729_297#_M1014_s 0.00216833f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_632_n N_A_729_297#_M1010_d 0.00216833f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_632_n N_A_729_297#_M1031_d 0.00216833f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_632_n N_A_1087_297#_M1010_s 0.0020932f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_519 N_VPWR_c_632_n N_A_1087_297#_M1015_s 0.00215203f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_632_n N_A_1087_297#_M1032_s 0.00246446f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_632_n N_A_1087_297#_M1004_d 0.00284632f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_632_n N_A_1087_297#_M1024_d 0.00260431f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_637_n N_A_1087_297#_c_1050_n 0.0330174f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_632_n N_A_1087_297#_c_1050_n 0.0204627f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_637_n N_A_1087_297#_c_1043_n 0.0198661f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_632_n N_A_1087_297#_c_1043_n 0.0117415f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_637_n N_A_1087_297#_c_1052_n 0.0330174f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_632_n N_A_1087_297#_c_1052_n 0.0204627f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_637_n N_A_1087_297#_c_1077_n 0.0143053f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_632_n N_A_1087_297#_c_1077_n 0.00962794f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_531 N_VPWR_M1001_s N_A_1087_297#_c_1045_n 0.00165831f $X=7.525 $Y=1.485 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_634_n N_A_1087_297#_c_1045_n 0.0126919f $X=7.66 $Y=1.96 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_638_n N_A_1087_297#_c_1081_n 0.0142343f $X=8.375 $Y=2.72 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_632_n N_A_1087_297#_c_1081_n 0.00955092f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_535 N_VPWR_M1016_s N_A_1087_297#_c_1046_n 0.00165831f $X=8.365 $Y=1.485 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_635_n N_A_1087_297#_c_1046_n 0.0126919f $X=8.5 $Y=1.96 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_639_n N_A_1087_297#_c_1048_n 0.0204682f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_632_n N_A_1087_297#_c_1048_n 0.0120542f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_637_n N_A_1087_297#_c_1087_n 0.0142933f $X=7.535 $Y=2.72 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_632_n N_A_1087_297#_c_1087_n 0.00962421f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_541 N_A_311_297#_c_738_n N_Y_M1003_s 0.00316492f $X=3.4 $Y=2.34 $X2=0 $Y2=0
cc_542 N_A_311_297#_c_738_n N_Y_M1023_s 0.00313257f $X=3.4 $Y=2.34 $X2=0 $Y2=0
cc_543 N_A_311_297#_M1008_d N_Y_c_803_n 0.00168993f $X=2.385 $Y=1.485 $X2=0
+ $Y2=0
cc_544 N_A_311_297#_c_753_n N_A_729_297#_M1000_s 0.00312348f $X=4.075 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_545 N_A_311_297#_c_739_n N_A_729_297#_M1014_s 0.00312348f $X=4.915 $Y=2.38
+ $X2=0 $Y2=0
cc_546 N_A_311_297#_M1009_d N_A_729_297#_c_984_n 0.00165831f $X=4.065 $Y=1.485
+ $X2=0 $Y2=0
cc_547 N_A_311_297#_c_753_n N_A_729_297#_c_984_n 0.00320918f $X=4.075 $Y=2.38
+ $X2=0 $Y2=0
cc_548 N_A_311_297#_c_778_p N_A_729_297#_c_984_n 0.0126766f $X=4.2 $Y=1.96 $X2=0
+ $Y2=0
cc_549 N_A_311_297#_c_739_n N_A_729_297#_c_984_n 0.00320918f $X=4.915 $Y=2.38
+ $X2=0 $Y2=0
cc_550 N_A_311_297#_M1030_d N_A_729_297#_c_985_n 0.00277342f $X=4.905 $Y=1.485
+ $X2=0 $Y2=0
cc_551 N_A_311_297#_c_739_n N_A_729_297#_c_985_n 0.00320918f $X=4.915 $Y=2.38
+ $X2=0 $Y2=0
cc_552 N_A_311_297#_c_740_n N_A_729_297#_c_985_n 0.0189421f $X=5.04 $Y=1.96
+ $X2=0 $Y2=0
cc_553 N_A_311_297#_c_753_n N_A_729_297#_c_987_n 0.0118729f $X=4.075 $Y=2.38
+ $X2=0 $Y2=0
cc_554 N_A_311_297#_c_739_n N_A_729_297#_c_988_n 0.0118729f $X=4.915 $Y=2.38
+ $X2=0 $Y2=0
cc_555 N_A_311_297#_c_740_n N_A_1087_297#_c_1042_n 0.0384365f $X=5.04 $Y=1.96
+ $X2=0 $Y2=0
cc_556 N_A_311_297#_c_739_n N_A_1087_297#_c_1043_n 0.0149966f $X=4.915 $Y=2.38
+ $X2=0 $Y2=0
cc_557 N_Y_c_792_n N_A_729_297#_c_985_n 0.00820983f $X=5.815 $Y=0.815 $X2=0
+ $Y2=0
cc_558 N_Y_c_794_n N_A_1087_297#_c_1044_n 0.00936521f $X=7.495 $Y=0.815 $X2=0
+ $Y2=0
cc_559 N_Y_c_794_n N_A_1087_297#_c_1045_n 3.18413e-19 $X=7.495 $Y=0.815 $X2=0
+ $Y2=0
cc_560 N_Y_c_787_n N_VGND_M1019_s 0.00162089f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_561 N_Y_c_790_n N_VGND_M1033_s 0.00162089f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_562 N_Y_c_791_n N_VGND_M1026_d 0.00162089f $X=4.455 $Y=0.815 $X2=0 $Y2=0
cc_563 N_Y_c_792_n N_VGND_M1034_d 0.0108248f $X=5.815 $Y=0.815 $X2=0 $Y2=0
cc_564 N_Y_c_793_n N_VGND_M1006_d 0.00162089f $X=6.655 $Y=0.815 $X2=0 $Y2=0
cc_565 N_Y_c_794_n N_VGND_M1021_d 0.00162089f $X=7.495 $Y=0.815 $X2=0 $Y2=0
cc_566 N_Y_c_795_n N_VGND_M1017_s 0.00162089f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_567 N_Y_c_787_n N_VGND_c_1108_n 0.0122559f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_568 N_Y_c_790_n N_VGND_c_1109_n 0.0122559f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_569 N_Y_c_791_n N_VGND_c_1110_n 0.0122559f $X=4.455 $Y=0.815 $X2=0 $Y2=0
cc_570 N_Y_c_793_n N_VGND_c_1111_n 0.0122559f $X=6.655 $Y=0.815 $X2=0 $Y2=0
cc_571 N_Y_c_794_n N_VGND_c_1112_n 0.0122559f $X=7.495 $Y=0.815 $X2=0 $Y2=0
cc_572 N_Y_c_794_n N_VGND_c_1113_n 0.00198695f $X=7.495 $Y=0.815 $X2=0 $Y2=0
cc_573 N_Y_c_887_n N_VGND_c_1113_n 0.0188551f $X=7.66 $Y=0.39 $X2=0 $Y2=0
cc_574 N_Y_c_795_n N_VGND_c_1113_n 0.00198695f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_575 N_Y_c_795_n N_VGND_c_1114_n 0.0122559f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_576 N_Y_c_795_n N_VGND_c_1116_n 0.00835456f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_577 N_Y_c_804_n N_VGND_c_1117_n 0.0188551f $X=2.1 $Y=0.39 $X2=0 $Y2=0
cc_578 N_Y_c_787_n N_VGND_c_1117_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_579 N_Y_c_787_n N_VGND_c_1119_n 0.00198695f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_580 N_Y_c_818_n N_VGND_c_1119_n 0.0188621f $X=2.94 $Y=0.39 $X2=0 $Y2=0
cc_581 N_Y_c_790_n N_VGND_c_1119_n 9.11858e-19 $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_582 N_Y_c_796_n N_VGND_c_1119_n 0.00118043f $X=2.98 $Y=0.815 $X2=0 $Y2=0
cc_583 N_Y_c_790_n N_VGND_c_1121_n 0.00198695f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_584 N_Y_c_828_n N_VGND_c_1121_n 0.0188551f $X=3.78 $Y=0.39 $X2=0 $Y2=0
cc_585 N_Y_c_791_n N_VGND_c_1121_n 0.00198695f $X=4.455 $Y=0.815 $X2=0 $Y2=0
cc_586 N_Y_c_792_n N_VGND_c_1123_n 0.00198695f $X=5.815 $Y=0.815 $X2=0 $Y2=0
cc_587 N_Y_c_875_n N_VGND_c_1123_n 0.0188551f $X=5.98 $Y=0.39 $X2=0 $Y2=0
cc_588 N_Y_c_793_n N_VGND_c_1123_n 0.00198695f $X=6.655 $Y=0.815 $X2=0 $Y2=0
cc_589 N_Y_c_793_n N_VGND_c_1125_n 0.00198695f $X=6.655 $Y=0.815 $X2=0 $Y2=0
cc_590 N_Y_c_882_n N_VGND_c_1125_n 0.0188551f $X=6.82 $Y=0.39 $X2=0 $Y2=0
cc_591 N_Y_c_794_n N_VGND_c_1125_n 0.00198695f $X=7.495 $Y=0.815 $X2=0 $Y2=0
cc_592 N_Y_c_795_n N_VGND_c_1127_n 0.00198695f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_593 N_Y_c_907_n N_VGND_c_1127_n 0.0188551f $X=8.5 $Y=0.39 $X2=0 $Y2=0
cc_594 N_Y_c_791_n N_VGND_c_1130_n 0.00198695f $X=4.455 $Y=0.815 $X2=0 $Y2=0
cc_595 N_Y_c_859_n N_VGND_c_1130_n 0.0188551f $X=4.62 $Y=0.39 $X2=0 $Y2=0
cc_596 N_Y_c_792_n N_VGND_c_1130_n 0.00198695f $X=5.815 $Y=0.815 $X2=0 $Y2=0
cc_597 N_Y_c_792_n N_VGND_c_1131_n 0.0528344f $X=5.815 $Y=0.815 $X2=0 $Y2=0
cc_598 N_Y_M1012_d N_VGND_c_1133_n 0.00215201f $X=1.965 $Y=0.235 $X2=0 $Y2=0
cc_599 N_Y_M1025_d N_VGND_c_1133_n 0.00215201f $X=2.805 $Y=0.235 $X2=0 $Y2=0
cc_600 N_Y_M1020_s N_VGND_c_1133_n 0.00215201f $X=3.645 $Y=0.235 $X2=0 $Y2=0
cc_601 N_Y_M1027_s N_VGND_c_1133_n 0.00215201f $X=4.485 $Y=0.235 $X2=0 $Y2=0
cc_602 N_Y_M1002_s N_VGND_c_1133_n 0.00215201f $X=5.845 $Y=0.235 $X2=0 $Y2=0
cc_603 N_Y_M1013_s N_VGND_c_1133_n 0.00215201f $X=6.685 $Y=0.235 $X2=0 $Y2=0
cc_604 N_Y_M1007_d N_VGND_c_1133_n 0.00215201f $X=7.525 $Y=0.235 $X2=0 $Y2=0
cc_605 N_Y_M1022_d N_VGND_c_1133_n 0.00215201f $X=8.365 $Y=0.235 $X2=0 $Y2=0
cc_606 N_Y_c_804_n N_VGND_c_1133_n 0.0122069f $X=2.1 $Y=0.39 $X2=0 $Y2=0
cc_607 N_Y_c_787_n N_VGND_c_1133_n 0.00835832f $X=2.775 $Y=0.815 $X2=0 $Y2=0
cc_608 N_Y_c_818_n N_VGND_c_1133_n 0.0122109f $X=2.94 $Y=0.39 $X2=0 $Y2=0
cc_609 N_Y_c_790_n N_VGND_c_1133_n 0.00663839f $X=3.615 $Y=0.815 $X2=0 $Y2=0
cc_610 N_Y_c_828_n N_VGND_c_1133_n 0.0122069f $X=3.78 $Y=0.39 $X2=0 $Y2=0
cc_611 N_Y_c_791_n N_VGND_c_1133_n 0.00835832f $X=4.455 $Y=0.815 $X2=0 $Y2=0
cc_612 N_Y_c_859_n N_VGND_c_1133_n 0.0122069f $X=4.62 $Y=0.39 $X2=0 $Y2=0
cc_613 N_Y_c_792_n N_VGND_c_1133_n 0.0103256f $X=5.815 $Y=0.815 $X2=0 $Y2=0
cc_614 N_Y_c_875_n N_VGND_c_1133_n 0.0122069f $X=5.98 $Y=0.39 $X2=0 $Y2=0
cc_615 N_Y_c_793_n N_VGND_c_1133_n 0.00835832f $X=6.655 $Y=0.815 $X2=0 $Y2=0
cc_616 N_Y_c_882_n N_VGND_c_1133_n 0.0122069f $X=6.82 $Y=0.39 $X2=0 $Y2=0
cc_617 N_Y_c_794_n N_VGND_c_1133_n 0.00835832f $X=7.495 $Y=0.815 $X2=0 $Y2=0
cc_618 N_Y_c_887_n N_VGND_c_1133_n 0.0122069f $X=7.66 $Y=0.39 $X2=0 $Y2=0
cc_619 N_Y_c_795_n N_VGND_c_1133_n 0.00835832f $X=8.335 $Y=0.815 $X2=0 $Y2=0
cc_620 N_Y_c_907_n N_VGND_c_1133_n 0.0122069f $X=8.5 $Y=0.39 $X2=0 $Y2=0
cc_621 N_Y_c_796_n N_VGND_c_1133_n 0.001841f $X=2.98 $Y=0.815 $X2=0 $Y2=0
cc_622 N_A_729_297#_c_985_n N_A_1087_297#_M1010_s 0.00277342f $X=5.855 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_623 N_A_729_297#_c_986_n N_A_1087_297#_M1015_s 0.00165831f $X=6.695 $Y=1.54
+ $X2=0 $Y2=0
cc_624 N_A_729_297#_c_985_n N_A_1087_297#_c_1042_n 0.021051f $X=5.855 $Y=1.54
+ $X2=0 $Y2=0
cc_625 N_A_729_297#_M1010_d N_A_1087_297#_c_1050_n 0.00312348f $X=5.845 $Y=1.485
+ $X2=0 $Y2=0
cc_626 N_A_729_297#_c_985_n N_A_1087_297#_c_1050_n 0.00320918f $X=5.855 $Y=1.54
+ $X2=0 $Y2=0
cc_627 N_A_729_297#_c_986_n N_A_1087_297#_c_1050_n 0.00320918f $X=6.695 $Y=1.54
+ $X2=0 $Y2=0
cc_628 N_A_729_297#_c_989_n N_A_1087_297#_c_1050_n 0.0118729f $X=5.98 $Y=1.62
+ $X2=0 $Y2=0
cc_629 N_A_729_297#_c_986_n N_A_1087_297#_c_1100_n 0.0126766f $X=6.695 $Y=1.54
+ $X2=0 $Y2=0
cc_630 N_A_729_297#_M1031_d N_A_1087_297#_c_1052_n 0.00312348f $X=6.685 $Y=1.485
+ $X2=0 $Y2=0
cc_631 N_A_729_297#_c_986_n N_A_1087_297#_c_1052_n 0.00320918f $X=6.695 $Y=1.54
+ $X2=0 $Y2=0
cc_632 N_A_729_297#_c_990_n N_A_1087_297#_c_1052_n 0.0118729f $X=6.82 $Y=1.62
+ $X2=0 $Y2=0
cc_633 N_A_729_297#_c_990_n N_A_1087_297#_c_1044_n 0.00271526f $X=6.82 $Y=1.62
+ $X2=0 $Y2=0

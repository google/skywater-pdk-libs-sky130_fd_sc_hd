* File: sky130_fd_sc_hd__a221oi_4.spice.SKY130_FD_SC_HD__A221OI_4.pxi
* Created: Thu Aug 27 14:02:12 2020
* 
x_PM_SKY130_FD_SC_HD__A221OI_4%C1 N_C1_c_127_n N_C1_M1014_g N_C1_M1011_g
+ N_C1_c_128_n N_C1_M1019_g N_C1_M1030_g N_C1_c_129_n N_C1_M1027_g N_C1_M1033_g
+ N_C1_c_130_n N_C1_M1028_g N_C1_M1037_g C1 N_C1_c_132_n
+ PM_SKY130_FD_SC_HD__A221OI_4%C1
x_PM_SKY130_FD_SC_HD__A221OI_4%B2 N_B2_c_207_n N_B2_M1000_g N_B2_c_208_n
+ N_B2_M1009_g N_B2_M1002_g N_B2_c_209_n N_B2_M1012_g N_B2_M1007_g N_B2_M1023_g
+ N_B2_c_210_n N_B2_M1025_g N_B2_M1026_g N_B2_c_211_n N_B2_c_212_n N_B2_c_213_n
+ N_B2_c_222_n B2 N_B2_c_214_n PM_SKY130_FD_SC_HD__A221OI_4%B2
x_PM_SKY130_FD_SC_HD__A221OI_4%B1 N_B1_c_331_n N_B1_M1004_g N_B1_M1008_g
+ N_B1_c_332_n N_B1_M1015_g N_B1_M1013_g N_B1_c_333_n N_B1_M1017_g N_B1_M1034_g
+ N_B1_c_334_n N_B1_M1020_g N_B1_M1038_g B1 N_B1_c_335_n N_B1_c_336_n
+ PM_SKY130_FD_SC_HD__A221OI_4%B1
x_PM_SKY130_FD_SC_HD__A221OI_4%A2 N_A2_c_395_n N_A2_M1005_g N_A2_M1016_g
+ N_A2_c_396_n N_A2_M1018_g N_A2_M1024_g N_A2_c_397_n N_A2_M1022_g N_A2_M1031_g
+ N_A2_c_398_n N_A2_M1029_g N_A2_M1036_g N_A2_c_399_n N_A2_c_400_n N_A2_c_411_n
+ N_A2_c_412_n N_A2_c_401_n N_A2_c_402_n A2 N_A2_c_403_n N_A2_c_404_n
+ PM_SKY130_FD_SC_HD__A221OI_4%A2
x_PM_SKY130_FD_SC_HD__A221OI_4%A1 N_A1_c_521_n N_A1_M1001_g N_A1_M1003_g
+ N_A1_c_522_n N_A1_M1006_g N_A1_M1032_g N_A1_c_523_n N_A1_M1010_g N_A1_M1035_g
+ N_A1_c_524_n N_A1_M1021_g N_A1_M1039_g A1 N_A1_c_539_n N_A1_c_525_n
+ PM_SKY130_FD_SC_HD__A221OI_4%A1
x_PM_SKY130_FD_SC_HD__A221OI_4%A_27_297# N_A_27_297#_M1011_s N_A_27_297#_M1030_s
+ N_A_27_297#_M1037_s N_A_27_297#_M1002_s N_A_27_297#_M1023_s
+ N_A_27_297#_M1013_d N_A_27_297#_M1038_d N_A_27_297#_c_579_n
+ N_A_27_297#_c_580_n N_A_27_297#_c_588_n N_A_27_297#_c_619_p
+ N_A_27_297#_c_590_n N_A_27_297#_c_581_n N_A_27_297#_c_582_n
+ N_A_27_297#_c_583_n N_A_27_297#_c_584_n N_A_27_297#_c_603_n
+ N_A_27_297#_c_604_n N_A_27_297#_c_605_n N_A_27_297#_c_652_p
+ PM_SKY130_FD_SC_HD__A221OI_4%A_27_297#
x_PM_SKY130_FD_SC_HD__A221OI_4%Y N_Y_M1014_d N_Y_M1027_d N_Y_M1004_d N_Y_M1017_d
+ N_Y_M1001_d N_Y_M1010_d N_Y_M1011_d N_Y_M1033_d N_Y_c_671_n N_Y_c_750_n
+ N_Y_c_667_n N_Y_c_668_n N_Y_c_658_n N_Y_c_659_n N_Y_c_689_n N_Y_c_754_n
+ N_Y_c_660_n N_Y_c_661_n N_Y_c_662_n N_Y_c_714_n N_Y_c_734_n N_Y_c_663_n
+ N_Y_c_669_n N_Y_c_670_n N_Y_c_716_n N_Y_c_664_n N_Y_c_665_n N_Y_c_666_n Y
+ PM_SKY130_FD_SC_HD__A221OI_4%Y
x_PM_SKY130_FD_SC_HD__A221OI_4%A_471_297# N_A_471_297#_M1002_d
+ N_A_471_297#_M1007_d N_A_471_297#_M1008_s N_A_471_297#_M1034_s
+ N_A_471_297#_M1026_d N_A_471_297#_M1003_d N_A_471_297#_M1035_d
+ N_A_471_297#_M1024_s N_A_471_297#_M1036_s N_A_471_297#_c_808_n
+ N_A_471_297#_c_809_n N_A_471_297#_c_815_n N_A_471_297#_c_820_n
+ N_A_471_297#_c_889_p N_A_471_297#_c_829_n N_A_471_297#_c_874_p
+ N_A_471_297#_c_834_n N_A_471_297#_c_810_n N_A_471_297#_c_811_n
+ N_A_471_297#_c_879_p N_A_471_297#_c_846_n
+ PM_SKY130_FD_SC_HD__A221OI_4%A_471_297#
x_PM_SKY130_FD_SC_HD__A221OI_4%VPWR N_VPWR_M1016_d N_VPWR_M1032_s N_VPWR_M1039_s
+ N_VPWR_M1031_d N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_901_n VPWR
+ N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_898_n N_VPWR_c_906_n
+ N_VPWR_c_907_n PM_SKY130_FD_SC_HD__A221OI_4%VPWR
x_PM_SKY130_FD_SC_HD__A221OI_4%VGND N_VGND_M1014_s N_VGND_M1019_s N_VGND_M1028_s
+ N_VGND_M1009_s N_VGND_M1025_s N_VGND_M1018_s N_VGND_M1029_s N_VGND_c_1003_n
+ N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n
+ N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n
+ N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n
+ N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n VGND N_VGND_c_1023_n
+ N_VGND_c_1024_n PM_SKY130_FD_SC_HD__A221OI_4%VGND
x_PM_SKY130_FD_SC_HD__A221OI_4%A_453_47# N_A_453_47#_M1000_d N_A_453_47#_M1012_d
+ N_A_453_47#_M1015_s N_A_453_47#_M1020_s N_A_453_47#_c_1141_n
+ N_A_453_47#_c_1143_n N_A_453_47#_c_1144_n N_A_453_47#_c_1146_n
+ PM_SKY130_FD_SC_HD__A221OI_4%A_453_47#
x_PM_SKY130_FD_SC_HD__A221OI_4%A_1241_47# N_A_1241_47#_M1005_d
+ N_A_1241_47#_M1006_s N_A_1241_47#_M1021_s N_A_1241_47#_M1022_d
+ N_A_1241_47#_c_1179_n N_A_1241_47#_c_1180_n N_A_1241_47#_c_1177_n
+ N_A_1241_47#_c_1178_n N_A_1241_47#_c_1191_n
+ PM_SKY130_FD_SC_HD__A221OI_4%A_1241_47#
cc_1 VNB N_C1_c_127_n 0.0216231f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_C1_c_128_n 0.0157805f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_C1_c_129_n 0.015776f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_C1_c_130_n 0.0159359f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB C1 0.0134887f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_6 VNB N_C1_c_132_n 0.0765267f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_B2_c_207_n 0.0159991f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B2_c_208_n 0.0156317f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_9 VNB N_B2_c_209_n 0.0199271f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.325
cc_10 VNB N_B2_c_210_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_11 VNB N_B2_c_211_n 0.00356333f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_12 VNB N_B2_c_212_n 0.0192987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B2_c_213_n 0.00525539f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_14 VNB N_B2_c_214_n 0.0775185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_331_n 0.0202009f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_16 VNB N_B1_c_332_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_17 VNB N_B1_c_333_n 0.0160051f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_18 VNB N_B1_c_334_n 0.0162456f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_19 VNB N_B1_c_335_n 0.00219191f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_20 VNB N_B1_c_336_n 0.061908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A2_c_395_n 0.0169414f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_22 VNB N_A2_c_396_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_23 VNB N_A2_c_397_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_24 VNB N_A2_c_398_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_25 VNB N_A2_c_399_n 0.00351686f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_26 VNB N_A2_c_400_n 0.0193115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A2_c_401_n 2.86539e-19 $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.16
cc_28 VNB N_A2_c_402_n 0.00189815f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.16
cc_29 VNB N_A2_c_403_n 0.0266502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A2_c_404_n 0.0569029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A1_c_521_n 0.016243f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_32 VNB N_A1_c_522_n 0.0160042f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_33 VNB N_A1_c_523_n 0.0160044f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_34 VNB N_A1_c_524_n 0.0162429f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_35 VNB N_A1_c_525_n 0.0642393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_658_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_37 VNB N_Y_c_659_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.16
cc_38 VNB N_Y_c_660_n 8.37691e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_661_n 0.00786616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_662_n 0.00157832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_663_n 0.0012664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_664_n 4.77184e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_665_n 0.00770891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_666_n 0.00270091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VPWR_c_898_n 0.402575f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_46 VNB N_VGND_c_1003_n 0.0106747f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_47 VNB N_VGND_c_1004_n 0.0311064f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_48 VNB N_VGND_c_1005_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_1006_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_50 VNB N_VGND_c_1007_n 0.00188409f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_51 VNB N_VGND_c_1008_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.16
cc_52 VNB N_VGND_c_1009_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.175
cc_53 VNB N_VGND_c_1010_n 0.0066043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1011_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1012_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1013_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1014_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1015_n 0.00153094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1016_n 0.00328829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1017_n 0.0863072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1018_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1019_n 0.0538896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1020_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1021_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1022_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1023_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1024_n 0.454569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1241_47#_c_1177_n 0.00325721f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_69 VNB N_A_1241_47#_c_1178_n 0.00440603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VPB N_C1_M1011_g 0.0249346f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_71 VPB N_C1_M1030_g 0.0181173f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_72 VPB N_C1_M1033_g 0.0180886f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_73 VPB N_C1_M1037_g 0.0242555f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_74 VPB N_C1_c_132_n 0.0138546f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_75 VPB N_B2_M1002_g 0.0250398f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.56
cc_76 VPB N_B2_M1007_g 0.0184839f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_77 VPB N_B2_M1023_g 0.017892f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_78 VPB N_B2_M1026_g 0.0181129f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_79 VPB N_B2_c_211_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_80 VPB N_B2_c_212_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_B2_c_213_n 0.00131588f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_82 VPB N_B2_c_222_n 0.01147f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_83 VPB N_B2_c_214_n 0.0223547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_B1_M1008_g 0.0183505f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_85 VPB N_B1_M1013_g 0.0181176f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_86 VPB N_B1_M1034_g 0.018119f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_87 VPB N_B1_M1038_g 0.0183572f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_88 VPB N_B1_c_336_n 0.0100566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A2_M1016_g 0.0178693f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_90 VPB N_A2_M1024_g 0.0176172f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_91 VPB N_A2_M1031_g 0.0181197f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_92 VPB N_A2_M1036_g 0.025044f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_93 VPB N_A2_c_399_n 0.00233749f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_94 VPB N_A2_c_400_n 0.00443023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A2_c_411_n 0.0133611f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_96 VPB N_A2_c_412_n 2.50157e-19 $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_97 VPB N_A2_c_401_n 0.00137341f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.16
cc_98 VPB N_A2_c_404_n 0.00910688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A1_M1003_g 0.0174125f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_100 VPB N_A1_M1032_g 0.0172192f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_101 VPB N_A1_M1035_g 0.0172196f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_102 VPB N_A1_M1039_g 0.0174156f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_103 VPB N_A1_c_525_n 0.0100821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_27_297#_c_579_n 0.00753428f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.995
cc_105 VPB N_A_27_297#_c_580_n 0.0360467f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_106 VPB N_A_27_297#_c_581_n 0.00181613f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_107 VPB N_A_27_297#_c_582_n 0.00652951f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.16
cc_108 VPB N_A_27_297#_c_583_n 0.013847f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.16
cc_109 VPB N_A_27_297#_c_584_n 0.00300568f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_110 VPB N_Y_c_667_n 0.00238525f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_111 VPB N_Y_c_668_n 0.00234506f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_112 VPB N_Y_c_669_n 0.00112006f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_Y_c_670_n 0.00112172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_471_297#_c_808_n 0.0025234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_471_297#_c_809_n 0.00400507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_471_297#_c_810_n 0.00619863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_471_297#_c_811_n 0.00138022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_899_n 0.00410258f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.995
cc_119 VPB N_VPWR_c_900_n 0.0150303f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_120 VPB N_VPWR_c_901_n 0.00324402f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_121 VPB N_VPWR_c_902_n 0.0188097f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_122 VPB N_VPWR_c_903_n 0.00417211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_904_n 0.0225629f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.16
cc_124 VPB N_VPWR_c_898_n 0.0586236f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_125 VPB N_VPWR_c_906_n 0.141577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_907_n 0.00408644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 N_C1_c_130_n N_B2_c_207_n 0.0191323f $X=1.75 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_128 N_C1_c_132_n N_B2_c_214_n 0.0191323f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C1_M1011_g N_A_27_297#_c_580_n 9.42064e-19 $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_130 C1 N_A_27_297#_c_580_n 0.0264267f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_131 N_C1_c_132_n N_A_27_297#_c_580_n 0.00195514f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_132 N_C1_M1011_g N_A_27_297#_c_588_n 0.0121747f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C1_M1030_g N_A_27_297#_c_588_n 0.0121747f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C1_M1033_g N_A_27_297#_c_590_n 0.0121747f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C1_M1037_g N_A_27_297#_c_590_n 0.0121747f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_136 N_C1_M1037_g N_A_27_297#_c_584_n 9.22601e-19 $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_137 N_C1_c_127_n N_Y_c_671_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C1_c_128_n N_Y_c_671_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C1_c_129_n N_Y_c_671_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C1_M1030_g N_Y_c_667_n 0.0133089f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_141 N_C1_M1033_g N_Y_c_667_n 0.0141417f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_142 C1 N_Y_c_667_n 0.0360189f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_143 N_C1_c_132_n N_Y_c_667_n 0.00214031f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_144 N_C1_M1011_g N_Y_c_668_n 3.45391e-19 $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_145 C1 N_Y_c_668_n 0.0203891f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_146 N_C1_c_132_n N_Y_c_668_n 0.00222344f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_147 N_C1_c_128_n N_Y_c_658_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_148 N_C1_c_129_n N_Y_c_658_n 0.00914727f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_149 C1 N_Y_c_658_n 0.0333876f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_150 N_C1_c_132_n N_Y_c_658_n 0.00222133f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_151 N_C1_c_127_n N_Y_c_659_n 0.00299247f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_152 N_C1_c_128_n N_Y_c_659_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_153 C1 N_Y_c_659_n 0.0265405f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_154 N_C1_c_132_n N_Y_c_659_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_155 N_C1_c_128_n N_Y_c_689_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_156 N_C1_c_129_n N_Y_c_689_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_157 N_C1_c_130_n N_Y_c_689_n 0.00513001f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_158 N_C1_c_129_n N_Y_c_660_n 0.00205955f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_159 N_C1_c_130_n N_Y_c_660_n 0.00210394f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_160 C1 N_Y_c_660_n 0.0014288f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_161 N_C1_c_132_n N_Y_c_660_n 0.00919607f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_162 N_C1_c_132_n N_Y_c_661_n 0.0147834f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_163 N_C1_c_129_n N_Y_c_663_n 0.00144031f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C1_c_130_n N_Y_c_663_n 0.00210928f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C1_c_132_n N_Y_c_663_n 3.16161e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_166 N_C1_M1033_g N_Y_c_669_n 0.00275378f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_167 N_C1_M1037_g N_Y_c_669_n 0.00579852f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_168 N_C1_c_132_n N_Y_c_669_n 0.00581264f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_169 N_C1_M1037_g N_Y_c_670_n 0.00378071f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_170 N_C1_c_132_n N_Y_c_670_n 3.04645e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_171 C1 Y 0.0151525f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_172 N_C1_c_132_n Y 0.00597684f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_173 N_C1_M1011_g N_VPWR_c_898_n 0.00619805f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_174 N_C1_M1030_g N_VPWR_c_898_n 0.00522516f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_175 N_C1_M1033_g N_VPWR_c_898_n 0.00522516f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_176 N_C1_M1037_g N_VPWR_c_898_n 0.00655123f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_177 N_C1_M1011_g N_VPWR_c_906_n 0.00357877f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_178 N_C1_M1030_g N_VPWR_c_906_n 0.00357877f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_179 N_C1_M1033_g N_VPWR_c_906_n 0.00357877f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_180 N_C1_M1037_g N_VPWR_c_906_n 0.00357877f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_181 N_C1_c_127_n N_VGND_c_1004_n 0.00343277f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_182 C1 N_VGND_c_1004_n 0.020187f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_183 N_C1_c_132_n N_VGND_c_1004_n 9.96531e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_184 N_C1_c_128_n N_VGND_c_1005_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_185 N_C1_c_129_n N_VGND_c_1005_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_186 N_C1_c_130_n N_VGND_c_1006_n 0.00175763f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_187 N_C1_c_130_n N_VGND_c_1007_n 0.00138226f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_188 N_C1_c_127_n N_VGND_c_1011_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_189 N_C1_c_128_n N_VGND_c_1011_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_190 N_C1_c_129_n N_VGND_c_1013_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_191 N_C1_c_130_n N_VGND_c_1013_n 0.00541359f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_192 N_C1_c_127_n N_VGND_c_1024_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_193 N_C1_c_128_n N_VGND_c_1024_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_194 N_C1_c_129_n N_VGND_c_1024_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_195 N_C1_c_130_n N_VGND_c_1024_n 0.00957732f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B2_M1023_g N_B1_M1008_g 0.0437142f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B2_c_222_n N_B1_M1008_g 0.0114737f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_198 N_B2_c_222_n N_B1_M1013_g 0.0106666f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_199 N_B2_c_222_n N_B1_M1034_g 0.0106666f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_200 N_B2_c_210_n N_B1_c_334_n 0.0265533f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B2_M1026_g N_B1_M1038_g 0.043506f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B2_c_222_n N_B1_M1038_g 0.0106225f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_203 N_B2_c_211_n N_B1_c_335_n 0.0159907f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B2_c_212_n N_B1_c_335_n 7.8248e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B2_c_213_n N_B1_c_335_n 0.0235459f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_206 N_B2_c_222_n N_B1_c_335_n 0.0981881f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_207 N_B2_c_214_n N_B1_c_335_n 2.46885e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B2_c_211_n N_B1_c_336_n 0.00461956f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B2_c_212_n N_B1_c_336_n 0.0213293f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_210 N_B2_c_213_n N_B1_c_336_n 0.00615921f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_211 N_B2_c_222_n N_B1_c_336_n 0.00642092f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_212 N_B2_c_214_n N_B1_c_336_n 0.0183261f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B2_c_210_n N_A2_c_395_n 0.0245777f $X=5.63 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_214 N_B2_M1026_g N_A2_M1016_g 0.02101f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B2_c_211_n N_A2_M1016_g 3.59226e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_216 N_B2_c_222_n N_A2_M1016_g 5.77655e-19 $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_217 N_B2_M1026_g N_A2_c_399_n 3.59226e-19 $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_218 N_B2_c_211_n N_A2_c_399_n 0.0307171f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B2_c_212_n N_A2_c_399_n 7.80994e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B2_c_211_n N_A2_c_400_n 7.80994e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B2_c_212_n N_A2_c_400_n 0.0197715f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B2_M1026_g N_A2_c_412_n 5.77655e-19 $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_223 N_B2_c_222_n N_A2_c_412_n 0.0154679f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_224 N_B2_c_213_n N_A_27_297#_M1023_s 0.00127619f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_225 N_B2_c_222_n N_A_27_297#_M1023_s 6.19991e-19 $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_226 N_B2_c_222_n N_A_27_297#_M1013_d 0.00185997f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_227 N_B2_c_222_n N_A_27_297#_M1038_d 0.00184938f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_228 N_B2_M1002_g N_A_27_297#_c_582_n 0.00317531f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_229 N_B2_M1002_g N_A_27_297#_c_583_n 0.0120804f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_230 N_B2_M1007_g N_A_27_297#_c_583_n 6.46788e-19 $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_231 N_B2_c_213_n N_A_27_297#_c_583_n 0.00343816f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B2_c_214_n N_A_27_297#_c_583_n 0.0158623f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B2_c_214_n N_A_27_297#_c_584_n 2.89127e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B2_M1002_g N_A_27_297#_c_603_n 0.00273231f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_235 N_B2_M1002_g N_A_27_297#_c_604_n 0.00427937f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_236 N_B2_M1007_g N_A_27_297#_c_605_n 0.0113231f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_237 N_B2_M1023_g N_A_27_297#_c_605_n 0.0110426f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_238 N_B2_M1026_g N_A_27_297#_c_605_n 0.00305585f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_239 N_B2_c_213_n N_A_27_297#_c_605_n 0.0123254f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B2_c_222_n N_A_27_297#_c_605_n 0.076777f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_241 N_B2_c_214_n N_A_27_297#_c_605_n 0.00242248f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B2_c_207_n N_Y_c_660_n 9.42752e-19 $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B2_c_213_n N_Y_c_661_n 0.0145048f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_244 N_B2_c_214_n N_Y_c_661_n 0.0523748f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B2_c_208_n N_Y_c_662_n 3.97882e-19 $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B2_c_209_n N_Y_c_662_n 0.00526285f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B2_c_213_n N_Y_c_662_n 0.00717854f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B2_c_214_n N_Y_c_662_n 0.0101555f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B2_c_209_n N_Y_c_714_n 0.0064824f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B2_c_214_n N_Y_c_669_n 2.91589e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B2_c_211_n N_Y_c_716_n 0.00229281f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B2_c_212_n N_Y_c_716_n 3.11223e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_253 N_B2_c_213_n N_Y_c_716_n 0.0266645f $X=3.5 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B2_c_222_n N_Y_c_716_n 0.00818214f $X=5.465 $Y=1.53 $X2=0 $Y2=0
cc_255 N_B2_c_214_n N_Y_c_716_n 0.00819446f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B2_c_210_n N_Y_c_664_n 0.0109527f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B2_c_211_n N_Y_c_664_n 0.022216f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B2_c_212_n N_Y_c_664_n 0.00112038f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B2_c_210_n N_Y_c_665_n 0.00366075f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_260 N_B2_c_212_n N_Y_c_665_n 0.001478f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B2_c_222_n N_A_471_297#_M1008_s 0.00185997f $X=5.465 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_B2_c_222_n N_A_471_297#_M1034_s 0.00185997f $X=5.465 $Y=1.53 $X2=0
+ $Y2=0
cc_263 N_B2_c_222_n N_A_471_297#_M1026_d 0.00151125f $X=5.465 $Y=1.53 $X2=0
+ $Y2=0
cc_264 N_B2_M1002_g N_A_471_297#_c_815_n 0.0113556f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B2_M1007_g N_A_471_297#_c_815_n 0.00970685f $X=3.11 $Y=1.985 $X2=0
+ $Y2=0
cc_266 N_B2_M1023_g N_A_471_297#_c_815_n 0.00964167f $X=3.53 $Y=1.985 $X2=0
+ $Y2=0
cc_267 N_B2_M1026_g N_A_471_297#_c_815_n 0.0112888f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B2_c_222_n N_A_471_297#_c_815_n 0.00322464f $X=5.465 $Y=1.53 $X2=0
+ $Y2=0
cc_269 N_B2_c_222_n N_A_471_297#_c_820_n 0.00292685f $X=5.465 $Y=1.53 $X2=0
+ $Y2=0
cc_270 N_B2_M1026_g N_VPWR_c_903_n 0.00104358f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B2_M1002_g N_VPWR_c_898_n 0.00655123f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B2_M1007_g N_VPWR_c_898_n 0.00522516f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B2_M1023_g N_VPWR_c_898_n 0.00525341f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B2_M1026_g N_VPWR_c_898_n 0.00546478f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B2_M1002_g N_VPWR_c_906_n 0.00357877f $X=2.69 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B2_M1007_g N_VPWR_c_906_n 0.00357877f $X=3.11 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B2_M1023_g N_VPWR_c_906_n 0.00357877f $X=3.53 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B2_M1026_g N_VPWR_c_906_n 0.00357877f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B2_c_207_n N_VGND_c_1006_n 0.00715825f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B2_c_210_n N_VGND_c_1008_n 0.00633616f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B2_c_209_n N_VGND_c_1015_n 3.09187e-19 $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B2_c_214_n N_VGND_c_1015_n 0.00266361f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B2_c_207_n N_VGND_c_1016_n 0.0150328f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B2_c_208_n N_VGND_c_1016_n 0.0116864f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B2_c_214_n N_VGND_c_1016_n 0.00230169f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_286 N_B2_c_207_n N_VGND_c_1017_n 0.00412827f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_208_n N_VGND_c_1017_n 0.00357877f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_209_n N_VGND_c_1017_n 0.00357877f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B2_c_210_n N_VGND_c_1017_n 0.00414934f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B2_c_207_n N_VGND_c_1024_n 0.00569493f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B2_c_208_n N_VGND_c_1024_n 0.00522516f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_209_n N_VGND_c_1024_n 0.00655123f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B2_c_210_n N_VGND_c_1024_n 0.00601858f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B2_c_209_n N_A_453_47#_c_1141_n 0.00412709f $X=3.03 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_B2_c_214_n N_A_453_47#_c_1141_n 6.24525e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_296 N_B2_c_210_n N_A_453_47#_c_1143_n 0.00337161f $X=5.63 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_B2_c_207_n N_A_453_47#_c_1144_n 0.00304268f $X=2.19 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_B2_c_208_n N_A_453_47#_c_1144_n 0.00376612f $X=2.61 $Y=0.995 $X2=0
+ $Y2=0
cc_299 N_B2_c_208_n N_A_453_47#_c_1146_n 0.00491253f $X=2.61 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_B2_c_209_n N_A_453_47#_c_1146_n 0.00615568f $X=3.03 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_B1_M1008_g N_A_27_297#_c_605_n 0.00972403f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_302 N_B1_M1013_g N_A_27_297#_c_605_n 0.00972403f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_303 N_B1_M1034_g N_A_27_297#_c_605_n 0.00972403f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_304 N_B1_M1038_g N_A_27_297#_c_605_n 0.00972403f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_305 N_B1_c_331_n N_Y_c_662_n 0.00370094f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_331_n N_Y_c_716_n 0.0115279f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_c_332_n N_Y_c_716_n 0.00852218f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_308 N_B1_c_333_n N_Y_c_716_n 0.00852218f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_c_334_n N_Y_c_716_n 0.00847671f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B1_c_335_n N_Y_c_716_n 0.082793f $X=5.12 $Y=1.16 $X2=0 $Y2=0
cc_311 N_B1_c_336_n N_Y_c_716_n 0.00603821f $X=5.21 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B1_c_334_n N_Y_c_664_n 6.55089e-19 $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_M1008_g N_A_471_297#_c_815_n 0.00964167f $X=3.95 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_B1_M1013_g N_A_471_297#_c_815_n 0.00970685f $X=4.37 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_B1_M1034_g N_A_471_297#_c_815_n 0.00970685f $X=4.79 $Y=1.985 $X2=0
+ $Y2=0
cc_316 N_B1_M1038_g N_A_471_297#_c_815_n 0.00964167f $X=5.21 $Y=1.985 $X2=0
+ $Y2=0
cc_317 N_B1_M1008_g N_VPWR_c_898_n 0.00525341f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_318 N_B1_M1013_g N_VPWR_c_898_n 0.00522516f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_319 N_B1_M1034_g N_VPWR_c_898_n 0.00522516f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_320 N_B1_M1038_g N_VPWR_c_898_n 0.00525341f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_321 N_B1_M1008_g N_VPWR_c_906_n 0.00357877f $X=3.95 $Y=1.985 $X2=0 $Y2=0
cc_322 N_B1_M1013_g N_VPWR_c_906_n 0.00357877f $X=4.37 $Y=1.985 $X2=0 $Y2=0
cc_323 N_B1_M1034_g N_VPWR_c_906_n 0.00357877f $X=4.79 $Y=1.985 $X2=0 $Y2=0
cc_324 N_B1_M1038_g N_VPWR_c_906_n 0.00357877f $X=5.21 $Y=1.985 $X2=0 $Y2=0
cc_325 N_B1_c_331_n N_VGND_c_1017_n 0.00357877f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B1_c_332_n N_VGND_c_1017_n 0.00357877f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B1_c_333_n N_VGND_c_1017_n 0.00357877f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B1_c_334_n N_VGND_c_1017_n 0.00357877f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_c_331_n N_VGND_c_1024_n 0.00655123f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_330 N_B1_c_332_n N_VGND_c_1024_n 0.00522516f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B1_c_333_n N_VGND_c_1024_n 0.00522516f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B1_c_334_n N_VGND_c_1024_n 0.00525237f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B1_c_331_n N_A_453_47#_c_1143_n 0.00892725f $X=3.95 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_B1_c_332_n N_A_453_47#_c_1143_n 0.00892725f $X=4.37 $Y=0.995 $X2=0
+ $Y2=0
cc_335 N_B1_c_333_n N_A_453_47#_c_1143_n 0.00892725f $X=4.79 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_B1_c_334_n N_A_453_47#_c_1143_n 0.00892725f $X=5.21 $Y=0.995 $X2=0
+ $Y2=0
cc_337 N_A2_c_395_n N_A1_c_521_n 0.0260114f $X=6.13 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_338 N_A2_M1016_g N_A1_M1003_g 0.0432959f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A2_c_411_n N_A1_M1003_g 0.0103037f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_340 N_A2_c_411_n N_A1_M1032_g 0.0103615f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_341 N_A2_c_411_n N_A1_M1035_g 0.0103615f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_342 N_A2_c_396_n N_A1_c_524_n 0.0241518f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A2_M1024_g N_A1_M1039_g 0.0241518f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A2_c_411_n N_A1_M1039_g 0.0103037f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_345 N_A2_c_399_n N_A1_c_539_n 0.0160038f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A2_c_400_n N_A1_c_539_n 2.34877e-19 $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A2_c_411_n N_A1_c_539_n 0.100214f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_348 N_A2_c_402_n N_A1_c_539_n 0.0151431f $X=8.265 $Y=1.175 $X2=0 $Y2=0
cc_349 N_A2_c_404_n N_A1_c_539_n 2.26155e-19 $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_350 N_A2_c_399_n N_A1_c_525_n 0.00518416f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A2_c_400_n N_A1_c_525_n 0.0228076f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A2_c_411_n N_A1_c_525_n 0.00641737f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_353 N_A2_c_401_n N_A1_c_525_n 0.00336014f $X=8.18 $Y=1.445 $X2=0 $Y2=0
cc_354 N_A2_c_402_n N_A1_c_525_n 0.001542f $X=8.265 $Y=1.175 $X2=0 $Y2=0
cc_355 N_A2_c_404_n N_A1_c_525_n 0.0241518f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_356 N_A2_c_411_n N_Y_c_734_n 2.51155e-19 $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_357 N_A2_c_395_n N_Y_c_664_n 3.31489e-19 $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A2_c_395_n N_Y_c_665_n 0.0120815f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A2_c_399_n N_Y_c_665_n 0.025402f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_360 N_A2_c_400_n N_Y_c_665_n 0.00295599f $X=6.13 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A2_c_395_n N_Y_c_666_n 0.00130466f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A2_c_411_n N_Y_c_666_n 0.00574656f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_363 N_A2_c_412_n N_A_471_297#_M1026_d 0.00151125f $X=6.295 $Y=1.53 $X2=0
+ $Y2=0
cc_364 N_A2_c_411_n N_A_471_297#_M1003_d 0.00166235f $X=8.095 $Y=1.53 $X2=0
+ $Y2=0
cc_365 N_A2_c_411_n N_A_471_297#_M1035_d 0.00166235f $X=8.095 $Y=1.53 $X2=0
+ $Y2=0
cc_366 N_A2_c_412_n N_A_471_297#_c_820_n 0.00292685f $X=6.295 $Y=1.53 $X2=0
+ $Y2=0
cc_367 N_A2_M1016_g N_A_471_297#_c_829_n 0.0118822f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A2_M1024_g N_A_471_297#_c_829_n 0.0123215f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A2_c_411_n N_A_471_297#_c_829_n 0.106315f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_370 N_A2_c_412_n N_A_471_297#_c_829_n 0.0142323f $X=6.295 $Y=1.53 $X2=0 $Y2=0
cc_371 N_A2_c_403_n N_A_471_297#_c_829_n 0.00183652f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_372 N_A2_M1024_g N_A_471_297#_c_834_n 0.00356696f $X=8.23 $Y=1.985 $X2=0
+ $Y2=0
cc_373 N_A2_M1031_g N_A_471_297#_c_834_n 0.0040777f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A2_M1036_g N_A_471_297#_c_834_n 4.65489e-19 $X=9.07 $Y=1.985 $X2=0
+ $Y2=0
cc_375 N_A2_M1031_g N_A_471_297#_c_810_n 0.0106747f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A2_M1036_g N_A_471_297#_c_810_n 0.0136443f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_377 N_A2_c_403_n N_A_471_297#_c_810_n 0.0599466f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A2_c_404_n N_A_471_297#_c_810_n 0.00324189f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A2_M1024_g N_A_471_297#_c_811_n 0.0011544f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_380 N_A2_M1031_g N_A_471_297#_c_811_n 0.002092f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_381 N_A2_c_411_n N_A_471_297#_c_811_n 0.0149285f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_382 N_A2_c_403_n N_A_471_297#_c_811_n 0.0136617f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A2_c_404_n N_A_471_297#_c_811_n 0.00123743f $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_384 N_A2_M1031_g N_A_471_297#_c_846_n 0.00349558f $X=8.65 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_A2_c_403_n N_A_471_297#_c_846_n 0.00258233f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_386 N_A2_c_404_n N_A_471_297#_c_846_n 7.86192e-19 $X=9.07 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A2_c_411_n N_VPWR_M1016_d 0.00130005f $X=8.095 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_388 N_A2_c_412_n N_VPWR_M1016_d 3.52503e-19 $X=6.295 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_389 N_A2_c_411_n N_VPWR_M1032_s 0.00166235f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_390 N_A2_c_411_n N_VPWR_M1039_s 0.00161973f $X=8.095 $Y=1.53 $X2=0 $Y2=0
cc_391 N_A2_M1031_g N_VPWR_c_899_n 0.00137298f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A2_M1036_g N_VPWR_c_899_n 0.00268723f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A2_M1024_g N_VPWR_c_900_n 0.00343969f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A2_M1031_g N_VPWR_c_900_n 0.00554458f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_395 N_A2_M1016_g N_VPWR_c_903_n 0.00834127f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_396 N_A2_M1036_g N_VPWR_c_904_n 0.00585385f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A2_M1016_g N_VPWR_c_898_n 0.00421719f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A2_M1024_g N_VPWR_c_898_n 0.00400583f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_399 N_A2_M1031_g N_VPWR_c_898_n 0.00960147f $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A2_M1036_g N_VPWR_c_898_n 0.0115882f $X=9.07 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A2_M1016_g N_VPWR_c_906_n 0.00343969f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A2_M1024_g N_VPWR_c_907_n 0.00725667f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_403 N_A2_M1031_g N_VPWR_c_907_n 5.72916e-19 $X=8.65 $Y=1.985 $X2=0 $Y2=0
cc_404 N_A2_c_395_n N_VGND_c_1008_n 0.00280412f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A2_c_396_n N_VGND_c_1009_n 0.00268723f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A2_c_397_n N_VGND_c_1009_n 0.00146448f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A2_c_398_n N_VGND_c_1010_n 0.00360182f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A2_c_403_n N_VGND_c_1010_n 0.0143482f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_409 N_A2_c_395_n N_VGND_c_1019_n 0.0042294f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A2_c_396_n N_VGND_c_1019_n 0.00421816f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A2_c_397_n N_VGND_c_1021_n 0.00423334f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_412 N_A2_c_398_n N_VGND_c_1021_n 0.00541359f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_413 N_A2_c_395_n N_VGND_c_1024_n 0.00598374f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A2_c_396_n N_VGND_c_1024_n 0.00575258f $X=8.23 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A2_c_397_n N_VGND_c_1024_n 0.0057163f $X=8.65 $Y=0.995 $X2=0 $Y2=0
cc_416 N_A2_c_398_n N_VGND_c_1024_n 0.0105526f $X=9.07 $Y=0.995 $X2=0 $Y2=0
cc_417 N_A2_c_395_n N_A_1241_47#_c_1179_n 0.00306567f $X=6.13 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A2_c_396_n N_A_1241_47#_c_1180_n 0.00255288f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_A2_c_396_n N_A_1241_47#_c_1177_n 0.00485712f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_420 N_A2_c_397_n N_A_1241_47#_c_1177_n 4.58193e-19 $X=8.65 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_A2_c_411_n N_A_1241_47#_c_1177_n 0.00600976f $X=8.095 $Y=1.53 $X2=0
+ $Y2=0
cc_422 N_A2_c_402_n N_A_1241_47#_c_1177_n 0.00799416f $X=8.265 $Y=1.175 $X2=0
+ $Y2=0
cc_423 N_A2_c_396_n N_A_1241_47#_c_1178_n 0.00870038f $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_424 N_A2_c_397_n N_A_1241_47#_c_1178_n 0.00978972f $X=8.65 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_A2_c_398_n N_A_1241_47#_c_1178_n 0.00262807f $X=9.07 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_A2_c_402_n N_A_1241_47#_c_1178_n 0.00596758f $X=8.265 $Y=1.175 $X2=0
+ $Y2=0
cc_427 N_A2_c_403_n N_A_1241_47#_c_1178_n 0.0571359f $X=9 $Y=1.16 $X2=0 $Y2=0
cc_428 N_A2_c_404_n N_A_1241_47#_c_1178_n 0.00452472f $X=9.07 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_A2_c_396_n N_A_1241_47#_c_1191_n 5.22228e-19 $X=8.23 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A2_c_397_n N_A_1241_47#_c_1191_n 0.00630972f $X=8.65 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A2_c_398_n N_A_1241_47#_c_1191_n 0.00539651f $X=9.07 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A1_c_521_n N_Y_c_734_n 0.0086237f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A1_c_522_n N_Y_c_734_n 0.00898061f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A1_c_523_n N_Y_c_734_n 0.00898061f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A1_c_524_n N_Y_c_734_n 0.00269582f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_436 N_A1_c_539_n N_Y_c_734_n 0.0569781f $X=6.64 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A1_c_525_n N_Y_c_734_n 0.00628291f $X=7.81 $Y=1.16 $X2=0 $Y2=0
cc_438 N_A1_c_521_n N_Y_c_666_n 8.89068e-19 $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_439 N_A1_M1003_g N_A_471_297#_c_829_n 0.0106608f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_440 N_A1_M1032_g N_A_471_297#_c_829_n 0.0107426f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_441 N_A1_M1035_g N_A_471_297#_c_829_n 0.0107426f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_442 N_A1_M1039_g N_A_471_297#_c_829_n 0.0106608f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_443 N_A1_M1003_g N_VPWR_c_902_n 0.0165646f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_444 N_A1_M1032_g N_VPWR_c_902_n 0.0165986f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_445 N_A1_M1035_g N_VPWR_c_902_n 0.0165986f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_446 N_A1_M1039_g N_VPWR_c_902_n 0.0165646f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_447 N_A1_c_521_n N_VGND_c_1019_n 0.00357877f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A1_c_522_n N_VGND_c_1019_n 0.00357877f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_449 N_A1_c_523_n N_VGND_c_1019_n 0.00357877f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_450 N_A1_c_524_n N_VGND_c_1019_n 0.00357877f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_451 N_A1_c_521_n N_VGND_c_1024_n 0.00525237f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A1_c_522_n N_VGND_c_1024_n 0.00522516f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_453 N_A1_c_523_n N_VGND_c_1024_n 0.00522516f $X=7.39 $Y=0.995 $X2=0 $Y2=0
cc_454 N_A1_c_524_n N_VGND_c_1024_n 0.00525237f $X=7.81 $Y=0.995 $X2=0 $Y2=0
cc_455 N_A1_c_521_n N_A_1241_47#_c_1179_n 0.00892725f $X=6.55 $Y=0.995 $X2=0
+ $Y2=0
cc_456 N_A1_c_522_n N_A_1241_47#_c_1179_n 0.00892725f $X=6.97 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_A1_c_523_n N_A_1241_47#_c_1179_n 0.00892725f $X=7.39 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A1_c_524_n N_A_1241_47#_c_1179_n 0.0105641f $X=7.81 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A1_c_539_n N_A_1241_47#_c_1179_n 0.00294252f $X=6.64 $Y=1.16 $X2=0
+ $Y2=0
cc_460 N_A1_c_524_n N_A_1241_47#_c_1177_n 6.06509e-19 $X=7.81 $Y=0.995 $X2=0
+ $Y2=0
cc_461 N_A_27_297#_c_588_n N_Y_M1011_d 0.00312348f $X=0.995 $Y=2.38 $X2=0 $Y2=0
cc_462 N_A_27_297#_c_590_n N_Y_M1033_d 0.00312348f $X=1.875 $Y=2.38 $X2=0 $Y2=0
cc_463 N_A_27_297#_c_588_n N_Y_c_750_n 0.0118865f $X=0.995 $Y=2.38 $X2=0 $Y2=0
cc_464 N_A_27_297#_M1030_s N_Y_c_667_n 0.00165831f $X=0.985 $Y=1.485 $X2=0 $Y2=0
cc_465 N_A_27_297#_c_619_p N_Y_c_667_n 0.0126919f $X=1.12 $Y=1.96 $X2=0 $Y2=0
cc_466 N_A_27_297#_c_580_n N_Y_c_668_n 0.00343604f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_467 N_A_27_297#_c_590_n N_Y_c_754_n 0.0118865f $X=1.875 $Y=2.38 $X2=0 $Y2=0
cc_468 N_A_27_297#_c_583_n N_Y_c_661_n 0.0667933f $X=2.735 $Y=1.53 $X2=0 $Y2=0
cc_469 N_A_27_297#_c_584_n N_Y_c_661_n 0.0211595f $X=2.125 $Y=1.53 $X2=0 $Y2=0
cc_470 N_A_27_297#_c_605_n N_Y_c_661_n 0.00518729f $X=5.42 $Y=1.96 $X2=0 $Y2=0
cc_471 N_A_27_297#_c_584_n N_Y_c_670_n 0.00902116f $X=2.125 $Y=1.53 $X2=0 $Y2=0
cc_472 N_A_27_297#_c_583_n N_A_471_297#_M1002_d 0.00278154f $X=2.735 $Y=1.53
+ $X2=-0.19 $Y2=1.305
cc_473 N_A_27_297#_c_605_n N_A_471_297#_M1007_d 0.00552169f $X=5.42 $Y=1.96
+ $X2=0 $Y2=0
cc_474 N_A_27_297#_c_605_n N_A_471_297#_M1008_s 0.00336868f $X=5.42 $Y=1.96
+ $X2=0 $Y2=0
cc_475 N_A_27_297#_c_605_n N_A_471_297#_M1034_s 0.00336868f $X=5.42 $Y=1.96
+ $X2=0 $Y2=0
cc_476 N_A_27_297#_c_581_n N_A_471_297#_c_808_n 0.0147157f $X=2 $Y=2.295 $X2=0
+ $Y2=0
cc_477 N_A_27_297#_c_582_n N_A_471_297#_c_808_n 0.00637684f $X=1.96 $Y=1.63
+ $X2=0 $Y2=0
cc_478 N_A_27_297#_c_582_n N_A_471_297#_c_809_n 0.0309727f $X=1.96 $Y=1.63 $X2=0
+ $Y2=0
cc_479 N_A_27_297#_c_583_n N_A_471_297#_c_809_n 0.0189646f $X=2.735 $Y=1.53
+ $X2=0 $Y2=0
cc_480 N_A_27_297#_M1002_s N_A_471_297#_c_815_n 0.00316082f $X=2.765 $Y=1.485
+ $X2=0 $Y2=0
cc_481 N_A_27_297#_M1023_s N_A_471_297#_c_815_n 0.00316492f $X=3.605 $Y=1.485
+ $X2=0 $Y2=0
cc_482 N_A_27_297#_M1013_d N_A_471_297#_c_815_n 0.00316492f $X=4.445 $Y=1.485
+ $X2=0 $Y2=0
cc_483 N_A_27_297#_M1038_d N_A_471_297#_c_815_n 0.00316492f $X=5.285 $Y=1.485
+ $X2=0 $Y2=0
cc_484 N_A_27_297#_c_583_n N_A_471_297#_c_815_n 0.00292909f $X=2.735 $Y=1.53
+ $X2=0 $Y2=0
cc_485 N_A_27_297#_c_603_n N_A_471_297#_c_815_n 0.0144726f $X=2.882 $Y=1.835
+ $X2=0 $Y2=0
cc_486 N_A_27_297#_c_605_n N_A_471_297#_c_815_n 0.130637f $X=5.42 $Y=1.96 $X2=0
+ $Y2=0
cc_487 N_A_27_297#_M1011_s N_VPWR_c_898_n 0.00225716f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_488 N_A_27_297#_M1030_s N_VPWR_c_898_n 0.00215203f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_489 N_A_27_297#_M1037_s N_VPWR_c_898_n 0.00209324f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_490 N_A_27_297#_M1002_s N_VPWR_c_898_n 0.00216833f $X=2.765 $Y=1.485 $X2=0
+ $Y2=0
cc_491 N_A_27_297#_M1023_s N_VPWR_c_898_n 0.00216833f $X=3.605 $Y=1.485 $X2=0
+ $Y2=0
cc_492 N_A_27_297#_M1013_d N_VPWR_c_898_n 0.00216833f $X=4.445 $Y=1.485 $X2=0
+ $Y2=0
cc_493 N_A_27_297#_M1038_d N_VPWR_c_898_n 0.00216833f $X=5.285 $Y=1.485 $X2=0
+ $Y2=0
cc_494 N_A_27_297#_c_579_n N_VPWR_c_898_n 0.012126f $X=0.247 $Y=2.295 $X2=0
+ $Y2=0
cc_495 N_A_27_297#_c_588_n N_VPWR_c_898_n 0.0204627f $X=0.995 $Y=2.38 $X2=0
+ $Y2=0
cc_496 N_A_27_297#_c_590_n N_VPWR_c_898_n 0.0219525f $X=1.875 $Y=2.38 $X2=0
+ $Y2=0
cc_497 N_A_27_297#_c_581_n N_VPWR_c_898_n 0.00962271f $X=2 $Y=2.295 $X2=0 $Y2=0
cc_498 N_A_27_297#_c_652_p N_VPWR_c_898_n 0.00962794f $X=1.12 $Y=2.38 $X2=0
+ $Y2=0
cc_499 N_A_27_297#_c_579_n N_VPWR_c_906_n 0.0205754f $X=0.247 $Y=2.295 $X2=0
+ $Y2=0
cc_500 N_A_27_297#_c_588_n N_VPWR_c_906_n 0.0330174f $X=0.995 $Y=2.38 $X2=0
+ $Y2=0
cc_501 N_A_27_297#_c_590_n N_VPWR_c_906_n 0.0344282f $X=1.875 $Y=2.38 $X2=0
+ $Y2=0
cc_502 N_A_27_297#_c_581_n N_VPWR_c_906_n 0.0173913f $X=2 $Y=2.295 $X2=0 $Y2=0
cc_503 N_A_27_297#_c_652_p N_VPWR_c_906_n 0.0143053f $X=1.12 $Y=2.38 $X2=0 $Y2=0
cc_504 N_Y_M1011_d N_VPWR_c_898_n 0.00216833f $X=0.565 $Y=1.485 $X2=0 $Y2=0
cc_505 N_Y_M1033_d N_VPWR_c_898_n 0.00216833f $X=1.405 $Y=1.485 $X2=0 $Y2=0
cc_506 N_Y_c_658_n N_VGND_M1019_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_507 N_Y_c_665_n N_VGND_M1025_s 0.00313716f $X=6.29 $Y=0.775 $X2=0 $Y2=0
cc_508 N_Y_c_659_n N_VGND_c_1004_n 0.00752165f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_509 N_Y_c_658_n N_VGND_c_1005_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_510 N_Y_c_660_n N_VGND_c_1007_n 0.00159575f $X=1.605 $Y=1.095 $X2=0 $Y2=0
cc_511 N_Y_c_661_n N_VGND_c_1007_n 0.0144144f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_512 N_Y_c_663_n N_VGND_c_1007_n 0.00850809f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_513 N_Y_c_665_n N_VGND_c_1008_n 0.012101f $X=6.29 $Y=0.775 $X2=0 $Y2=0
cc_514 N_Y_c_671_n N_VGND_c_1011_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_515 N_Y_c_658_n N_VGND_c_1011_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_516 N_Y_c_658_n N_VGND_c_1013_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_517 N_Y_c_689_n N_VGND_c_1013_n 0.0188877f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_518 N_Y_c_662_n N_VGND_c_1015_n 0.00527882f $X=3.16 $Y=1.095 $X2=0 $Y2=0
cc_519 N_Y_c_661_n N_VGND_c_1016_n 0.0634759f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_520 N_Y_c_664_n N_VGND_c_1017_n 0.00156038f $X=5.68 $Y=0.775 $X2=0 $Y2=0
cc_521 N_Y_c_665_n N_VGND_c_1017_n 0.00178152f $X=6.29 $Y=0.775 $X2=0 $Y2=0
cc_522 N_Y_c_665_n N_VGND_c_1019_n 0.00194318f $X=6.29 $Y=0.775 $X2=0 $Y2=0
cc_523 N_Y_M1014_d N_VGND_c_1024_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_524 N_Y_M1027_d N_VGND_c_1024_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_525 N_Y_M1004_d N_VGND_c_1024_n 0.00216833f $X=4.025 $Y=0.235 $X2=0 $Y2=0
cc_526 N_Y_M1017_d N_VGND_c_1024_n 0.00216833f $X=4.865 $Y=0.235 $X2=0 $Y2=0
cc_527 N_Y_M1001_d N_VGND_c_1024_n 0.00216833f $X=6.625 $Y=0.235 $X2=0 $Y2=0
cc_528 N_Y_M1010_d N_VGND_c_1024_n 0.00216833f $X=7.465 $Y=0.235 $X2=0 $Y2=0
cc_529 N_Y_c_671_n N_VGND_c_1024_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_530 N_Y_c_658_n N_VGND_c_1024_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_531 N_Y_c_689_n N_VGND_c_1024_n 0.0122159f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_532 N_Y_c_716_n N_VGND_c_1024_n 0.00650641f $X=5.51 $Y=0.775 $X2=0 $Y2=0
cc_533 N_Y_c_665_n N_VGND_c_1024_n 0.00870024f $X=6.29 $Y=0.775 $X2=0 $Y2=0
cc_534 N_Y_c_662_n N_A_453_47#_M1012_d 0.00109912f $X=3.16 $Y=1.095 $X2=0 $Y2=0
cc_535 N_Y_c_714_n N_A_453_47#_M1012_d 8.85226e-19 $X=3.245 $Y=0.732 $X2=0 $Y2=0
cc_536 N_Y_c_716_n N_A_453_47#_M1012_d 0.0160298f $X=5.51 $Y=0.775 $X2=0 $Y2=0
cc_537 N_Y_c_716_n N_A_453_47#_M1015_s 0.00307941f $X=5.51 $Y=0.775 $X2=0 $Y2=0
cc_538 N_Y_c_716_n N_A_453_47#_M1020_s 0.00447855f $X=5.51 $Y=0.775 $X2=0 $Y2=0
cc_539 N_Y_c_661_n N_A_453_47#_c_1141_n 9.37998e-19 $X=3.075 $Y=1.185 $X2=0
+ $Y2=0
cc_540 N_Y_c_714_n N_A_453_47#_c_1141_n 0.00862495f $X=3.245 $Y=0.732 $X2=0
+ $Y2=0
cc_541 N_Y_c_716_n N_A_453_47#_c_1141_n 0.062885f $X=5.51 $Y=0.775 $X2=0 $Y2=0
cc_542 N_Y_M1004_d N_A_453_47#_c_1143_n 0.00305026f $X=4.025 $Y=0.235 $X2=0
+ $Y2=0
cc_543 N_Y_M1017_d N_A_453_47#_c_1143_n 0.00305026f $X=4.865 $Y=0.235 $X2=0
+ $Y2=0
cc_544 N_Y_c_664_n N_A_453_47#_c_1143_n 0.062885f $X=5.68 $Y=0.775 $X2=0 $Y2=0
cc_545 N_Y_c_661_n N_A_453_47#_c_1146_n 0.0022631f $X=3.075 $Y=1.185 $X2=0 $Y2=0
cc_546 N_Y_c_665_n N_A_1241_47#_M1005_d 3.3779e-19 $X=6.29 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_547 N_Y_c_666_n N_A_1241_47#_M1005_d 0.00249059f $X=6.46 $Y=0.775 $X2=-0.19
+ $Y2=-0.24
cc_548 N_Y_c_734_n N_A_1241_47#_M1006_s 0.0033322f $X=7.6 $Y=0.73 $X2=0 $Y2=0
cc_549 N_Y_M1001_d N_A_1241_47#_c_1179_n 0.00305026f $X=6.625 $Y=0.235 $X2=0
+ $Y2=0
cc_550 N_Y_M1010_d N_A_1241_47#_c_1179_n 0.00305026f $X=7.465 $Y=0.235 $X2=0
+ $Y2=0
cc_551 N_Y_c_665_n N_A_1241_47#_c_1179_n 0.00268596f $X=6.29 $Y=0.775 $X2=0
+ $Y2=0
cc_552 N_Y_c_666_n N_A_1241_47#_c_1179_n 0.0737736f $X=6.46 $Y=0.775 $X2=0 $Y2=0
cc_553 N_A_471_297#_c_829_n N_VPWR_M1016_d 0.00328256f $X=8.355 $Y=1.915
+ $X2=-0.19 $Y2=1.305
cc_554 N_A_471_297#_c_829_n N_VPWR_M1032_s 0.00319635f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_555 N_A_471_297#_c_829_n N_VPWR_M1039_s 0.00328335f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_556 N_A_471_297#_c_810_n N_VPWR_M1031_d 0.00169858f $X=9.155 $Y=1.53 $X2=0
+ $Y2=0
cc_557 N_A_471_297#_c_810_n N_VPWR_c_899_n 0.0121607f $X=9.155 $Y=1.53 $X2=0
+ $Y2=0
cc_558 N_A_471_297#_c_829_n N_VPWR_c_900_n 0.0022675f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_559 N_A_471_297#_c_874_p N_VPWR_c_900_n 0.0113958f $X=8.44 $Y=2.3 $X2=0 $Y2=0
cc_560 N_A_471_297#_c_846_n N_VPWR_c_900_n 9.22958e-19 $X=8.44 $Y=1.96 $X2=0
+ $Y2=0
cc_561 N_A_471_297#_M1003_d N_VPWR_c_902_n 0.00172715f $X=6.625 $Y=1.485 $X2=0
+ $Y2=0
cc_562 N_A_471_297#_M1035_d N_VPWR_c_902_n 0.00172715f $X=7.465 $Y=1.485 $X2=0
+ $Y2=0
cc_563 N_A_471_297#_c_829_n N_VPWR_c_903_n 0.110047f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_564 N_A_471_297#_c_879_p N_VPWR_c_904_n 0.0158369f $X=9.28 $Y=1.62 $X2=0
+ $Y2=0
cc_565 N_A_471_297#_M1002_d N_VPWR_c_898_n 0.00209324f $X=2.355 $Y=1.485 $X2=0
+ $Y2=0
cc_566 N_A_471_297#_M1007_d N_VPWR_c_898_n 0.00215227f $X=3.185 $Y=1.485 $X2=0
+ $Y2=0
cc_567 N_A_471_297#_M1008_s N_VPWR_c_898_n 0.00215227f $X=4.025 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_A_471_297#_M1034_s N_VPWR_c_898_n 0.00215227f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_569 N_A_471_297#_M1026_d N_VPWR_c_898_n 0.00300176f $X=5.705 $Y=1.485 $X2=0
+ $Y2=0
cc_570 N_A_471_297#_M1024_s N_VPWR_c_898_n 0.00254985f $X=8.305 $Y=1.485 $X2=0
+ $Y2=0
cc_571 N_A_471_297#_M1036_s N_VPWR_c_898_n 0.00397704f $X=9.145 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_471_297#_c_808_n N_VPWR_c_898_n 0.00962421f $X=2.44 $Y=2.215 $X2=0
+ $Y2=0
cc_573 N_A_471_297#_c_815_n N_VPWR_c_898_n 0.113773f $X=5.755 $Y=2.34 $X2=0
+ $Y2=0
cc_574 N_A_471_297#_c_889_p N_VPWR_c_898_n 0.00962271f $X=5.88 $Y=2.215 $X2=0
+ $Y2=0
cc_575 N_A_471_297#_c_829_n N_VPWR_c_898_n 0.0165668f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_576 N_A_471_297#_c_874_p N_VPWR_c_898_n 0.00646998f $X=8.44 $Y=2.3 $X2=0
+ $Y2=0
cc_577 N_A_471_297#_c_879_p N_VPWR_c_898_n 0.00955092f $X=9.28 $Y=1.62 $X2=0
+ $Y2=0
cc_578 N_A_471_297#_c_846_n N_VPWR_c_898_n 0.00211648f $X=8.44 $Y=1.96 $X2=0
+ $Y2=0
cc_579 N_A_471_297#_c_808_n N_VPWR_c_906_n 0.0173726f $X=2.44 $Y=2.215 $X2=0
+ $Y2=0
cc_580 N_A_471_297#_c_815_n N_VPWR_c_906_n 0.178242f $X=5.755 $Y=2.34 $X2=0
+ $Y2=0
cc_581 N_A_471_297#_c_889_p N_VPWR_c_906_n 0.0170924f $X=5.88 $Y=2.215 $X2=0
+ $Y2=0
cc_582 N_A_471_297#_c_829_n N_VPWR_c_906_n 0.0022675f $X=8.355 $Y=1.915 $X2=0
+ $Y2=0
cc_583 N_VGND_c_1016_n N_A_453_47#_M1000_d 0.00162688f $X=2.735 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_584 N_VGND_c_1024_n N_A_453_47#_M1000_d 0.00215227f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_585 N_VGND_c_1024_n N_A_453_47#_M1012_d 0.00623662f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_1024_n N_A_453_47#_M1015_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_1024_n N_A_453_47#_M1020_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1008_n N_A_453_47#_c_1143_n 0.0127119f $X=5.92 $Y=0.39 $X2=0
+ $Y2=0
cc_589 N_VGND_c_1006_n N_A_453_47#_c_1144_n 0.0155499f $X=1.96 $Y=0.39 $X2=0
+ $Y2=0
cc_590 N_VGND_c_1016_n N_A_453_47#_c_1144_n 0.0184859f $X=2.735 $Y=0.76 $X2=0
+ $Y2=0
cc_591 N_VGND_c_1017_n N_A_453_47#_c_1144_n 0.190267f $X=5.835 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_1024_n N_A_453_47#_c_1144_n 0.120434f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_M1009_s N_A_453_47#_c_1146_n 0.00303853f $X=2.685 $Y=0.235 $X2=0
+ $Y2=0
cc_594 N_VGND_c_1015_n N_A_453_47#_c_1146_n 0.0111953f $X=2.82 $Y=0.76 $X2=0
+ $Y2=0
cc_595 N_VGND_c_1016_n N_A_453_47#_c_1146_n 0.00387778f $X=2.735 $Y=0.76 $X2=0
+ $Y2=0
cc_596 N_VGND_c_1024_n N_A_1241_47#_M1005_d 0.00215227f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_597 N_VGND_c_1024_n N_A_1241_47#_M1006_s 0.00215227f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_1024_n N_A_1241_47#_M1021_s 0.00215206f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_c_1024_n N_A_1241_47#_M1022_d 0.00215201f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_600 N_VGND_c_1019_n N_A_1241_47#_c_1179_n 0.0973818f $X=8.355 $Y=0 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1024_n N_A_1241_47#_c_1179_n 0.0626919f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1019_n N_A_1241_47#_c_1180_n 0.0152108f $X=8.355 $Y=0 $X2=0
+ $Y2=0
cc_603 N_VGND_c_1024_n N_A_1241_47#_c_1180_n 0.00940698f $X=9.43 $Y=0 $X2=0
+ $Y2=0
cc_604 N_VGND_M1018_s N_A_1241_47#_c_1178_n 0.00162089f $X=8.305 $Y=0.235 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1009_n N_A_1241_47#_c_1178_n 0.0122559f $X=8.44 $Y=0.39 $X2=0
+ $Y2=0
cc_606 N_VGND_c_1010_n N_A_1241_47#_c_1178_n 0.00830019f $X=9.28 $Y=0.39 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1019_n N_A_1241_47#_c_1178_n 0.00198695f $X=8.355 $Y=0 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1021_n N_A_1241_47#_c_1178_n 0.00198695f $X=9.195 $Y=0 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1024_n N_A_1241_47#_c_1178_n 0.00835832f $X=9.43 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1021_n N_A_1241_47#_c_1191_n 0.0188551f $X=9.195 $Y=0 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1024_n N_A_1241_47#_c_1191_n 0.0122069f $X=9.43 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nor2b_2.pex.spice
* Created: Tue Sep  1 19:18:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR2B_2%A 1 3 6 8 10 13 15 22
r37 20 22 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.645 $Y=1.16
+ $X2=0.91 $Y2=1.16
r38 17 20 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.645 $Y2=1.16
r39 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r40 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r41 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r42 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r43 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r44 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r45 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r46 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r47 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%A_251_21# 1 2 7 9 12 14 16 19 21 25 28 31 33
+ 34 39 43 45 48
c84 31 0 2.92742e-20 $X=2.322 $Y=1.075
r85 46 48 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.345 $Y=1.53
+ $X2=2.48 $Y2=1.53
r86 37 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=1.615
+ $X2=2.48 $Y2=1.53
r87 37 39 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.48 $Y=1.615
+ $X2=2.48 $Y2=2.28
r88 34 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.725
+ $X2=2.48 $Y2=0.81
r89 34 36 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=2.48 $Y=0.725
+ $X2=2.48 $Y2=0.68
r90 33 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=1.445
+ $X2=2.345 $Y2=1.53
r91 32 45 4.65272 $w=1.92e-07 $l=9.58123e-08 $layer=LI1_cond $X=2.345 $Y=1.245
+ $X2=2.322 $Y2=1.16
r92 32 33 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.345 $Y=1.245
+ $X2=2.345 $Y2=1.445
r93 31 45 4.65272 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=2.322 $Y=1.075
+ $X2=2.322 $Y2=1.16
r94 30 43 10.308 $w=1.68e-07 $l=1.58e-07 $layer=LI1_cond $X=2.322 $Y=0.81
+ $X2=2.48 $Y2=0.81
r95 30 31 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=2.322 $Y=0.895
+ $X2=2.322 $Y2=1.075
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.16 $X2=2.04 $Y2=1.16
r97 25 45 1.79375 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.215 $Y=1.16
+ $X2=2.322 $Y2=1.16
r98 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.215 $Y=1.16
+ $X2=2.04 $Y2=1.16
r99 22 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.33 $Y=1.16
+ $X2=1.75 $Y2=1.16
r100 21 28 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.825 $Y=1.16
+ $X2=2.04 $Y2=1.16
r101 21 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.825 $Y=1.16
+ $X2=1.75 $Y2=1.16
r102 17 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r103 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r104 14 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r105 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r106 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r107 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r108 7 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r109 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r110 2 39 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=2.065 $X2=2.48 $Y2=2.28
r111 1 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.465 $X2=2.48 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%B_N 3 6 8 9 10 17 19
c35 17 0 2.92742e-20 $X=2.765 $Y=1.16
r36 17 20 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=2.757 $Y=1.16
+ $X2=2.757 $Y2=1.325
r37 17 19 48.1214 $w=2.85e-07 $l=1.65e-07 $layer=POLY_cond $X=2.757 $Y=1.16
+ $X2=2.757 $Y2=0.995
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.16 $X2=2.765 $Y2=1.16
r39 9 10 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=3.017 $Y=1.53
+ $X2=3.017 $Y2=1.87
r40 8 18 6.68646 $w=3.78e-07 $l=1.45e-07 $layer=LI1_cond $X=2.91 $Y=1.17
+ $X2=2.765 $Y2=1.17
r41 8 9 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.017 $Y=1.275
+ $X2=3.017 $Y2=1.53
r42 6 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.69 $Y=2.275
+ $X2=2.69 $Y2=1.325
r43 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.69 $Y=0.675
+ $X2=2.69 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%A_27_297# 1 2 3 10 12 14 16 17 18 22 24 25
r44 25 34 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.295
+ $X2=1.98 $Y2=2.38
r45 24 32 5.95937 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.98 $Y=2.035
+ $X2=1.98 $Y2=1.89
r46 24 25 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=1.98 $Y=2.035
+ $X2=1.98 $Y2=2.295
r47 22 32 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=1.962 $Y=1.63
+ $X2=1.962 $Y2=1.89
r48 19 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.38
+ $X2=1.12 $Y2=2.38
r49 18 34 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.835 $Y=2.38
+ $X2=1.98 $Y2=2.38
r50 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.835 $Y=2.38
+ $X2=1.245 $Y2=2.38
r51 17 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.295
+ $X2=1.12 $Y2=2.38
r52 16 29 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.12 $Y=1.655
+ $X2=1.12 $Y2=1.55
r53 16 17 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=1.12 $Y=1.655
+ $X2=1.12 $Y2=2.295
r54 15 27 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=0.405 $Y=1.55
+ $X2=0.245 $Y2=1.55
r55 14 29 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=1.55
+ $X2=1.12 $Y2=1.55
r56 14 15 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=0.995 $Y=1.55
+ $X2=0.405 $Y2=1.55
r57 10 27 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=1.55
r58 10 12 23.2289 $w=3.18e-07 $l=6.45e-07 $layer=LI1_cond $X=0.245 $Y=1.655
+ $X2=0.245 $Y2=2.3
r59 3 34 400 $w=1.7e-07 $l=8.89944e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=2.31
r60 3 22 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.485 $X2=1.96 $Y2=1.63
r61 2 31 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=2.3
r62 2 29 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r63 1 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r64 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%VPWR 1 2 9 11 13 15 17 22 31 35
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 23 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=0.7 $Y2=2.72
r50 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.825 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 22 34 3.9252 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.997 $Y2=2.72
r52 22 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.53 $Y2=2.72
r53 17 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.7 $Y2=2.72
r54 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.575 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 11 34 3.21796 $w=2.5e-07 $l=1.32868e-07 $layer=LI1_cond $X=2.9 $Y=2.635
+ $X2=2.997 $Y2=2.72
r58 11 13 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=2.9 $Y=2.635
+ $X2=2.9 $Y2=2.31
r59 7 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.72
r60 7 9 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2
r61 2 13 600 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=2.065 $X2=2.9 $Y2=2.31
r62 1 9 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%Y 1 2 3 12 14 15 18 21 22 25
r50 22 25 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.54 $Y=0.51 $X2=1.54
+ $Y2=0.39
r51 20 22 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.51
r52 20 21 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.725
+ $X2=1.54 $Y2=0.81
r53 16 21 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=0.895
+ $X2=1.54 $Y2=0.81
r54 16 18 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=1.54 $Y=0.895
+ $X2=1.54 $Y2=1.62
r55 14 21 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.81
+ $X2=1.54 $Y2=0.81
r56 14 15 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.375 $Y=0.81
+ $X2=0.865 $Y2=0.81
r57 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.7 $Y=0.725
+ $X2=0.865 $Y2=0.81
r58 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=0.725 $X2=0.7
+ $Y2=0.39
r59 3 18 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r60 2 25 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.39
r61 1 12 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR2B_2%VGND 1 2 3 4 13 15 19 23 25 27 30 31 33 34
+ 35 44 53
r53 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r54 47 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r56 44 52 3.96354 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.997
+ $Y2=0
r57 44 46 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.53
+ $Y2=0
r58 43 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r59 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r60 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r61 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r62 37 49 4.33083 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r63 37 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r64 35 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 35 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 33 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.61
+ $Y2=0
r67 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.96
+ $Y2=0
r68 32 46 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.045 $Y=0 $X2=2.53
+ $Y2=0
r69 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0 $X2=1.96
+ $Y2=0
r70 30 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r71 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.12
+ $Y2=0
r72 29 42 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.61
+ $Y2=0
r73 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.12
+ $Y2=0
r74 25 52 3.21368 $w=2.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.902 $Y=0.085
+ $X2=2.997 $Y2=0
r75 25 27 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=2.902 $Y=0.085
+ $X2=2.902 $Y2=0.68
r76 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r77 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.39
r78 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r79 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r80 13 49 3.02922 $w=2.8e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.182 $Y2=0
r81 13 15 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.39
r82 4 27 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.465 $X2=2.9 $Y2=0.68
r83 3 23 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r84 2 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r85 1 15 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__o2bb2ai_4.pxi.spice
* Created: Tue Sep  1 19:24:14 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A2_N N_A2_N_c_156_n N_A2_N_M1008_g
+ N_A2_N_M1005_g N_A2_N_c_157_n N_A2_N_M1012_g N_A2_N_M1021_g N_A2_N_c_158_n
+ N_A2_N_M1017_g N_A2_N_M1025_g N_A2_N_c_159_n N_A2_N_M1019_g N_A2_N_M1034_g
+ A2_N N_A2_N_c_160_n N_A2_N_c_161_n PM_SKY130_FD_SC_HD__O2BB2AI_4%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A1_N N_A1_N_c_218_n N_A1_N_M1014_g
+ N_A1_N_M1004_g N_A1_N_c_219_n N_A1_N_M1020_g N_A1_N_M1015_g N_A1_N_c_220_n
+ N_A1_N_M1023_g N_A1_N_M1016_g N_A1_N_c_221_n N_A1_N_M1027_g N_A1_N_M1026_g
+ A1_N N_A1_N_c_222_n N_A1_N_c_223_n PM_SKY130_FD_SC_HD__O2BB2AI_4%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A_113_47# N_A_113_47#_M1008_d
+ N_A_113_47#_M1017_d N_A_113_47#_M1005_d N_A_113_47#_M1025_d
+ N_A_113_47#_M1004_s N_A_113_47#_M1016_s N_A_113_47#_M1001_g
+ N_A_113_47#_c_296_n N_A_113_47#_M1007_g N_A_113_47#_M1006_g
+ N_A_113_47#_c_297_n N_A_113_47#_M1009_g N_A_113_47#_M1022_g
+ N_A_113_47#_c_298_n N_A_113_47#_M1011_g N_A_113_47#_M1028_g
+ N_A_113_47#_c_299_n N_A_113_47#_M1013_g N_A_113_47#_c_300_n
+ N_A_113_47#_c_301_n N_A_113_47#_c_302_n N_A_113_47#_c_312_n
+ N_A_113_47#_c_313_n N_A_113_47#_c_382_p N_A_113_47#_c_314_n
+ N_A_113_47#_c_378_p N_A_113_47#_c_315_n N_A_113_47#_c_379_p
+ N_A_113_47#_c_316_n N_A_113_47#_c_383_p N_A_113_47#_c_317_n
+ N_A_113_47#_c_303_n N_A_113_47#_c_304_n N_A_113_47#_c_305_n
+ N_A_113_47#_c_319_n N_A_113_47#_c_320_n N_A_113_47#_c_321_n
+ N_A_113_47#_c_322_n N_A_113_47#_c_306_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%A_113_47#
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%B2 N_B2_c_452_n N_B2_M1024_g N_B2_M1003_g
+ N_B2_c_453_n N_B2_M1031_g N_B2_M1010_g N_B2_c_454_n N_B2_M1032_g N_B2_M1033_g
+ N_B2_c_455_n N_B2_M1038_g N_B2_M1036_g B2 N_B2_c_464_p N_B2_c_456_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%B2
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%B1 N_B1_c_533_n N_B1_M1000_g N_B1_M1018_g
+ N_B1_c_534_n N_B1_M1002_g N_B1_M1029_g N_B1_c_535_n N_B1_M1035_g N_B1_M1030_g
+ N_B1_c_536_n N_B1_M1039_g N_B1_M1037_g B1 N_B1_c_537_n N_B1_c_538_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%B1
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%VPWR N_VPWR_M1005_s N_VPWR_M1021_s
+ N_VPWR_M1034_s N_VPWR_M1015_d N_VPWR_M1026_d N_VPWR_M1006_d N_VPWR_M1028_d
+ N_VPWR_M1018_s N_VPWR_M1030_s N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n
+ N_VPWR_c_612_n N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n
+ N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n N_VPWR_c_621_n
+ N_VPWR_c_622_n N_VPWR_c_623_n N_VPWR_c_624_n N_VPWR_c_625_n N_VPWR_c_626_n
+ N_VPWR_c_627_n N_VPWR_c_628_n N_VPWR_c_629_n VPWR N_VPWR_c_630_n
+ N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_608_n N_VPWR_c_634_n N_VPWR_c_635_n
+ N_VPWR_c_636_n VPWR PM_SKY130_FD_SC_HD__O2BB2AI_4%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%Y N_Y_M1007_s N_Y_M1011_s N_Y_M1001_s
+ N_Y_M1022_s N_Y_M1003_s N_Y_M1033_s N_Y_c_758_n N_Y_c_760_n N_Y_c_811_n
+ N_Y_c_761_n N_Y_c_815_n N_Y_c_762_n N_Y_c_759_n N_Y_c_764_n N_Y_c_765_n
+ N_Y_c_766_n N_Y_c_767_n N_Y_c_768_n N_Y_c_769_n Y
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%Y
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A_1241_297# N_A_1241_297#_M1003_d
+ N_A_1241_297#_M1010_d N_A_1241_297#_M1036_d N_A_1241_297#_M1029_d
+ N_A_1241_297#_M1037_d N_A_1241_297#_c_844_n N_A_1241_297#_c_852_n
+ N_A_1241_297#_c_845_n N_A_1241_297#_c_901_n N_A_1241_297#_c_854_n
+ N_A_1241_297#_c_846_n N_A_1241_297#_c_882_n N_A_1241_297#_c_847_n
+ N_A_1241_297#_c_886_n N_A_1241_297#_c_848_n N_A_1241_297#_c_849_n
+ N_A_1241_297#_c_850_n N_A_1241_297#_c_892_n N_A_1241_297#_c_851_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%A_1241_297#
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1012_s
+ N_A_27_47#_M1019_s N_A_27_47#_M1020_d N_A_27_47#_M1027_d N_A_27_47#_c_907_n
+ N_A_27_47#_c_918_n N_A_27_47#_c_908_n N_A_27_47#_c_909_n N_A_27_47#_c_926_n
+ N_A_27_47#_c_910_n N_A_27_47#_c_911_n N_A_27_47#_c_912_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%A_27_47#
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%VGND N_VGND_M1014_s N_VGND_M1023_s
+ N_VGND_M1024_d N_VGND_M1032_d N_VGND_M1000_s N_VGND_M1035_s N_VGND_c_980_n
+ N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n N_VGND_c_984_n N_VGND_c_985_n
+ N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n
+ N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n VGND N_VGND_c_994_n
+ N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n N_VGND_c_999_n
+ VGND PM_SKY130_FD_SC_HD__O2BB2AI_4%VGND
x_PM_SKY130_FD_SC_HD__O2BB2AI_4%A_807_47# N_A_807_47#_M1007_d
+ N_A_807_47#_M1009_d N_A_807_47#_M1013_d N_A_807_47#_M1031_s
+ N_A_807_47#_M1038_s N_A_807_47#_M1002_d N_A_807_47#_M1039_d
+ N_A_807_47#_c_1131_n N_A_807_47#_c_1132_n N_A_807_47#_c_1197_n
+ N_A_807_47#_c_1139_n N_A_807_47#_c_1137_n N_A_807_47#_c_1122_n
+ N_A_807_47#_c_1123_n N_A_807_47#_c_1148_n N_A_807_47#_c_1124_n
+ N_A_807_47#_c_1156_n N_A_807_47#_c_1125_n N_A_807_47#_c_1170_n
+ N_A_807_47#_c_1126_n N_A_807_47#_c_1127_n N_A_807_47#_c_1128_n
+ N_A_807_47#_c_1129_n N_A_807_47#_c_1130_n
+ PM_SKY130_FD_SC_HD__O2BB2AI_4%A_807_47#
cc_1 VNB N_A2_N_c_156_n 0.0192294f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A2_N_c_157_n 0.0157856f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A2_N_c_158_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A2_N_c_159_n 0.0161471f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A2_N_c_160_n 0.00156728f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_6 VNB N_A2_N_c_161_n 0.0654289f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_A1_N_c_218_n 0.0159983f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_A1_N_c_219_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_9 VNB N_A1_N_c_220_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_10 VNB N_A1_N_c_221_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_11 VNB N_A1_N_c_222_n 0.00378123f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_12 VNB N_A1_N_c_223_n 0.0683205f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_13 VNB N_A_113_47#_c_296_n 0.0215042f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_14 VNB N_A_113_47#_c_297_n 0.0158044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_113_47#_c_298_n 0.0157858f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.16
cc_16 VNB N_A_113_47#_c_299_n 0.0192404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_113_47#_c_300_n 0.0190401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_113_47#_c_301_n 0.0116419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_113_47#_c_302_n 0.0087143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_113_47#_c_303_n 5.22495e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_113_47#_c_304_n 0.00772394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_113_47#_c_305_n 0.0159479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_113_47#_c_306_n 0.0744578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_B2_c_452_n 0.0194674f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_25 VNB N_B2_c_453_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_26 VNB N_B2_c_454_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_27 VNB N_B2_c_455_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_28 VNB N_B2_c_456_n 0.0676368f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_29 VNB N_B1_c_533_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_30 VNB N_B1_c_534_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_31 VNB N_B1_c_535_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_32 VNB N_B1_c_536_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_33 VNB N_B1_c_537_n 0.029244f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_34 VNB N_B1_c_538_n 0.0689339f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_35 VNB N_VPWR_c_608_n 0.421552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_758_n 0.00917992f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_37 VNB N_Y_c_759_n 0.0110217f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_38 VNB N_A_27_47#_c_907_n 0.00973351f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_39 VNB N_A_27_47#_c_908_n 0.00356055f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_40 VNB N_A_27_47#_c_909_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_41 VNB N_A_27_47#_c_910_n 0.00855566f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_911_n 0.00481776f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_43 VNB N_A_27_47#_c_912_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_44 VNB N_VGND_c_980_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_981_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.325
cc_46 VNB N_VGND_c_982_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.105
cc_47 VNB N_VGND_c_983_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_48 VNB N_VGND_c_984_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.16
cc_49 VNB N_VGND_c_985_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_50 VNB N_VGND_c_986_n 0.0548409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_987_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=1.14 $Y2=1.18
cc_52 VNB N_VGND_c_988_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.18
cc_53 VNB N_VGND_c_989_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_990_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_991_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_992_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_993_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_994_n 0.0788726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_995_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_996_n 0.0226353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_997_n 0.48415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_998_n 0.00323594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_999_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_807_47#_c_1122_n 0.00217448f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_807_47#_c_1123_n 0.00233699f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_66 VNB N_A_807_47#_c_1124_n 0.00217664f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.16
cc_67 VNB N_A_807_47#_c_1125_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_807_47#_c_1126_n 0.0126428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_807_47#_c_1127_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_807_47#_c_1128_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_807_47#_c_1129_n 0.00384439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_807_47#_c_1130_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VPB N_A2_N_M1005_g 0.0220093f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_74 VPB N_A2_N_M1021_g 0.0182022f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_75 VPB N_A2_N_M1025_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_76 VPB N_A2_N_M1034_g 0.0185045f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_77 VPB N_A2_N_c_161_n 0.0102949f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_78 VPB N_A1_N_M1004_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_79 VPB N_A1_N_M1015_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_80 VPB N_A1_N_M1016_g 0.0182034f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_81 VPB N_A1_N_M1026_g 0.0221564f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_82 VPB N_A1_N_c_223_n 0.0103216f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_83 VPB N_A_113_47#_M1001_g 0.0225066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_113_47#_M1006_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_113_47#_M1022_g 0.0182029f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_86 VPB N_A_113_47#_M1028_g 0.0220777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_113_47#_c_300_n 0.00736047f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_113_47#_c_312_n 0.00221293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_113_47#_c_313_n 0.00934466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_113_47#_c_314_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_113_47#_c_315_n 0.00522373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_113_47#_c_316_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_113_47#_c_317_n 0.00426889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_113_47#_c_303_n 0.00409746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_113_47#_c_319_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_113_47#_c_320_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_113_47#_c_321_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_113_47#_c_322_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_113_47#_c_306_n 0.0115076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_B2_M1003_g 0.0223128f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_101 VPB N_B2_M1010_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_102 VPB N_B2_M1033_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_103 VPB N_B2_M1036_g 0.018818f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_104 VPB N_B2_c_456_n 0.0103501f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_105 VPB N_B1_M1018_g 0.0185045f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_106 VPB N_B1_M1029_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_107 VPB N_B1_M1030_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_108 VPB N_B1_M1037_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_109 VPB N_B1_c_538_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_110 VPB N_VPWR_c_609_n 0.011928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_610_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_611_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_113 VPB N_VPWR_c_612_n 0.00393015f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.16
cc_114 VPB N_VPWR_c_613_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_614_n 0.00663054f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_615_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_616_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_617_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_618_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_619_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_620_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_621_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_622_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_623_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_624_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_625_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_626_n 0.056414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_627_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_628_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_629_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_630_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_631_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_632_n 0.0223167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_608_n 0.0626094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_634_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_635_n 0.0142078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_636_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_Y_c_760_n 0.00236072f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.325
cc_139 VPB N_Y_c_761_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.105
cc_140 VPB N_Y_c_762_n 0.00253896f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_141 VPB N_Y_c_759_n 0.00473618f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.16
cc_142 VPB N_Y_c_764_n 0.00935741f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.16
cc_143 VPB N_Y_c_765_n 0.00234634f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.18
cc_144 VPB N_Y_c_766_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_Y_c_767_n 0.0103659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_Y_c_768_n 0.0020229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_Y_c_769_n 0.00224497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_1241_297#_c_844_n 0.00485118f $X=-0.19 $Y=1.305 $X2=1.33
+ $Y2=1.325
cc_149 VPB N_A_1241_297#_c_845_n 0.00179695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_1241_297#_c_846_n 0.00357073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_1241_297#_c_847_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_1241_297#_c_848_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_153 VPB N_A_1241_297#_c_849_n 0.0101972f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.16
cc_154 VPB N_A_1241_297#_c_850_n 0.032524f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=1.16
cc_155 VPB N_A_1241_297#_c_851_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 N_A2_N_c_159_n N_A1_N_c_218_n 0.0193361f $X=1.75 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_157 N_A2_N_M1034_g N_A1_N_M1004_g 0.0193361f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A2_N_c_160_n N_A1_N_c_222_n 0.0121231f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A2_N_c_161_n N_A1_N_c_222_n 2.62535e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A2_N_c_160_n N_A1_N_c_223_n 2.62535e-19 $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A2_N_c_161_n N_A1_N_c_223_n 0.0193361f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_N_c_156_n N_A_113_47#_c_300_n 0.0182079f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A2_N_c_160_n N_A_113_47#_c_300_n 0.0166223f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A2_N_c_156_n N_A_113_47#_c_302_n 0.0133993f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A2_N_c_157_n N_A_113_47#_c_302_n 0.0109625f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A2_N_c_158_n N_A_113_47#_c_302_n 0.0109625f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A2_N_c_159_n N_A_113_47#_c_302_n 0.00372684f $X=1.75 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A2_N_c_160_n N_A_113_47#_c_302_n 0.0943373f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A2_N_c_161_n N_A_113_47#_c_302_n 0.00672641f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_170 N_A2_N_M1005_g N_A_113_47#_c_312_n 0.0149006f $X=0.49 $Y=1.985 $X2=0
+ $Y2=0
cc_171 N_A2_N_c_160_n N_A_113_47#_c_312_n 0.0103349f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A2_N_M1021_g N_A_113_47#_c_314_n 0.0132714f $X=0.91 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A2_N_M1025_g N_A_113_47#_c_314_n 0.0132714f $X=1.33 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A2_N_c_160_n N_A_113_47#_c_314_n 0.0416643f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A2_N_c_161_n N_A_113_47#_c_314_n 0.00211509f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A2_N_M1034_g N_A_113_47#_c_315_n 0.0132273f $X=1.75 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A2_N_c_160_n N_A_113_47#_c_315_n 0.0110239f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A2_N_c_160_n N_A_113_47#_c_319_n 0.0204549f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A2_N_c_161_n N_A_113_47#_c_319_n 0.00220041f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A2_N_c_160_n N_A_113_47#_c_320_n 0.0204549f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A2_N_c_161_n N_A_113_47#_c_320_n 0.00220041f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_182 N_A2_N_M1005_g N_VPWR_c_610_n 0.00338128f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_N_M1021_g N_VPWR_c_611_n 0.00157837f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A2_N_M1025_g N_VPWR_c_611_n 0.00157837f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A2_N_M1034_g N_VPWR_c_612_n 0.00157837f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A2_N_M1025_g N_VPWR_c_620_n 0.00585385f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_N_M1034_g N_VPWR_c_620_n 0.00585385f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_N_M1005_g N_VPWR_c_630_n 0.00585385f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A2_N_M1021_g N_VPWR_c_630_n 0.00585385f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_N_M1005_g N_VPWR_c_608_n 0.0114096f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A2_N_M1021_g N_VPWR_c_608_n 0.0104367f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A2_N_M1025_g N_VPWR_c_608_n 0.0104367f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A2_N_M1034_g N_VPWR_c_608_n 0.010464f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A2_N_c_156_n N_A_27_47#_c_907_n 0.00892725f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_195 N_A2_N_c_157_n N_A_27_47#_c_907_n 0.00892725f $X=0.91 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_158_n N_A_27_47#_c_907_n 0.00892725f $X=1.33 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A2_N_c_159_n N_A_27_47#_c_907_n 0.0105669f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_N_c_160_n N_A_27_47#_c_907_n 0.00295908f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A2_N_c_156_n N_VGND_c_986_n 0.00357877f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_N_c_157_n N_VGND_c_986_n 0.00357877f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A2_N_c_158_n N_VGND_c_986_n 0.00357877f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A2_N_c_159_n N_VGND_c_986_n 0.00357877f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A2_N_c_156_n N_VGND_c_997_n 0.00619805f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A2_N_c_157_n N_VGND_c_997_n 0.00522516f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_N_c_158_n N_VGND_c_997_n 0.00522516f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_206 N_A2_N_c_159_n N_VGND_c_997_n 0.00525237f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A1_N_M1004_g N_A_113_47#_c_315_n 0.0132273f $X=2.17 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A1_N_c_222_n N_A_113_47#_c_315_n 0.0110239f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A1_N_M1015_g N_A_113_47#_c_316_n 0.0132714f $X=2.59 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A1_N_M1016_g N_A_113_47#_c_316_n 0.0132714f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A1_N_c_222_n N_A_113_47#_c_316_n 0.0416643f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A1_N_c_223_n N_A_113_47#_c_316_n 0.00211509f $X=3.43 $Y=1.16 $X2=0
+ $Y2=0
cc_213 N_A1_N_M1026_g N_A_113_47#_c_317_n 0.0149576f $X=3.43 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A1_N_c_222_n N_A_113_47#_c_317_n 0.0110239f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A1_N_c_223_n N_A_113_47#_c_303_n 0.00562056f $X=3.43 $Y=1.16 $X2=0
+ $Y2=0
cc_216 N_A1_N_c_222_n N_A_113_47#_c_304_n 0.0143012f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A1_N_c_223_n N_A_113_47#_c_304_n 0.00156252f $X=3.43 $Y=1.16 $X2=0
+ $Y2=0
cc_218 N_A1_N_c_222_n N_A_113_47#_c_321_n 0.0204549f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A1_N_c_223_n N_A_113_47#_c_321_n 0.00220041f $X=3.43 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A1_N_c_222_n N_A_113_47#_c_322_n 0.0204549f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A1_N_c_223_n N_A_113_47#_c_322_n 0.00220041f $X=3.43 $Y=1.16 $X2=0
+ $Y2=0
cc_222 N_A1_N_M1004_g N_VPWR_c_612_n 0.00157837f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A1_N_M1015_g N_VPWR_c_613_n 0.00157837f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A1_N_M1016_g N_VPWR_c_613_n 0.00157837f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A1_N_M1026_g N_VPWR_c_614_n 0.00352998f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A1_N_M1004_g N_VPWR_c_622_n 0.00585385f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A1_N_M1015_g N_VPWR_c_622_n 0.00585385f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A1_N_M1016_g N_VPWR_c_631_n 0.00585385f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A1_N_M1026_g N_VPWR_c_631_n 0.00585385f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_230 N_A1_N_M1004_g N_VPWR_c_608_n 0.010464f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A1_N_M1015_g N_VPWR_c_608_n 0.0104367f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A1_N_M1016_g N_VPWR_c_608_n 0.0104367f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A1_N_M1026_g N_VPWR_c_608_n 0.0117628f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A1_N_c_218_n N_A_27_47#_c_918_n 0.00255288f $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A1_N_c_218_n N_A_27_47#_c_908_n 0.0048497f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A1_N_c_219_n N_A_27_47#_c_908_n 4.58193e-19 $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A1_N_c_222_n N_A_27_47#_c_908_n 0.00231036f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A1_N_c_218_n N_A_27_47#_c_909_n 0.00870364f $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_239 N_A1_N_c_219_n N_A_27_47#_c_909_n 0.00865686f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_240 N_A1_N_c_222_n N_A_27_47#_c_909_n 0.0362443f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A1_N_c_223_n N_A_27_47#_c_909_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A1_N_c_218_n N_A_27_47#_c_926_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A1_N_c_219_n N_A_27_47#_c_926_n 0.00630972f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A1_N_c_220_n N_A_27_47#_c_926_n 0.00630972f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A1_N_c_221_n N_A_27_47#_c_926_n 5.22228e-19 $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A1_N_c_220_n N_A_27_47#_c_910_n 0.00870364f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A1_N_c_221_n N_A_27_47#_c_910_n 0.00999903f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A1_N_c_222_n N_A_27_47#_c_910_n 0.038555f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_N_c_223_n N_A_27_47#_c_910_n 0.00222133f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A1_N_c_220_n N_A_27_47#_c_911_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A1_N_c_221_n N_A_27_47#_c_911_n 0.00630972f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A1_N_c_219_n N_A_27_47#_c_912_n 0.00113286f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A1_N_c_220_n N_A_27_47#_c_912_n 0.00113286f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A1_N_c_222_n N_A_27_47#_c_912_n 0.0266272f $X=3.28 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A1_N_c_223_n N_A_27_47#_c_912_n 0.00230339f $X=3.43 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A1_N_c_218_n N_VGND_c_980_n 0.00268723f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A1_N_c_219_n N_VGND_c_980_n 0.00146448f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A1_N_c_220_n N_VGND_c_981_n 0.00146448f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_N_c_221_n N_VGND_c_981_n 0.00268723f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A1_N_c_218_n N_VGND_c_986_n 0.00421816f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A1_N_c_219_n N_VGND_c_988_n 0.00423334f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A1_N_c_220_n N_VGND_c_988_n 0.00423334f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A1_N_c_221_n N_VGND_c_994_n 0.00423334f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A1_N_c_218_n N_VGND_c_997_n 0.00575258f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A1_N_c_219_n N_VGND_c_997_n 0.0057163f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A1_N_c_220_n N_VGND_c_997_n 0.0057163f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_N_c_221_n N_VGND_c_997_n 0.00704237f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_113_47#_c_312_n N_VPWR_M1005_s 0.00108428f $X=0.575 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_269 N_A_113_47#_c_313_n N_VPWR_M1005_s 0.00281778f $X=0.255 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_270 N_A_113_47#_c_314_n N_VPWR_M1021_s 0.00165831f $X=1.415 $Y=1.54 $X2=0
+ $Y2=0
cc_271 N_A_113_47#_c_315_n N_VPWR_M1034_s 0.00165831f $X=2.255 $Y=1.54 $X2=0
+ $Y2=0
cc_272 N_A_113_47#_c_316_n N_VPWR_M1015_d 0.00165831f $X=3.095 $Y=1.54 $X2=0
+ $Y2=0
cc_273 N_A_113_47#_c_317_n N_VPWR_M1026_d 0.00768298f $X=3.745 $Y=1.54 $X2=0
+ $Y2=0
cc_274 N_A_113_47#_c_312_n N_VPWR_c_610_n 0.00834345f $X=0.575 $Y=1.54 $X2=0
+ $Y2=0
cc_275 N_A_113_47#_c_313_n N_VPWR_c_610_n 0.00892602f $X=0.255 $Y=1.54 $X2=0
+ $Y2=0
cc_276 N_A_113_47#_c_314_n N_VPWR_c_611_n 0.0126919f $X=1.415 $Y=1.54 $X2=0
+ $Y2=0
cc_277 N_A_113_47#_c_315_n N_VPWR_c_612_n 0.0126919f $X=2.255 $Y=1.54 $X2=0
+ $Y2=0
cc_278 N_A_113_47#_c_316_n N_VPWR_c_613_n 0.0126919f $X=3.095 $Y=1.54 $X2=0
+ $Y2=0
cc_279 N_A_113_47#_M1001_g N_VPWR_c_614_n 0.00352998f $X=4.34 $Y=1.985 $X2=0
+ $Y2=0
cc_280 N_A_113_47#_c_317_n N_VPWR_c_614_n 0.0299422f $X=3.745 $Y=1.54 $X2=0
+ $Y2=0
cc_281 N_A_113_47#_c_305_n N_VPWR_c_614_n 0.0119603f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_113_47#_M1006_g N_VPWR_c_615_n 0.00157837f $X=4.76 $Y=1.985 $X2=0
+ $Y2=0
cc_283 N_A_113_47#_M1022_g N_VPWR_c_615_n 0.00157837f $X=5.18 $Y=1.985 $X2=0
+ $Y2=0
cc_284 N_A_113_47#_M1022_g N_VPWR_c_616_n 0.00585385f $X=5.18 $Y=1.985 $X2=0
+ $Y2=0
cc_285 N_A_113_47#_M1028_g N_VPWR_c_616_n 0.00585385f $X=5.6 $Y=1.985 $X2=0
+ $Y2=0
cc_286 N_A_113_47#_M1028_g N_VPWR_c_617_n 0.00338128f $X=5.6 $Y=1.985 $X2=0
+ $Y2=0
cc_287 N_A_113_47#_c_378_p N_VPWR_c_620_n 0.0142343f $X=1.54 $Y=2.3 $X2=0 $Y2=0
cc_288 N_A_113_47#_c_379_p N_VPWR_c_622_n 0.0142343f $X=2.38 $Y=2.3 $X2=0 $Y2=0
cc_289 N_A_113_47#_M1001_g N_VPWR_c_624_n 0.00585385f $X=4.34 $Y=1.985 $X2=0
+ $Y2=0
cc_290 N_A_113_47#_M1006_g N_VPWR_c_624_n 0.00585385f $X=4.76 $Y=1.985 $X2=0
+ $Y2=0
cc_291 N_A_113_47#_c_382_p N_VPWR_c_630_n 0.0142343f $X=0.7 $Y=2.3 $X2=0 $Y2=0
cc_292 N_A_113_47#_c_383_p N_VPWR_c_631_n 0.0142343f $X=3.22 $Y=2.3 $X2=0 $Y2=0
cc_293 N_A_113_47#_M1005_d N_VPWR_c_608_n 0.00284632f $X=0.565 $Y=1.485 $X2=0
+ $Y2=0
cc_294 N_A_113_47#_M1025_d N_VPWR_c_608_n 0.00284632f $X=1.405 $Y=1.485 $X2=0
+ $Y2=0
cc_295 N_A_113_47#_M1004_s N_VPWR_c_608_n 0.00284632f $X=2.245 $Y=1.485 $X2=0
+ $Y2=0
cc_296 N_A_113_47#_M1016_s N_VPWR_c_608_n 0.00284632f $X=3.085 $Y=1.485 $X2=0
+ $Y2=0
cc_297 N_A_113_47#_M1001_g N_VPWR_c_608_n 0.0117628f $X=4.34 $Y=1.985 $X2=0
+ $Y2=0
cc_298 N_A_113_47#_M1006_g N_VPWR_c_608_n 0.0104367f $X=4.76 $Y=1.985 $X2=0
+ $Y2=0
cc_299 N_A_113_47#_M1022_g N_VPWR_c_608_n 0.0104367f $X=5.18 $Y=1.985 $X2=0
+ $Y2=0
cc_300 N_A_113_47#_M1028_g N_VPWR_c_608_n 0.0117628f $X=5.6 $Y=1.985 $X2=0 $Y2=0
cc_301 N_A_113_47#_c_382_p N_VPWR_c_608_n 0.00955092f $X=0.7 $Y=2.3 $X2=0 $Y2=0
cc_302 N_A_113_47#_c_378_p N_VPWR_c_608_n 0.00955092f $X=1.54 $Y=2.3 $X2=0 $Y2=0
cc_303 N_A_113_47#_c_379_p N_VPWR_c_608_n 0.00955092f $X=2.38 $Y=2.3 $X2=0 $Y2=0
cc_304 N_A_113_47#_c_383_p N_VPWR_c_608_n 0.00955092f $X=3.22 $Y=2.3 $X2=0 $Y2=0
cc_305 N_A_113_47#_c_296_n N_Y_c_758_n 0.00460086f $X=4.37 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_113_47#_c_297_n N_Y_c_758_n 0.0109625f $X=4.79 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_113_47#_c_298_n N_Y_c_758_n 0.0109625f $X=5.21 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_113_47#_c_299_n N_Y_c_758_n 0.0136645f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_113_47#_c_305_n N_Y_c_758_n 0.0950491f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_113_47#_c_306_n N_Y_c_758_n 0.00711324f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_113_47#_M1001_g N_Y_c_760_n 4.51254e-19 $X=4.34 $Y=1.985 $X2=0 $Y2=0
cc_312 N_A_113_47#_c_317_n N_Y_c_760_n 0.00405228f $X=3.745 $Y=1.54 $X2=0 $Y2=0
cc_313 N_A_113_47#_c_305_n N_Y_c_760_n 0.0204549f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_113_47#_c_306_n N_Y_c_760_n 0.00232398f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_113_47#_M1006_g N_Y_c_761_n 0.0132131f $X=4.76 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_113_47#_M1022_g N_Y_c_761_n 0.0132273f $X=5.18 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A_113_47#_c_305_n N_Y_c_761_n 0.0416643f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_113_47#_c_306_n N_Y_c_761_n 0.00223852f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_113_47#_M1028_g N_Y_c_762_n 0.0153744f $X=5.6 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_113_47#_c_305_n N_Y_c_762_n 0.0132031f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_113_47#_c_306_n N_Y_c_762_n 8.28465e-19 $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_113_47#_M1028_g N_Y_c_759_n 0.00453969f $X=5.6 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_113_47#_c_299_n N_Y_c_759_n 0.00676796f $X=5.63 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_113_47#_c_305_n N_Y_c_759_n 0.0172409f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_113_47#_c_306_n N_Y_c_759_n 0.00329028f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_113_47#_c_305_n N_Y_c_766_n 0.0204549f $X=5.48 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_113_47#_c_306_n N_Y_c_766_n 0.00232398f $X=5.63 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_113_47#_c_301_n N_A_27_47#_M1008_s 0.00261124f $X=0.255 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_329 N_A_113_47#_c_302_n N_A_27_47#_M1008_s 0.00106131f $X=1.54 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_330 N_A_113_47#_c_302_n N_A_27_47#_M1012_s 0.00162317f $X=1.54 $Y=0.73 $X2=0
+ $Y2=0
cc_331 N_A_113_47#_M1008_d N_A_27_47#_c_907_n 0.00305026f $X=0.565 $Y=0.235
+ $X2=0 $Y2=0
cc_332 N_A_113_47#_M1017_d N_A_27_47#_c_907_n 0.00305026f $X=1.405 $Y=0.235
+ $X2=0 $Y2=0
cc_333 N_A_113_47#_c_301_n N_A_27_47#_c_907_n 0.0122591f $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_334 N_A_113_47#_c_302_n N_A_27_47#_c_907_n 0.0737784f $X=1.54 $Y=0.73 $X2=0
+ $Y2=0
cc_335 N_A_113_47#_c_302_n N_A_27_47#_c_908_n 0.00841895f $X=1.54 $Y=0.73 $X2=0
+ $Y2=0
cc_336 N_A_113_47#_c_315_n N_A_27_47#_c_908_n 0.00817864f $X=2.255 $Y=1.54 $X2=0
+ $Y2=0
cc_337 N_A_113_47#_c_296_n N_A_27_47#_c_910_n 0.00149957f $X=4.37 $Y=0.995 $X2=0
+ $Y2=0
cc_338 N_A_113_47#_c_317_n N_A_27_47#_c_910_n 0.00890545f $X=3.745 $Y=1.54 $X2=0
+ $Y2=0
cc_339 N_A_113_47#_c_304_n N_A_27_47#_c_910_n 0.00551491f $X=3.915 $Y=1.18 $X2=0
+ $Y2=0
cc_340 N_A_113_47#_c_296_n N_A_27_47#_c_911_n 7.52656e-19 $X=4.37 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_113_47#_c_301_n N_VGND_c_986_n 2.98364e-19 $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_342 N_A_113_47#_c_296_n N_VGND_c_994_n 0.00357877f $X=4.37 $Y=0.995 $X2=0
+ $Y2=0
cc_343 N_A_113_47#_c_297_n N_VGND_c_994_n 0.00357877f $X=4.79 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_113_47#_c_298_n N_VGND_c_994_n 0.00357877f $X=5.21 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_113_47#_c_299_n N_VGND_c_994_n 0.00357877f $X=5.63 $Y=0.995 $X2=0
+ $Y2=0
cc_346 N_A_113_47#_M1008_d N_VGND_c_997_n 0.00216833f $X=0.565 $Y=0.235 $X2=0
+ $Y2=0
cc_347 N_A_113_47#_M1017_d N_VGND_c_997_n 0.00216833f $X=1.405 $Y=0.235 $X2=0
+ $Y2=0
cc_348 N_A_113_47#_c_296_n N_VGND_c_997_n 0.00664112f $X=4.37 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_113_47#_c_297_n N_VGND_c_997_n 0.00522516f $X=4.79 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_113_47#_c_298_n N_VGND_c_997_n 0.00522516f $X=5.21 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_113_47#_c_299_n N_VGND_c_997_n 0.00655123f $X=5.63 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_113_47#_c_301_n N_VGND_c_997_n 8.363e-19 $X=0.255 $Y=0.775 $X2=0
+ $Y2=0
cc_353 N_A_113_47#_c_305_n N_A_807_47#_c_1131_n 0.0116182f $X=5.48 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_A_113_47#_c_296_n N_A_807_47#_c_1132_n 0.0130436f $X=4.37 $Y=0.995
+ $X2=0 $Y2=0
cc_355 N_A_113_47#_c_297_n N_A_807_47#_c_1132_n 0.00886996f $X=4.79 $Y=0.995
+ $X2=0 $Y2=0
cc_356 N_A_113_47#_c_298_n N_A_807_47#_c_1132_n 0.00892725f $X=5.21 $Y=0.995
+ $X2=0 $Y2=0
cc_357 N_A_113_47#_c_299_n N_A_807_47#_c_1132_n 0.00892725f $X=5.63 $Y=0.995
+ $X2=0 $Y2=0
cc_358 N_A_113_47#_c_305_n N_A_807_47#_c_1132_n 0.00365276f $X=5.48 $Y=1.16
+ $X2=0 $Y2=0
cc_359 N_A_113_47#_c_299_n N_A_807_47#_c_1137_n 0.00274112f $X=5.63 $Y=0.995
+ $X2=0 $Y2=0
cc_360 N_A_113_47#_c_299_n N_A_807_47#_c_1123_n 5.50017e-19 $X=5.63 $Y=0.995
+ $X2=0 $Y2=0
cc_361 N_B2_c_455_n N_B1_c_533_n 0.015126f $X=7.8 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_362 N_B2_M1036_g N_B1_M1018_g 0.015126f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_363 N_B2_c_464_p N_B1_c_537_n 0.0184614f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_364 N_B2_c_456_n N_B1_c_537_n 0.00159737f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_365 N_B2_c_464_p N_B1_c_538_n 2.16609e-19 $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_366 N_B2_c_456_n N_B1_c_538_n 0.015126f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_367 N_B2_M1003_g N_VPWR_c_617_n 0.00214918f $X=6.54 $Y=1.985 $X2=0 $Y2=0
cc_368 N_B2_M1003_g N_VPWR_c_626_n 0.00357877f $X=6.54 $Y=1.985 $X2=0 $Y2=0
cc_369 N_B2_M1010_g N_VPWR_c_626_n 0.00357877f $X=6.96 $Y=1.985 $X2=0 $Y2=0
cc_370 N_B2_M1033_g N_VPWR_c_626_n 0.00357877f $X=7.38 $Y=1.985 $X2=0 $Y2=0
cc_371 N_B2_M1036_g N_VPWR_c_626_n 0.00357877f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_372 N_B2_M1003_g N_VPWR_c_608_n 0.00655123f $X=6.54 $Y=1.985 $X2=0 $Y2=0
cc_373 N_B2_M1010_g N_VPWR_c_608_n 0.00522516f $X=6.96 $Y=1.985 $X2=0 $Y2=0
cc_374 N_B2_M1033_g N_VPWR_c_608_n 0.00522516f $X=7.38 $Y=1.985 $X2=0 $Y2=0
cc_375 N_B2_M1036_g N_VPWR_c_608_n 0.00525237f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_376 N_B2_c_452_n N_Y_c_758_n 0.00149512f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_377 N_B2_c_452_n N_Y_c_759_n 0.0163848f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_378 N_B2_c_464_p N_Y_c_759_n 0.0110646f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_379 N_B2_M1003_g N_Y_c_764_n 0.0130673f $X=6.54 $Y=1.985 $X2=0 $Y2=0
cc_380 N_B2_c_464_p N_Y_c_764_n 0.011015f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_381 N_B2_M1010_g N_Y_c_765_n 0.0109338f $X=6.96 $Y=1.985 $X2=0 $Y2=0
cc_382 N_B2_M1033_g N_Y_c_765_n 0.0109196f $X=7.38 $Y=1.985 $X2=0 $Y2=0
cc_383 N_B2_c_464_p N_Y_c_765_n 0.0418862f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_384 N_B2_c_456_n N_Y_c_765_n 0.00211393f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_385 N_B2_c_464_p N_Y_c_768_n 0.020533f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_386 N_B2_c_456_n N_Y_c_768_n 0.00219397f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B2_M1036_g N_Y_c_769_n 2.57315e-19 $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_388 N_B2_c_464_p N_Y_c_769_n 0.020533f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_389 N_B2_c_456_n N_Y_c_769_n 0.00219397f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_390 N_B2_M1003_g N_A_1241_297#_c_852_n 0.00988743f $X=6.54 $Y=1.985 $X2=0
+ $Y2=0
cc_391 N_B2_M1010_g N_A_1241_297#_c_852_n 0.00984328f $X=6.96 $Y=1.985 $X2=0
+ $Y2=0
cc_392 N_B2_M1033_g N_A_1241_297#_c_854_n 0.00984328f $X=7.38 $Y=1.985 $X2=0
+ $Y2=0
cc_393 N_B2_M1036_g N_A_1241_297#_c_854_n 0.0121747f $X=7.8 $Y=1.985 $X2=0 $Y2=0
cc_394 N_B2_M1036_g N_A_1241_297#_c_846_n 2.57315e-19 $X=7.8 $Y=1.985 $X2=0
+ $Y2=0
cc_395 N_B2_c_452_n N_VGND_c_982_n 0.00268723f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_396 N_B2_c_453_n N_VGND_c_982_n 0.00146448f $X=6.96 $Y=0.995 $X2=0 $Y2=0
cc_397 N_B2_c_454_n N_VGND_c_983_n 0.00146448f $X=7.38 $Y=0.995 $X2=0 $Y2=0
cc_398 N_B2_c_455_n N_VGND_c_983_n 0.00146448f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B2_c_455_n N_VGND_c_990_n 0.00423334f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_400 N_B2_c_452_n N_VGND_c_994_n 0.00422898f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_401 N_B2_c_453_n N_VGND_c_995_n 0.00424416f $X=6.96 $Y=0.995 $X2=0 $Y2=0
cc_402 N_B2_c_454_n N_VGND_c_995_n 0.00423334f $X=7.38 $Y=0.995 $X2=0 $Y2=0
cc_403 N_B2_c_452_n N_VGND_c_997_n 0.00707121f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_404 N_B2_c_453_n N_VGND_c_997_n 0.00573607f $X=6.96 $Y=0.995 $X2=0 $Y2=0
cc_405 N_B2_c_454_n N_VGND_c_997_n 0.0057163f $X=7.38 $Y=0.995 $X2=0 $Y2=0
cc_406 N_B2_c_455_n N_VGND_c_997_n 0.0057435f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B2_c_452_n N_A_807_47#_c_1139_n 0.00255288f $X=6.54 $Y=0.995 $X2=0
+ $Y2=0
cc_408 N_B2_c_452_n N_A_807_47#_c_1137_n 0.0065045f $X=6.54 $Y=0.995 $X2=0 $Y2=0
cc_409 N_B2_c_453_n N_A_807_47#_c_1137_n 4.89212e-19 $X=6.96 $Y=0.995 $X2=0
+ $Y2=0
cc_410 N_B2_c_452_n N_A_807_47#_c_1122_n 0.00849697f $X=6.54 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_B2_c_453_n N_A_807_47#_c_1122_n 0.00845282f $X=6.96 $Y=0.995 $X2=0
+ $Y2=0
cc_412 N_B2_c_464_p N_A_807_47#_c_1122_n 0.036276f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_413 N_B2_c_456_n N_A_807_47#_c_1122_n 0.00221699f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_414 N_B2_c_452_n N_A_807_47#_c_1123_n 0.00381348f $X=6.54 $Y=0.995 $X2=0
+ $Y2=0
cc_415 N_B2_c_464_p N_A_807_47#_c_1123_n 0.00224551f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_416 N_B2_c_452_n N_A_807_47#_c_1148_n 5.22228e-19 $X=6.54 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_B2_c_453_n N_A_807_47#_c_1148_n 0.00630972f $X=6.96 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_B2_c_454_n N_A_807_47#_c_1148_n 0.00630972f $X=7.38 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_B2_c_455_n N_A_807_47#_c_1148_n 5.22228e-19 $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_420 N_B2_c_454_n N_A_807_47#_c_1124_n 0.00869873f $X=7.38 $Y=0.995 $X2=0
+ $Y2=0
cc_421 N_B2_c_455_n N_A_807_47#_c_1124_n 0.00869873f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_422 N_B2_c_464_p N_A_807_47#_c_1124_n 0.0364367f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_423 N_B2_c_456_n N_A_807_47#_c_1124_n 0.00222006f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_424 N_B2_c_454_n N_A_807_47#_c_1156_n 5.22228e-19 $X=7.38 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_B2_c_455_n N_A_807_47#_c_1156_n 0.00630972f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_426 N_B2_c_453_n N_A_807_47#_c_1128_n 0.00127881f $X=6.96 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_B2_c_454_n N_A_807_47#_c_1128_n 0.00113159f $X=7.38 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_B2_c_464_p N_A_807_47#_c_1128_n 0.0267643f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_429 N_B2_c_456_n N_A_807_47#_c_1128_n 0.00230167f $X=7.8 $Y=1.16 $X2=0 $Y2=0
cc_430 N_B2_c_455_n N_A_807_47#_c_1129_n 0.00111217f $X=7.8 $Y=0.995 $X2=0 $Y2=0
cc_431 N_B2_c_464_p N_A_807_47#_c_1129_n 0.0022458f $X=6.63 $Y=1.16 $X2=0 $Y2=0
cc_432 N_B1_M1018_g N_VPWR_c_618_n 0.00302074f $X=8.22 $Y=1.985 $X2=0 $Y2=0
cc_433 N_B1_M1029_g N_VPWR_c_618_n 0.00157837f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_434 N_B1_M1030_g N_VPWR_c_619_n 0.00157837f $X=9.06 $Y=1.985 $X2=0 $Y2=0
cc_435 N_B1_M1037_g N_VPWR_c_619_n 0.00302074f $X=9.48 $Y=1.985 $X2=0 $Y2=0
cc_436 N_B1_M1018_g N_VPWR_c_626_n 0.00585385f $X=8.22 $Y=1.985 $X2=0 $Y2=0
cc_437 N_B1_M1029_g N_VPWR_c_628_n 0.00585385f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_438 N_B1_M1030_g N_VPWR_c_628_n 0.00585385f $X=9.06 $Y=1.985 $X2=0 $Y2=0
cc_439 N_B1_M1037_g N_VPWR_c_632_n 0.00585385f $X=9.48 $Y=1.985 $X2=0 $Y2=0
cc_440 N_B1_M1018_g N_VPWR_c_608_n 0.010464f $X=8.22 $Y=1.985 $X2=0 $Y2=0
cc_441 N_B1_M1029_g N_VPWR_c_608_n 0.0104367f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_442 N_B1_M1030_g N_VPWR_c_608_n 0.0104367f $X=9.06 $Y=1.985 $X2=0 $Y2=0
cc_443 N_B1_M1037_g N_VPWR_c_608_n 0.0115188f $X=9.48 $Y=1.985 $X2=0 $Y2=0
cc_444 N_B1_c_537_n N_A_1241_297#_c_846_n 0.00771248f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_445 N_B1_M1018_g N_A_1241_297#_c_847_n 0.0132131f $X=8.22 $Y=1.985 $X2=0
+ $Y2=0
cc_446 N_B1_M1029_g N_A_1241_297#_c_847_n 0.0132273f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_447 N_B1_c_537_n N_A_1241_297#_c_847_n 0.041703f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_448 N_B1_c_538_n N_A_1241_297#_c_847_n 0.00211509f $X=9.48 $Y=1.16 $X2=0
+ $Y2=0
cc_449 N_B1_M1030_g N_A_1241_297#_c_848_n 0.0132714f $X=9.06 $Y=1.985 $X2=0
+ $Y2=0
cc_450 N_B1_M1037_g N_A_1241_297#_c_848_n 0.0135194f $X=9.48 $Y=1.985 $X2=0
+ $Y2=0
cc_451 N_B1_c_537_n N_A_1241_297#_c_848_n 0.041703f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_452 N_B1_c_538_n N_A_1241_297#_c_848_n 0.00211509f $X=9.48 $Y=1.16 $X2=0
+ $Y2=0
cc_453 N_B1_c_537_n N_A_1241_297#_c_849_n 0.0265652f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_454 N_B1_c_537_n N_A_1241_297#_c_851_n 0.0204549f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_455 N_B1_c_538_n N_A_1241_297#_c_851_n 0.00220041f $X=9.48 $Y=1.16 $X2=0
+ $Y2=0
cc_456 N_B1_c_533_n N_VGND_c_984_n 0.00146448f $X=8.22 $Y=0.995 $X2=0 $Y2=0
cc_457 N_B1_c_534_n N_VGND_c_984_n 0.00146448f $X=8.64 $Y=0.995 $X2=0 $Y2=0
cc_458 N_B1_c_535_n N_VGND_c_985_n 0.00146448f $X=9.06 $Y=0.995 $X2=0 $Y2=0
cc_459 N_B1_c_536_n N_VGND_c_985_n 0.00268723f $X=9.48 $Y=0.995 $X2=0 $Y2=0
cc_460 N_B1_c_533_n N_VGND_c_990_n 0.00423334f $X=8.22 $Y=0.995 $X2=0 $Y2=0
cc_461 N_B1_c_534_n N_VGND_c_992_n 0.00423334f $X=8.64 $Y=0.995 $X2=0 $Y2=0
cc_462 N_B1_c_535_n N_VGND_c_992_n 0.00423334f $X=9.06 $Y=0.995 $X2=0 $Y2=0
cc_463 N_B1_c_536_n N_VGND_c_996_n 0.00423334f $X=9.48 $Y=0.995 $X2=0 $Y2=0
cc_464 N_B1_c_533_n N_VGND_c_997_n 0.0057435f $X=8.22 $Y=0.995 $X2=0 $Y2=0
cc_465 N_B1_c_534_n N_VGND_c_997_n 0.0057163f $X=8.64 $Y=0.995 $X2=0 $Y2=0
cc_466 N_B1_c_535_n N_VGND_c_997_n 0.0057163f $X=9.06 $Y=0.995 $X2=0 $Y2=0
cc_467 N_B1_c_536_n N_VGND_c_997_n 0.00679836f $X=9.48 $Y=0.995 $X2=0 $Y2=0
cc_468 N_B1_c_533_n N_A_807_47#_c_1156_n 0.00630972f $X=8.22 $Y=0.995 $X2=0
+ $Y2=0
cc_469 N_B1_c_534_n N_A_807_47#_c_1156_n 5.22228e-19 $X=8.64 $Y=0.995 $X2=0
+ $Y2=0
cc_470 N_B1_c_533_n N_A_807_47#_c_1125_n 0.00870364f $X=8.22 $Y=0.995 $X2=0
+ $Y2=0
cc_471 N_B1_c_534_n N_A_807_47#_c_1125_n 0.00870364f $X=8.64 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_B1_c_537_n N_A_807_47#_c_1125_n 0.0362443f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_473 N_B1_c_538_n N_A_807_47#_c_1125_n 0.00222133f $X=9.48 $Y=1.16 $X2=0 $Y2=0
cc_474 N_B1_c_533_n N_A_807_47#_c_1170_n 5.22228e-19 $X=8.22 $Y=0.995 $X2=0
+ $Y2=0
cc_475 N_B1_c_534_n N_A_807_47#_c_1170_n 0.00630972f $X=8.64 $Y=0.995 $X2=0
+ $Y2=0
cc_476 N_B1_c_535_n N_A_807_47#_c_1170_n 0.00630972f $X=9.06 $Y=0.995 $X2=0
+ $Y2=0
cc_477 N_B1_c_536_n N_A_807_47#_c_1170_n 5.22228e-19 $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_B1_c_535_n N_A_807_47#_c_1126_n 0.00870364f $X=9.06 $Y=0.995 $X2=0
+ $Y2=0
cc_479 N_B1_c_536_n N_A_807_47#_c_1126_n 0.00999903f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_B1_c_537_n N_A_807_47#_c_1126_n 0.0641689f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_481 N_B1_c_538_n N_A_807_47#_c_1126_n 0.00222133f $X=9.48 $Y=1.16 $X2=0 $Y2=0
cc_482 N_B1_c_535_n N_A_807_47#_c_1127_n 5.22228e-19 $X=9.06 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_B1_c_536_n N_A_807_47#_c_1127_n 0.00630972f $X=9.48 $Y=0.995 $X2=0
+ $Y2=0
cc_484 N_B1_c_533_n N_A_807_47#_c_1129_n 0.00112787f $X=8.22 $Y=0.995 $X2=0
+ $Y2=0
cc_485 N_B1_c_537_n N_A_807_47#_c_1129_n 0.0108485f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_486 N_B1_c_534_n N_A_807_47#_c_1130_n 0.00113286f $X=8.64 $Y=0.995 $X2=0
+ $Y2=0
cc_487 N_B1_c_535_n N_A_807_47#_c_1130_n 0.00113286f $X=9.06 $Y=0.995 $X2=0
+ $Y2=0
cc_488 N_B1_c_537_n N_A_807_47#_c_1130_n 0.0266272f $X=9.3 $Y=1.16 $X2=0 $Y2=0
cc_489 N_B1_c_538_n N_A_807_47#_c_1130_n 0.00230339f $X=9.48 $Y=1.16 $X2=0 $Y2=0
cc_490 N_VPWR_c_608_n N_Y_M1001_s 0.00284632f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_491 N_VPWR_c_608_n N_Y_M1022_s 0.00284632f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_492 N_VPWR_c_608_n N_Y_M1003_s 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_493 N_VPWR_c_608_n N_Y_M1033_s 0.00216833f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_494 N_VPWR_c_624_n N_Y_c_811_n 0.0142343f $X=4.845 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_c_608_n N_Y_c_811_n 0.00955092f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_496 N_VPWR_M1006_d N_Y_c_761_n 0.00165831f $X=4.835 $Y=1.485 $X2=0 $Y2=0
cc_497 N_VPWR_c_615_n N_Y_c_761_n 0.0126919f $X=4.97 $Y=1.96 $X2=0 $Y2=0
cc_498 N_VPWR_c_616_n N_Y_c_815_n 0.0142343f $X=5.685 $Y=2.72 $X2=0 $Y2=0
cc_499 N_VPWR_c_608_n N_Y_c_815_n 0.00955092f $X=9.89 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_M1028_d N_Y_c_762_n 0.00165567f $X=5.675 $Y=1.485 $X2=0 $Y2=0
cc_501 N_VPWR_c_617_n N_Y_c_762_n 0.0115978f $X=5.81 $Y=1.96 $X2=0 $Y2=0
cc_502 N_VPWR_M1028_d N_Y_c_767_n 0.00111785f $X=5.675 $Y=1.485 $X2=0 $Y2=0
cc_503 N_VPWR_c_617_n N_Y_c_767_n 0.00531954f $X=5.81 $Y=1.96 $X2=0 $Y2=0
cc_504 N_VPWR_c_608_n N_A_1241_297#_M1003_d 0.0020932f $X=9.89 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_505 N_VPWR_c_608_n N_A_1241_297#_M1010_d 0.00215203f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_608_n N_A_1241_297#_M1036_d 0.00246446f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_608_n N_A_1241_297#_M1029_d 0.00284632f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_608_n N_A_1241_297#_M1037_d 0.00260431f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_617_n N_A_1241_297#_c_844_n 0.0308495f $X=5.81 $Y=1.96 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_626_n N_A_1241_297#_c_852_n 0.0330174f $X=8.305 $Y=2.72 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_608_n N_A_1241_297#_c_852_n 0.0204627f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_617_n N_A_1241_297#_c_845_n 0.0113145f $X=5.81 $Y=1.96 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_626_n N_A_1241_297#_c_845_n 0.0180757f $X=8.305 $Y=2.72 $X2=0
+ $Y2=0
cc_514 N_VPWR_c_608_n N_A_1241_297#_c_845_n 0.0107791f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_626_n N_A_1241_297#_c_854_n 0.0330174f $X=8.305 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_608_n N_A_1241_297#_c_854_n 0.0204627f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_626_n N_A_1241_297#_c_882_n 0.0143053f $X=8.305 $Y=2.72 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_608_n N_A_1241_297#_c_882_n 0.00962794f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_519 N_VPWR_M1018_s N_A_1241_297#_c_847_n 0.00165831f $X=8.295 $Y=1.485 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_618_n N_A_1241_297#_c_847_n 0.0126919f $X=8.43 $Y=1.96 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_628_n N_A_1241_297#_c_886_n 0.0142343f $X=9.145 $Y=2.72 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_608_n N_A_1241_297#_c_886_n 0.00955092f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_523 N_VPWR_M1030_s N_A_1241_297#_c_848_n 0.00165831f $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_619_n N_A_1241_297#_c_848_n 0.0126919f $X=9.27 $Y=1.96 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_632_n N_A_1241_297#_c_850_n 0.0201098f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_608_n N_A_1241_297#_c_850_n 0.0118616f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_626_n N_A_1241_297#_c_892_n 0.0142933f $X=8.305 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_608_n N_A_1241_297#_c_892_n 0.00962421f $X=9.89 $Y=2.72 $X2=0
+ $Y2=0
cc_529 N_Y_c_764_n N_A_1241_297#_M1003_d 0.00277342f $X=6.625 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_530 N_Y_c_765_n N_A_1241_297#_M1010_d 0.00165831f $X=7.465 $Y=1.54 $X2=0
+ $Y2=0
cc_531 N_Y_c_764_n N_A_1241_297#_c_844_n 0.0189421f $X=6.625 $Y=1.54 $X2=0 $Y2=0
cc_532 N_Y_M1003_s N_A_1241_297#_c_852_n 0.00312348f $X=6.615 $Y=1.485 $X2=0
+ $Y2=0
cc_533 N_Y_c_764_n N_A_1241_297#_c_852_n 0.00320918f $X=6.625 $Y=1.54 $X2=0
+ $Y2=0
cc_534 N_Y_c_765_n N_A_1241_297#_c_852_n 0.00320918f $X=7.465 $Y=1.54 $X2=0
+ $Y2=0
cc_535 N_Y_c_768_n N_A_1241_297#_c_852_n 0.0118729f $X=6.75 $Y=1.62 $X2=0 $Y2=0
cc_536 N_Y_c_765_n N_A_1241_297#_c_901_n 0.0126766f $X=7.465 $Y=1.54 $X2=0 $Y2=0
cc_537 N_Y_M1033_s N_A_1241_297#_c_854_n 0.00312348f $X=7.455 $Y=1.485 $X2=0
+ $Y2=0
cc_538 N_Y_c_765_n N_A_1241_297#_c_854_n 0.00320918f $X=7.465 $Y=1.54 $X2=0
+ $Y2=0
cc_539 Y N_A_1241_297#_c_854_n 0.0118729f $X=7.505 $Y=1.785 $X2=0 $Y2=0
cc_540 N_Y_c_769_n N_A_1241_297#_c_846_n 0.00271526f $X=7.59 $Y=1.625 $X2=0
+ $Y2=0
cc_541 N_Y_c_758_n N_A_27_47#_c_910_n 0.00232529f $X=5.875 $Y=0.775 $X2=0 $Y2=0
cc_542 N_Y_M1007_s N_VGND_c_997_n 0.00216833f $X=4.445 $Y=0.235 $X2=0 $Y2=0
cc_543 N_Y_M1011_s N_VGND_c_997_n 0.00216833f $X=5.285 $Y=0.235 $X2=0 $Y2=0
cc_544 N_Y_c_758_n N_A_807_47#_M1009_d 0.00162317f $X=5.875 $Y=0.775 $X2=0 $Y2=0
cc_545 N_Y_c_758_n N_A_807_47#_M1013_d 0.00994839f $X=5.875 $Y=0.775 $X2=0 $Y2=0
cc_546 N_Y_M1007_s N_A_807_47#_c_1132_n 0.00305026f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_Y_M1011_s N_A_807_47#_c_1132_n 0.00305026f $X=5.285 $Y=0.235 $X2=0
+ $Y2=0
cc_548 N_Y_c_758_n N_A_807_47#_c_1132_n 0.0964603f $X=5.875 $Y=0.775 $X2=0 $Y2=0
cc_549 N_Y_c_758_n N_A_807_47#_c_1137_n 0.00728575f $X=5.875 $Y=0.775 $X2=0
+ $Y2=0
cc_550 N_Y_c_758_n N_A_807_47#_c_1123_n 0.015398f $X=5.875 $Y=0.775 $X2=0 $Y2=0
cc_551 N_Y_c_764_n N_A_807_47#_c_1123_n 0.00523344f $X=6.625 $Y=1.54 $X2=0 $Y2=0
cc_552 N_A_1241_297#_c_846_n N_A_807_47#_c_1129_n 0.00658191f $X=8.01 $Y=1.625
+ $X2=0 $Y2=0
cc_553 N_A_27_47#_c_909_n N_VGND_M1014_s 0.00162089f $X=2.635 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_554 N_A_27_47#_c_910_n N_VGND_M1023_s 0.00162089f $X=3.475 $Y=0.815 $X2=0
+ $Y2=0
cc_555 N_A_27_47#_c_909_n N_VGND_c_980_n 0.0122559f $X=2.635 $Y=0.815 $X2=0
+ $Y2=0
cc_556 N_A_27_47#_c_910_n N_VGND_c_981_n 0.0122559f $X=3.475 $Y=0.815 $X2=0
+ $Y2=0
cc_557 N_A_27_47#_c_907_n N_VGND_c_986_n 0.100139f $X=1.875 $Y=0.365 $X2=0 $Y2=0
cc_558 N_A_27_47#_c_918_n N_VGND_c_986_n 0.0152108f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_559 N_A_27_47#_c_909_n N_VGND_c_986_n 0.00198695f $X=2.635 $Y=0.815 $X2=0
+ $Y2=0
cc_560 N_A_27_47#_c_909_n N_VGND_c_988_n 0.00198695f $X=2.635 $Y=0.815 $X2=0
+ $Y2=0
cc_561 N_A_27_47#_c_926_n N_VGND_c_988_n 0.0188551f $X=2.8 $Y=0.39 $X2=0 $Y2=0
cc_562 N_A_27_47#_c_910_n N_VGND_c_988_n 0.00198695f $X=3.475 $Y=0.815 $X2=0
+ $Y2=0
cc_563 N_A_27_47#_c_910_n N_VGND_c_994_n 0.00198695f $X=3.475 $Y=0.815 $X2=0
+ $Y2=0
cc_564 N_A_27_47#_c_911_n N_VGND_c_994_n 0.0209752f $X=3.64 $Y=0.39 $X2=0 $Y2=0
cc_565 N_A_27_47#_M1008_s N_VGND_c_997_n 0.00225742f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_566 N_A_27_47#_M1012_s N_VGND_c_997_n 0.00215227f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_567 N_A_27_47#_M1019_s N_VGND_c_997_n 0.00215206f $X=1.825 $Y=0.235 $X2=0
+ $Y2=0
cc_568 N_A_27_47#_M1020_d N_VGND_c_997_n 0.00215201f $X=2.665 $Y=0.235 $X2=0
+ $Y2=0
cc_569 N_A_27_47#_M1027_d N_VGND_c_997_n 0.00209319f $X=3.505 $Y=0.235 $X2=0
+ $Y2=0
cc_570 N_A_27_47#_c_907_n N_VGND_c_997_n 0.0634607f $X=1.875 $Y=0.365 $X2=0
+ $Y2=0
cc_571 N_A_27_47#_c_918_n N_VGND_c_997_n 0.00940698f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_572 N_A_27_47#_c_909_n N_VGND_c_997_n 0.00835832f $X=2.635 $Y=0.815 $X2=0
+ $Y2=0
cc_573 N_A_27_47#_c_926_n N_VGND_c_997_n 0.0122069f $X=2.8 $Y=0.39 $X2=0 $Y2=0
cc_574 N_A_27_47#_c_910_n N_VGND_c_997_n 0.00835832f $X=3.475 $Y=0.815 $X2=0
+ $Y2=0
cc_575 N_A_27_47#_c_911_n N_VGND_c_997_n 0.0124119f $X=3.64 $Y=0.39 $X2=0 $Y2=0
cc_576 N_A_27_47#_c_910_n N_A_807_47#_c_1131_n 0.00687335f $X=3.475 $Y=0.815
+ $X2=0 $Y2=0
cc_577 N_A_27_47#_c_911_n N_A_807_47#_c_1131_n 0.01461f $X=3.64 $Y=0.39 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_c_911_n N_A_807_47#_c_1197_n 0.0142381f $X=3.64 $Y=0.39 $X2=0
+ $Y2=0
cc_579 N_VGND_c_997_n N_A_807_47#_M1007_d 0.00296916f $X=9.89 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_580 N_VGND_c_997_n N_A_807_47#_M1009_d 0.00215227f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_c_997_n N_A_807_47#_M1013_d 0.00615449f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_997_n N_A_807_47#_M1031_s 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_997_n N_A_807_47#_M1038_s 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_c_997_n N_A_807_47#_M1002_d 0.00215201f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_997_n N_A_807_47#_M1039_d 0.00209319f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_994_n N_A_807_47#_c_1132_n 0.119771f $X=6.665 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_997_n N_A_807_47#_c_1132_n 0.07495f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_994_n N_A_807_47#_c_1197_n 0.0126217f $X=6.665 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_997_n N_A_807_47#_c_1197_n 0.00709554f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_994_n N_A_807_47#_c_1139_n 0.00984597f $X=6.665 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_997_n N_A_807_47#_c_1139_n 0.00632969f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_M1024_d N_A_807_47#_c_1122_n 0.00165819f $X=6.615 $Y=0.235 $X2=0
+ $Y2=0
cc_593 N_VGND_c_982_n N_A_807_47#_c_1122_n 0.0116528f $X=6.75 $Y=0.39 $X2=0
+ $Y2=0
cc_594 N_VGND_c_994_n N_A_807_47#_c_1122_n 0.00193763f $X=6.665 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_995_n N_A_807_47#_c_1122_n 0.00193763f $X=7.505 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_997_n N_A_807_47#_c_1122_n 0.00827287f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_995_n N_A_807_47#_c_1148_n 0.0188551f $X=7.505 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_c_997_n N_A_807_47#_c_1148_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_599 N_VGND_M1032_d N_A_807_47#_c_1124_n 0.00162089f $X=7.455 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_VGND_c_983_n N_A_807_47#_c_1124_n 0.0122559f $X=7.59 $Y=0.39 $X2=0
+ $Y2=0
cc_601 N_VGND_c_990_n N_A_807_47#_c_1124_n 0.00198695f $X=8.345 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_995_n N_A_807_47#_c_1124_n 0.00198695f $X=7.505 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_997_n N_A_807_47#_c_1124_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_990_n N_A_807_47#_c_1156_n 0.0188551f $X=8.345 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_997_n N_A_807_47#_c_1156_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_M1000_s N_A_807_47#_c_1125_n 0.00162089f $X=8.295 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_VGND_c_984_n N_A_807_47#_c_1125_n 0.0122559f $X=8.43 $Y=0.39 $X2=0
+ $Y2=0
cc_608 N_VGND_c_990_n N_A_807_47#_c_1125_n 0.00198695f $X=8.345 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_c_992_n N_A_807_47#_c_1125_n 0.00198695f $X=9.185 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_997_n N_A_807_47#_c_1125_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_992_n N_A_807_47#_c_1170_n 0.0188551f $X=9.185 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_c_997_n N_A_807_47#_c_1170_n 0.0122069f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_M1035_s N_A_807_47#_c_1126_n 0.00162089f $X=9.135 $Y=0.235 $X2=0
+ $Y2=0
cc_614 N_VGND_c_985_n N_A_807_47#_c_1126_n 0.0122559f $X=9.27 $Y=0.39 $X2=0
+ $Y2=0
cc_615 N_VGND_c_992_n N_A_807_47#_c_1126_n 0.00198695f $X=9.185 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_996_n N_A_807_47#_c_1126_n 0.00198695f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_617 N_VGND_c_997_n N_A_807_47#_c_1126_n 0.00835832f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_996_n N_A_807_47#_c_1127_n 0.0209752f $X=9.89 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_997_n N_A_807_47#_c_1127_n 0.0124119f $X=9.89 $Y=0 $X2=0 $Y2=0

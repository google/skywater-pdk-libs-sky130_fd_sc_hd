* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
M1000 VPWR a_244_47# a_355_47# VPB phighvt w=820000u l=250000u
+  ad=9.305e+11p pd=6.05e+06u as=2.173e+11p ps=2.17e+06u
M1001 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=6.168e+11p pd=4.65e+06u as=1.134e+11p ps=1.38e+06u
M1002 VGND a_244_47# a_355_47# VNB nshort w=650000u l=250000u
+  ad=0p pd=0u as=1.7225e+11p ps=1.83e+06u
M1003 X a_355_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=4.95e+11p pd=2.99e+06u as=0p ps=0u
M1004 VPWR A a_27_47# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1005 a_244_47# a_27_47# VGND VNB nshort w=650000u l=250000u
+  ad=1.7225e+11p pd=1.83e+06u as=0p ps=0u
M1006 X a_355_47# VGND VNB nshort w=420000u l=150000u
+  ad=2.079e+11p pd=1.83e+06u as=0p ps=0u
M1007 a_244_47# a_27_47# VPWR VPB phighvt w=820000u l=250000u
+  ad=2.173e+11p pd=2.17e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__o22a_2.spice.pex
* Created: Thu Aug 27 14:37:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O22A_2%A_81_21# 1 2 7 9 12 14 16 19 24 25 27 28 29
+ 30 32 35 36
c80 35 0 8.67224e-20 $X=2.05 $Y=0.73
c81 24 0 1.48555e-19 $X=1.135 $Y=1.16
r82 43 44 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.9 $Y=1.16 $X2=0.91
+ $Y2=1.16
r83 42 43 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.49 $Y=1.16 $X2=0.9
+ $Y2=1.16
r84 40 42 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.48 $Y=1.16 $X2=0.49
+ $Y2=1.16
r85 35 36 10.1417 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=2.05 $Y=0.77 $X2=1.85
+ $Y2=0.77
r86 30 39 2.69144 $w=3.85e-07 $l=1.05e-07 $layer=LI1_cond $X=2.382 $Y=1.705
+ $X2=2.382 $Y2=1.6
r87 30 32 17.8105 $w=3.83e-07 $l=5.95e-07 $layer=LI1_cond $X=2.382 $Y=1.705
+ $X2=2.382 $Y2=2.3
r88 28 39 4.92149 $w=2.1e-07 $l=1.92e-07 $layer=LI1_cond $X=2.19 $Y=1.6
+ $X2=2.382 $Y2=1.6
r89 28 29 49.381 $w=2.08e-07 $l=9.35e-07 $layer=LI1_cond $X=2.19 $Y=1.6
+ $X2=1.255 $Y2=1.6
r90 27 36 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=1.255 $Y=0.805
+ $X2=1.85 $Y2=0.805
r91 25 44 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.135 $Y=1.16
+ $X2=0.91 $Y2=1.16
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.16 $X2=1.135 $Y2=1.16
r93 22 29 6.999 $w=2.1e-07 $l=1.85203e-07 $layer=LI1_cond $X=1.115 $Y=1.495
+ $X2=1.255 $Y2=1.6
r94 22 24 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.115 $Y=1.495
+ $X2=1.115 $Y2=1.16
r95 21 27 7.24404 $w=1.8e-07 $l=1.79444e-07 $layer=LI1_cond $X=1.115 $Y=0.895
+ $X2=1.255 $Y2=0.805
r96 21 24 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.115 $Y=0.895
+ $X2=1.115 $Y2=1.16
r97 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r98 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r99 14 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=1.16
r100 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.9 $Y2=0.56
r101 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r102 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.985
r103 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r104 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=0.56
r105 2 39 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.485 $X2=2.41 $Y2=1.62
r106 2 32 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.485 $X2=2.41 $Y2=2.3
r107 1 35 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.05 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%B1 1 3 6 8 14
c32 14 0 2.66047e-20 $X=1.84 $Y=1.16
c33 8 0 1.88537e-19 $X=1.605 $Y=1.19
r34 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.625 $Y=1.16
+ $X2=1.84 $Y2=1.16
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.16 $X2=1.625 $Y2=1.16
r36 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.16
r37 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.84 $Y=1.325 $X2=1.84
+ $Y2=1.985
r38 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.84 $Y=0.995 $X2=1.84
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%B2 3 5 7 8 11 12
c36 11 0 3.01914e-19 $X=2.26 $Y=1.16
r37 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.26 $Y2=1.325
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r39 8 12 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=2.065 $Y=1.2
+ $X2=2.26 $Y2=1.2
r40 5 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.995
+ $X2=2.26 $Y2=1.16
r41 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.26 $Y=0.995 $X2=2.26
+ $Y2=0.56
r42 3 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.2 $Y=1.985 $X2=2.2
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%A2 3 6 8 11 12 15
c39 15 0 8.67224e-20 $X=2.75 $Y=0.995
c40 11 0 4.78532e-20 $X=2.76 $Y=1.16
c41 8 0 2.66047e-20 $X=3 $Y=1.615
r42 11 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=1.325
r43 11 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.16
+ $X2=2.75 $Y2=0.995
r44 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.16 $X2=2.76 $Y2=1.16
r45 8 12 15.555 $w=2e-07 $l=2.55e-07 $layer=LI1_cond $X=3 $Y=1.615 $X2=3
+ $Y2=1.87
r46 8 10 19.6881 $w=3.04e-07 $l=5.25966e-07 $layer=LI1_cond $X=3 $Y=1.615
+ $X2=2.847 $Y2=1.16
r47 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.82 $Y=1.985
+ $X2=2.82 $Y2=1.325
r48 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.79 $Y=0.56 $X2=2.79
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%A1 3 7 8 9 14 16 27
c29 9 0 4.78532e-20 $X=3.36 $Y=1.445
r30 14 17 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.16
+ $X2=3.275 $Y2=1.325
r31 14 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.16
+ $X2=3.275 $Y2=0.995
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.16 $X2=3.29 $Y2=1.16
r33 8 27 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.445 $Y=1.175
+ $X2=3.45 $Y2=1.175
r34 8 15 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=3.43 $Y=1.175
+ $X2=3.29 $Y2=1.175
r35 8 9 7.66305 $w=4.88e-07 $l=2.55e-07 $layer=LI1_cond $X=3.43 $Y=1.275
+ $X2=3.43 $Y2=1.53
r36 7 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.56 $X2=3.21
+ $Y2=0.995
r37 3 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.18 $Y=1.985
+ $X2=3.18 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%VPWR 1 2 3 10 12 16 18 20 22 27 39 47 51
c47 2 0 1.48555e-19 $X=0.985 $Y=1.485
r48 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r49 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 39 42 11.3627 $w=7.98e-07 $l=7.6e-07 $layer=LI1_cond $X=1.395 $Y=1.96
+ $X2=1.395 $Y2=2.72
r51 36 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 31 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 30 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 28 42 10.2089 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=1.795 $Y=2.72 $X2=1.395
+ $Y2=2.72
r59 28 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 27 46 4.70099 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=3.475 $Y2=2.72
r61 27 33 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 26 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 26 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 23 36 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r66 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 22 42 10.2089 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=0.995 $Y=2.72 $X2=1.395
+ $Y2=2.72
r68 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 20 51 0.00426813 $w=4.8e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 16 46 2.98112 $w=3.2e-07 $l=1.05119e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.475 $Y2=2.72
r71 16 18 24.3093 $w=3.18e-07 $l=6.75e-07 $layer=LI1_cond $X=3.43 $Y=2.635
+ $X2=3.43 $Y2=1.96
r72 12 15 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.24 $Y2=2.3
r73 10 36 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.182 $Y2=2.72
r74 10 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.3
r75 3 18 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=1.485 $X2=3.39 $Y2=1.96
r76 2 39 150 $w=1.7e-07 $l=8.49941e-07 $layer=licon1_PDIFF $count=4 $X=0.985
+ $Y=1.485 $X2=1.63 $Y2=1.96
r77 1 15 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r78 1 12 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%X 1 2 7 10
r16 10 13 54.9421 $w=2.13e-07 $l=1.025e-06 $layer=LI1_cond $X=0.697 $Y=0.595
+ $X2=0.697 $Y2=1.62
r17 7 17 4.82418 $w=2.13e-07 $l=9e-08 $layer=LI1_cond $X=0.697 $Y=2.21 $X2=0.697
+ $Y2=2.3
r18 7 13 31.6252 $w=2.13e-07 $l=5.9e-07 $layer=LI1_cond $X=0.697 $Y=2.21
+ $X2=0.697 $Y2=1.62
r19 2 17 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.3
r20 2 13 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.62
r21 1 10 182 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.69 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%VGND 1 2 3 10 12 16 18 22 24 26 33 34 40 43
+ 48
r54 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 41 44 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r56 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r57 37 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 34 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r59 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r60 31 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0 $X2=3
+ $Y2=0
r61 31 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.45
+ $Y2=0
r62 30 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r63 30 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r64 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 27 37 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r66 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r67 26 40 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.115
+ $Y2=0
r68 26 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.69
+ $Y2=0
r69 24 48 0.00426813 $w=4.8e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=0
+ $X2=0.23 $Y2=0
r70 20 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0
r71 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0.36
r72 19 40 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.115
+ $Y2=0
r73 18 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0 $X2=3
+ $Y2=0
r74 18 19 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=1.205 $Y2=0
r75 14 40 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r76 14 16 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.38
r77 10 37 3.40825 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.177 $Y2=0
r78 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r79 3 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3 $Y2=0.36
r80 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=1.11 $Y2=0.38
r81 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O22A_2%A_301_47# 1 2 3 10 14 15 16 20
c41 15 0 1.13378e-19 $X=2.56 $Y=0.695
r42 18 20 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=3.422 $Y=0.695
+ $X2=3.422 $Y2=0.39
r43 17 25 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.73 $Y=0.78 $X2=2.56
+ $Y2=0.78
r44 16 18 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=3.422 $Y2=0.695
r45 16 17 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.255 $Y=0.78
+ $X2=2.73 $Y2=0.78
r46 15 25 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.695
+ $X2=2.56 $Y2=0.78
r47 14 23 2.66241 $w=3.4e-07 $l=9e-08 $layer=LI1_cond $X=2.56 $Y=0.475 $X2=2.56
+ $Y2=0.385
r48 14 15 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=2.56 $Y=0.475
+ $X2=2.56 $Y2=0.695
r49 10 23 5.02899 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.39 $Y=0.385
+ $X2=2.56 $Y2=0.385
r50 10 12 46.8283 $w=1.78e-07 $l=7.6e-07 $layer=LI1_cond $X=2.39 $Y=0.385
+ $X2=1.63 $Y2=0.385
r51 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.39
r52 2 25 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.555 $Y2=0.73
r53 2 23 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.555 $Y2=0.39
r54 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.63 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__nand3b_1.spice.SKY130_FD_SC_HD__NAND3B_1.pxi
* Created: Thu Aug 27 14:29:46 2020
* 
x_PM_SKY130_FD_SC_HD__NAND3B_1%A_N N_A_N_M1004_g N_A_N_M1003_g A_N N_A_N_c_49_n
+ N_A_N_c_50_n PM_SKY130_FD_SC_HD__NAND3B_1%A_N
x_PM_SKY130_FD_SC_HD__NAND3B_1%C N_C_M1002_g N_C_M1007_g C N_C_c_79_n N_C_c_80_n
+ PM_SKY130_FD_SC_HD__NAND3B_1%C
x_PM_SKY130_FD_SC_HD__NAND3B_1%B N_B_M1000_g N_B_M1001_g B N_B_c_110_n
+ N_B_c_111_n PM_SKY130_FD_SC_HD__NAND3B_1%B
x_PM_SKY130_FD_SC_HD__NAND3B_1%A_53_93# N_A_53_93#_M1004_s N_A_53_93#_M1003_s
+ N_A_53_93#_M1006_g N_A_53_93#_M1005_g N_A_53_93#_c_145_n N_A_53_93#_c_159_n
+ N_A_53_93#_c_146_n N_A_53_93#_c_147_n N_A_53_93#_c_148_n N_A_53_93#_c_154_n
+ N_A_53_93#_c_149_n PM_SKY130_FD_SC_HD__NAND3B_1%A_53_93#
x_PM_SKY130_FD_SC_HD__NAND3B_1%VPWR N_VPWR_M1003_d N_VPWR_M1001_d N_VPWR_c_217_n
+ N_VPWR_c_218_n N_VPWR_c_219_n N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n
+ VPWR N_VPWR_c_223_n N_VPWR_c_216_n PM_SKY130_FD_SC_HD__NAND3B_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND3B_1%Y N_Y_M1006_d N_Y_M1007_d N_Y_M1005_d N_Y_c_255_n
+ N_Y_c_257_n N_Y_c_261_n N_Y_c_264_n Y Y Y Y Y Y N_Y_c_250_n Y
+ PM_SKY130_FD_SC_HD__NAND3B_1%Y
x_PM_SKY130_FD_SC_HD__NAND3B_1%VGND N_VGND_M1004_d N_VGND_c_298_n N_VGND_c_299_n
+ N_VGND_c_300_n VGND N_VGND_c_301_n N_VGND_c_302_n
+ PM_SKY130_FD_SC_HD__NAND3B_1%VGND
cc_1 VNB A_N 0.00282198f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_2 VNB N_A_N_c_49_n 0.02557f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_3 VNB N_A_N_c_50_n 0.0211638f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_4 VNB C 0.00213592f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_5 VNB N_C_c_79_n 0.0234632f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_6 VNB N_C_c_80_n 0.0185094f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_7 VNB B 0.00161387f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.105
cc_8 VNB N_B_c_110_n 0.0261171f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_9 VNB N_B_c_111_n 0.017476f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_10 VNB N_A_53_93#_c_145_n 0.023339f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_11 VNB N_A_53_93#_c_146_n 0.00101052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_53_93#_c_147_n 0.0285487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_53_93#_c_148_n 0.0228497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_53_93#_c_149_n 0.0211747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_216_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Y_c_250_n 0.0135475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.0410378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_298_n 0.00795355f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.695
cc_19 VNB N_VGND_c_299_n 0.0211377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_300_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_21 VNB N_VGND_c_301_n 0.0457124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_302_n 0.169053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VPB N_A_N_M1003_g 0.0253918f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_24 VPB A_N 0.0020516f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_25 VPB N_A_N_c_49_n 0.00638382f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_26 VPB N_C_M1007_g 0.0221988f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_27 VPB C 3.0539e-19 $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_28 VPB N_C_c_79_n 0.00692673f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_29 VPB N_B_M1001_g 0.0203709f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.695
cc_30 VPB B 0.00161387f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_31 VPB N_B_c_110_n 0.00632297f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_32 VPB N_A_53_93#_M1005_g 0.0238175f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_33 VPB N_A_53_93#_c_145_n 0.0149536f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_34 VPB N_A_53_93#_c_146_n 9.27585e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_53_93#_c_147_n 0.00628489f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_53_93#_c_154_n 0.0236179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_217_n 0.022704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_218_n 0.00474998f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_39 VPB N_VPWR_c_219_n 0.0247369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_220_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_221_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_222_n 0.00544936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_223_n 0.0233753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_216_n 0.0554244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB Y 0.00868423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB Y 0.0422471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB Y 0.0107819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 N_A_N_M1003_g N_C_M1007_g 0.0143222f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_49 A_N C 0.0238604f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_N_c_49_n C 3.00886e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_51 A_N N_C_c_79_n 0.00219735f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_52 N_A_N_c_49_n N_C_c_79_n 0.0204854f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_N_c_50_n N_C_c_80_n 0.0203883f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_N_M1003_g N_A_53_93#_c_145_n 0.0067114f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_55 A_N N_A_53_93#_c_145_n 0.0248817f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_N_c_49_n N_A_53_93#_c_145_n 0.00816168f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_N_c_50_n N_A_53_93#_c_145_n 0.00521379f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A_N_c_50_n N_A_53_93#_c_159_n 0.0102212f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_59 A_N N_A_53_93#_c_148_n 0.0219504f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_60 N_A_N_c_49_n N_A_53_93#_c_148_n 0.00542336f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_N_c_50_n N_A_53_93#_c_148_n 4.58643e-19 $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_N_M1003_g N_A_53_93#_c_154_n 4.58643e-19 $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_63 A_N N_A_53_93#_c_154_n 0.00343051f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_N_c_49_n N_A_53_93#_c_154_n 0.00458826f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_N_M1003_g N_VPWR_c_217_n 0.0052717f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_66 A_N N_VPWR_c_217_n 0.00460569f $X=0.605 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_N_M1003_g N_VPWR_c_219_n 0.00327927f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_68 N_A_N_M1003_g N_VPWR_c_216_n 0.00417489f $X=0.6 $Y=1.695 $X2=0 $Y2=0
cc_69 N_A_N_c_50_n N_VGND_c_298_n 0.00343738f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_N_c_50_n N_VGND_c_299_n 0.00393318f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_N_c_50_n N_VGND_c_302_n 0.00512902f $X=0.51 $Y=0.995 $X2=0 $Y2=0
cc_72 N_C_M1007_g N_B_M1001_g 0.0151563f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_73 C B 0.0236096f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_74 N_C_c_79_n B 3.96006e-19 $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_75 C N_B_c_110_n 0.00182429f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_76 N_C_c_79_n N_B_c_110_n 0.0207134f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_c_80_n N_B_c_111_n 0.0444797f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_78 C N_A_53_93#_c_159_n 0.0159505f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_79 N_C_c_79_n N_A_53_93#_c_159_n 0.00301183f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_80 N_C_c_80_n N_A_53_93#_c_159_n 0.0117968f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_81 N_C_M1007_g N_VPWR_c_217_n 0.00321269f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_82 N_C_c_79_n N_VPWR_c_217_n 0.00217348f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_M1007_g N_VPWR_c_221_n 0.00541359f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_84 N_C_M1007_g N_VPWR_c_216_n 0.0108548f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_85 N_C_M1007_g N_Y_c_255_n 0.0022193f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_86 C N_Y_c_255_n 0.0060702f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_87 N_C_M1007_g N_Y_c_257_n 0.00885586f $X=1.085 $Y=1.985 $X2=0 $Y2=0
cc_88 N_C_c_80_n N_VGND_c_298_n 0.0110169f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_89 N_C_c_80_n N_VGND_c_301_n 0.00341689f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C_c_80_n N_VGND_c_302_n 0.00405445f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B_M1001_g N_A_53_93#_M1005_g 0.0198628f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_92 B N_A_53_93#_c_159_n 0.0217525f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B_c_110_n N_A_53_93#_c_159_n 0.00110224f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B_c_111_n N_A_53_93#_c_159_n 0.0123433f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_95 B N_A_53_93#_c_146_n 0.0153762f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B_c_110_n N_A_53_93#_c_146_n 0.00102339f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_c_111_n N_A_53_93#_c_146_n 8.52962e-19 $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_98 B N_A_53_93#_c_147_n 0.00122018f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B_c_110_n N_A_53_93#_c_147_n 0.0204065f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B_c_111_n N_A_53_93#_c_149_n 0.0298473f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B_M1001_g N_VPWR_c_218_n 0.0016963f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B_M1001_g N_VPWR_c_221_n 0.00541359f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B_M1001_g N_VPWR_c_216_n 0.00981263f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B_M1001_g N_Y_c_255_n 8.8334e-19 $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_105 B N_Y_c_255_n 0.00251657f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_106 N_B_M1001_g N_Y_c_257_n 0.010277f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B_M1001_g N_Y_c_261_n 0.0112741f $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_108 B N_Y_c_261_n 0.0194139f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B_c_110_n N_Y_c_261_n 0.00110224f $X=1.59 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B_c_111_n N_Y_c_264_n 0.00106258f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_M1001_g Y 5.92331e-19 $X=1.505 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B_c_111_n N_VGND_c_298_n 0.00227626f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_111_n N_VGND_c_301_n 0.00428022f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B_c_111_n N_VGND_c_302_n 0.00624857f $X=1.59 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_53_93#_c_159_n N_VPWR_c_217_n 0.00511975f $X=2.045 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_53_93#_c_154_n N_VPWR_c_217_n 0.00133957f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_117 N_A_53_93#_M1005_g N_VPWR_c_218_n 0.00299999f $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_118 N_A_53_93#_M1005_g N_VPWR_c_223_n 0.00541359f $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_53_93#_M1005_g N_VPWR_c_216_n 0.0109082f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_53_93#_c_154_n N_VPWR_c_216_n 0.0161088f $X=0.39 $Y=1.76 $X2=0 $Y2=0
cc_121 N_A_53_93#_c_159_n N_Y_M1006_d 0.00233548f $X=2.045 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_53_93#_c_146_n N_Y_M1006_d 6.2871e-19 $X=2.13 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_53_93#_c_159_n N_Y_c_255_n 0.00398354f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_53_93#_M1005_g N_Y_c_257_n 5.96051e-19 $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_53_93#_M1005_g N_Y_c_261_n 0.012479f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_53_93#_c_159_n N_Y_c_261_n 0.00569346f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_53_93#_c_146_n N_Y_c_261_n 0.00293308f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_53_93#_c_159_n N_Y_c_264_n 0.00556146f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_53_93#_c_147_n N_Y_c_264_n 0.00246454f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_53_93#_c_149_n N_Y_c_264_n 0.00555535f $X=2.13 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_53_93#_M1005_g Y 8.8334e-19 $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_53_93#_c_146_n Y 0.00856844f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_53_93#_c_147_n Y 0.00421057f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_53_93#_M1005_g Y 0.010277f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_53_93#_M1005_g Y 0.00539085f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_53_93#_c_159_n Y 0.0143469f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_53_93#_c_146_n Y 0.0377835f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_53_93#_c_147_n Y 0.00824505f $X=2.13 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_53_93#_c_149_n Y 0.0061565f $X=2.13 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_53_93#_c_159_n N_VGND_M1004_d 0.00605005f $X=2.045 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_53_93#_c_159_n N_VGND_c_298_n 0.0190084f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A_53_93#_c_148_n N_VGND_c_298_n 0.00136717f $X=0.51 $Y=0.635 $X2=0
+ $Y2=0
cc_143 N_A_53_93#_c_159_n N_VGND_c_299_n 0.00279278f $X=2.045 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_53_93#_c_148_n N_VGND_c_299_n 0.01312f $X=0.51 $Y=0.635 $X2=0 $Y2=0
cc_145 N_A_53_93#_c_159_n N_VGND_c_301_n 0.0154117f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_53_93#_c_149_n N_VGND_c_301_n 0.00413954f $X=2.13 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_53_93#_c_159_n N_VGND_c_302_n 0.0344387f $X=2.045 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_53_93#_c_148_n N_VGND_c_302_n 0.0143027f $X=0.51 $Y=0.635 $X2=0 $Y2=0
cc_149 N_A_53_93#_c_149_n N_VGND_c_302_n 0.00717131f $X=2.13 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_53_93#_c_159_n A_232_47# 0.00588528f $X=2.045 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_53_93#_c_159_n A_316_47# 0.0092823f $X=2.045 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_152 N_VPWR_c_216_n N_Y_M1007_d 0.00215201f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_153 N_VPWR_c_216_n N_Y_M1005_d 0.00225715f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_221_n N_Y_c_257_n 0.0189039f $X=1.63 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_216_n N_Y_c_257_n 0.0122217f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_M1001_d N_Y_c_261_n 0.00732793f $X=1.58 $Y=1.485 $X2=0 $Y2=0
cc_157 N_VPWR_c_218_n N_Y_c_261_n 0.0220482f $X=1.775 $Y=2 $X2=0 $Y2=0
cc_158 N_VPWR_c_223_n Y 0.0396514f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_c_216_n Y 0.0224398f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_160 N_Y_c_264_n N_VGND_c_301_n 0.0176166f $X=2.385 $Y=0.37 $X2=0 $Y2=0
cc_161 N_Y_c_250_n N_VGND_c_301_n 0.0207779f $X=2.53 $Y=0.485 $X2=0 $Y2=0
cc_162 N_Y_M1006_d N_VGND_c_302_n 0.00225741f $X=2.115 $Y=0.235 $X2=0 $Y2=0
cc_163 N_Y_c_264_n N_VGND_c_302_n 0.0110356f $X=2.385 $Y=0.37 $X2=0 $Y2=0
cc_164 N_Y_c_250_n N_VGND_c_302_n 0.0111684f $X=2.53 $Y=0.485 $X2=0 $Y2=0
cc_165 N_VGND_c_302_n A_232_47# 0.00323135f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_166 N_VGND_c_302_n A_316_47# 0.00460767f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 a_1031_413# a_27_47# a_938_413# VPB phighvt w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.323e+11p ps=1.47e+06u
M1001 a_1097_183# a_938_413# VGND VNB nshort w=640000u l=150000u
+  ad=1.978e+11p pd=1.99e+06u as=1.5361e+12p ps=1.571e+07u
M1002 VPWR a_2049_47# Q_N VPB phighvt w=1e+06u l=150000u
+  ad=2.17125e+12p pd=1.991e+07u as=2.7e+11p ps=2.54e+06u
M1003 VGND a_1525_315# a_1483_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1004 VPWR SCD a_644_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.016e+11p ps=1.91e+06u
M1005 VPWR a_1525_315# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VGND a_2049_47# Q_N VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1007 a_644_369# a_299_47# a_560_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.841e+11p ps=3.19e+06u
M1008 a_1438_413# a_193_47# a_1354_413# VPB phighvt w=420000u l=150000u
+  ad=1.827e+11p pd=1.71e+06u as=1.134e+11p ps=1.38e+06u
M1009 Q_N a_2049_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_560_369# D a_466_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1011 VGND SCD a_661_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1012 VPWR CLK a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1013 VPWR a_1097_183# a_1031_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Q_N a_2049_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_938_413# a_193_47# a_560_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_487_47# a_299_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1017 a_560_369# D a_487_47# VNB nshort w=420000u l=150000u
+  ad=2.394e+11p pd=2.78e+06u as=0p ps=0u
M1018 a_1354_413# a_27_47# a_1097_183# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.19e+11p ps=2.15e+06u
M1019 Q a_1525_315# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1035_47# a_193_47# a_938_413# VNB nshort w=360000u l=150000u
+  ad=1.374e+11p pd=1.52e+06u as=1.188e+11p ps=1.38e+06u
M1021 a_661_47# SCE a_560_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1354_413# a_193_47# a_1097_183# VNB nshort w=360000u l=150000u
+  ad=1.314e+11p pd=1.45e+06u as=0p ps=0u
M1023 a_1483_47# a_27_47# a_1354_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_938_413# a_27_47# a_560_369# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_1525_315# a_2049_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1026 a_466_369# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1028 VGND a_1525_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1029 Q a_1525_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR SCE a_299_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1031 VPWR a_1525_315# a_1438_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_1354_413# a_1525_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1033 a_1097_183# a_938_413# VPWR VPB phighvt w=750000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_1097_183# a_1035_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_1354_413# a_1525_315# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
M1036 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=0p ps=0u
M1037 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1038 VPWR a_1525_315# a_2049_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1039 VGND SCE a_299_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
.ends

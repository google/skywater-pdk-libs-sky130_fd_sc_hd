* File: sky130_fd_sc_hd__nand4bb_2.pxi.spice
* Created: Thu Aug 27 14:30:56 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4BB_2%B_N N_B_N_c_116_n N_B_N_c_111_n N_B_N_M1017_g
+ N_B_N_M1004_g N_B_N_c_112_n N_B_N_c_118_n B_N B_N N_B_N_c_114_n N_B_N_c_115_n
+ PM_SKY130_FD_SC_HD__NAND4BB_2%B_N
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_N N_A_N_M1006_g N_A_N_M1019_g A_N A_N
+ N_A_N_c_153_n PM_SKY130_FD_SC_HD__NAND4BB_2%A_N
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_193_47# N_A_193_47#_M1006_d
+ N_A_193_47#_M1019_d N_A_193_47#_c_189_n N_A_193_47#_M1009_g
+ N_A_193_47#_M1005_g N_A_193_47#_c_190_n N_A_193_47#_M1015_g
+ N_A_193_47#_M1008_g N_A_193_47#_c_193_n N_A_193_47#_c_194_n
+ N_A_193_47#_c_202_n N_A_193_47#_c_195_n N_A_193_47#_c_196_n
+ N_A_193_47#_c_203_n N_A_193_47#_c_197_n N_A_193_47#_c_204_n
+ PM_SKY130_FD_SC_HD__NAND4BB_2%A_193_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_27_47# N_A_27_47#_M1017_s N_A_27_47#_M1004_s
+ N_A_27_47#_M1014_g N_A_27_47#_M1000_g N_A_27_47#_M1018_g N_A_27_47#_M1001_g
+ N_A_27_47#_c_272_n N_A_27_47#_c_281_n N_A_27_47#_c_273_n N_A_27_47#_c_274_n
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_c_275_n N_A_27_47#_c_276_n
+ N_A_27_47#_c_277_n N_A_27_47#_c_278_n PM_SKY130_FD_SC_HD__NAND4BB_2%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_2%C N_C_M1010_g N_C_M1011_g N_C_M1016_g
+ N_C_M1013_g C C N_C_c_386_n N_C_c_387_n PM_SKY130_FD_SC_HD__NAND4BB_2%C
x_PM_SKY130_FD_SC_HD__NAND4BB_2%D N_D_M1003_g N_D_M1002_g N_D_M1007_g
+ N_D_M1012_g N_D_c_432_n D D N_D_c_434_n PM_SKY130_FD_SC_HD__NAND4BB_2%D
x_PM_SKY130_FD_SC_HD__NAND4BB_2%VPWR N_VPWR_M1004_d N_VPWR_M1005_d
+ N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1013_d N_VPWR_M1012_s N_VPWR_c_481_n
+ N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_492_n VPWR N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_480_n
+ PM_SKY130_FD_SC_HD__NAND4BB_2%VPWR
x_PM_SKY130_FD_SC_HD__NAND4BB_2%Y N_Y_M1009_d N_Y_M1005_s N_Y_M1000_s
+ N_Y_M1011_s N_Y_M1002_d N_Y_c_576_n N_Y_c_584_n N_Y_c_569_n N_Y_c_586_n
+ N_Y_c_570_n N_Y_c_571_n N_Y_c_612_n N_Y_c_572_n N_Y_c_573_n N_Y_c_615_n
+ N_Y_c_587_n N_Y_c_574_n Y Y PM_SKY130_FD_SC_HD__NAND4BB_2%Y
x_PM_SKY130_FD_SC_HD__NAND4BB_2%VGND N_VGND_M1017_d N_VGND_M1003_s
+ N_VGND_c_660_n N_VGND_c_661_n VGND N_VGND_c_662_n N_VGND_c_663_n
+ N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ PM_SKY130_FD_SC_HD__NAND4BB_2%VGND
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_341_47# N_A_341_47#_M1009_s
+ N_A_341_47#_M1015_s N_A_341_47#_M1018_s N_A_341_47#_c_728_n
+ N_A_341_47#_c_732_n PM_SKY130_FD_SC_HD__NAND4BB_2%A_341_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_591_47# N_A_591_47#_M1014_d
+ N_A_591_47#_M1010_d N_A_591_47#_c_752_n
+ PM_SKY130_FD_SC_HD__NAND4BB_2%A_591_47#
x_PM_SKY130_FD_SC_HD__NAND4BB_2%A_781_47# N_A_781_47#_M1010_s
+ N_A_781_47#_M1016_s N_A_781_47#_M1007_d N_A_781_47#_c_778_n
+ N_A_781_47#_c_784_n N_A_781_47#_c_779_n N_A_781_47#_c_780_n
+ N_A_781_47#_c_781_n PM_SKY130_FD_SC_HD__NAND4BB_2%A_781_47#
cc_1 VNB N_B_N_c_111_n 0.017179f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_2 VNB N_B_N_c_112_n 0.0209321f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_3 VNB B_N 0.00978855f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_B_N_c_114_n 0.0211912f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_B_N_c_115_n 0.0159684f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_N_M1006_g 0.0394842f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_7 VNB A_N 0.00329807f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_8 VNB N_A_N_c_153_n 0.022609f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_9 VNB N_A_193_47#_c_189_n 0.019205f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_10 VNB N_A_193_47#_c_190_n 0.0258549f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_11 VNB N_A_193_47#_M1015_g 0.017202f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.86
cc_12 VNB N_A_193_47#_M1008_g 3.79881e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB N_A_193_47#_c_193_n 0.047002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_193_47#_c_194_n 0.00468706f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_15 VNB N_A_193_47#_c_195_n 0.00219447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_193_47#_c_196_n 0.00326686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_193_47#_c_197_n 0.00315598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1014_g 0.017695f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_19 VNB N_A_27_47#_M1000_g 3.81135e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_M1018_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_M1001_g 5.54454e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_22 VNB N_A_27_47#_c_272_n 0.0187453f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_23 VNB N_A_27_47#_c_273_n 0.0167625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_274_n 0.00786701f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_25 VNB N_A_27_47#_c_275_n 0.00625044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_276_n 0.00614679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_277_n 0.0011775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_278_n 0.0356874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_C_M1010_g 0.0238956f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_30 VNB N_C_M1011_g 5.70974e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_31 VNB N_C_M1016_g 0.0176998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_C_M1013_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB C 0.00338482f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_34 VNB N_C_c_386_n 0.0304245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_C_c_387_n 0.0251087f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_36 VNB N_D_M1003_g 0.017551f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.4
cc_37 VNB N_D_M1002_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_38 VNB N_D_M1007_g 0.0230765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_D_c_432_n 0.0289271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB D 0.00962113f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_41 VNB N_D_c_434_n 0.0268068f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_42 VNB N_VPWR_c_480_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB Y 0.00327973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_660_n 0.00231024f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_45 VNB N_VGND_c_661_n 0.00462218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_662_n 0.0144236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_663_n 0.103045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_664_n 0.017368f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.19
cc_49 VNB N_VGND_c_665_n 0.30499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_666_n 0.00353477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_667_n 0.00323621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_341_47#_c_728_n 0.00271098f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.805
cc_53 VNB N_A_591_47#_c_752_n 0.0177036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_781_47#_c_778_n 0.00263528f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_55 VNB N_A_781_47#_c_779_n 0.00295923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_781_47#_c_780_n 0.0115894f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.86
cc_57 VNB N_A_781_47#_c_781_n 0.0194553f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_58 VPB N_B_N_c_116_n 0.0293096f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.785
cc_59 VPB N_B_N_M1004_g 0.0203205f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_60 VPB N_B_N_c_118_n 0.0248783f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.86
cc_61 VPB B_N 0.0124835f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_62 VPB N_B_N_c_114_n 0.0106323f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_63 VPB N_A_N_M1019_g 0.051109f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_64 VPB A_N 0.00399757f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_65 VPB N_A_N_c_153_n 0.0153927f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_66 VPB N_A_193_47#_M1005_g 0.0219362f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.805
cc_67 VPB N_A_193_47#_c_190_n 5.75634e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.805
cc_68 VPB N_A_193_47#_M1008_g 0.0186154f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_69 VPB N_A_193_47#_c_193_n 0.0240707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_193_47#_c_202_n 0.00481164f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_71 VPB N_A_193_47#_c_203_n 0.0142533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_193_47#_c_204_n 0.00144621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_M1000_g 0.0194255f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_M1001_g 0.0240955f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_75 VPB N_A_27_47#_c_281_n 0.0185621f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_76 VPB N_A_27_47#_c_282_n 0.0124615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_283_n 0.00897929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_275_n 0.00996251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_276_n 0.00865004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_C_M1011_g 0.0243476f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_81 VPB N_C_M1013_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_D_M1002_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_83 VPB N_D_M1012_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_D_c_434_n 0.00835978f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_85 VPB N_VPWR_c_481_n 0.00230843f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_86 VPB N_VPWR_c_482_n 0.00407299f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_87 VPB N_VPWR_c_483_n 0.0152056f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.19
cc_88 VPB N_VPWR_c_484_n 0.00171127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_485_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_486_n 0.00645473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_487_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_488_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_489_n 0.0100765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_490_n 0.046934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_491_n 0.0243819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_492_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_493_n 0.0151232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_494_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_495_n 0.00320131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_496_n 0.00353672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_497_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_498_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_480_n 0.0501142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_Y_c_569_n 0.00260929f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_105 VPB N_Y_c_570_n 0.00611787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_Y_c_571_n 0.00307011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_Y_c_572_n 0.00455314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_Y_c_573_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_574_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB Y 0.00262866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 N_B_N_c_111_n N_A_N_M1006_g 0.0209954f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_112 N_B_N_c_115_n N_A_N_M1006_g 0.00598582f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_113 N_B_N_c_116_n N_A_N_M1019_g 0.009307f $X=0.305 $Y=1.785 $X2=0 $Y2=0
cc_114 N_B_N_c_118_n N_A_N_M1019_g 0.0244503f $X=0.47 $Y=1.86 $X2=0 $Y2=0
cc_115 N_B_N_c_116_n A_N 0.00152699f $X=0.305 $Y=1.785 $X2=0 $Y2=0
cc_116 B_N A_N 0.0297095f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_117 N_B_N_c_114_n A_N 0.00175932f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_118 B_N N_A_N_c_153_n 7.2408e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B_N_c_114_n N_A_N_c_153_n 0.0202651f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_120 N_B_N_c_111_n N_A_27_47#_c_272_n 0.00320911f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_121 N_B_N_M1004_g N_A_27_47#_c_281_n 0.00387938f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_122 N_B_N_c_112_n N_A_27_47#_c_273_n 0.011081f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_123 N_B_N_c_115_n N_A_27_47#_c_273_n 0.00185237f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_124 N_B_N_c_112_n N_A_27_47#_c_274_n 0.00675396f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_125 B_N N_A_27_47#_c_274_n 0.020875f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B_N_c_114_n N_A_27_47#_c_274_n 9.79955e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_127 N_B_N_c_115_n N_A_27_47#_c_274_n 0.00273512f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_128 N_B_N_M1004_g N_A_27_47#_c_282_n 0.00569569f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_129 N_B_N_c_118_n N_A_27_47#_c_282_n 0.0110175f $X=0.47 $Y=1.86 $X2=0 $Y2=0
cc_130 N_B_N_c_118_n N_A_27_47#_c_283_n 0.0111984f $X=0.47 $Y=1.86 $X2=0 $Y2=0
cc_131 B_N N_A_27_47#_c_283_n 0.0214513f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B_N_c_114_n N_A_27_47#_c_283_n 6.00486e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_133 N_B_N_M1004_g N_VPWR_c_481_n 0.00768947f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_134 N_B_N_M1004_g N_VPWR_c_493_n 0.00424408f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_135 N_B_N_M1004_g N_VPWR_c_480_n 0.00594309f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_136 N_B_N_c_111_n N_VGND_c_660_n 0.00885865f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_137 N_B_N_c_111_n N_VGND_c_662_n 0.00350026f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_138 N_B_N_c_112_n N_VGND_c_662_n 0.00101953f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_139 N_B_N_c_111_n N_VGND_c_665_n 0.00516659f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_140 N_B_N_c_112_n N_VGND_c_665_n 0.00128537f $X=0.47 $Y=0.805 $X2=0 $Y2=0
cc_141 N_A_N_M1006_g N_A_193_47#_c_193_n 0.0093032f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_N_M1006_g N_A_193_47#_c_194_n 0.00416584f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_N_M1019_g N_A_193_47#_c_202_n 0.00428252f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_144 N_A_N_M1006_g N_A_193_47#_c_195_n 6.64042e-19 $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_145 N_A_N_M1019_g N_A_193_47#_c_203_n 0.00498747f $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_146 N_A_N_M1006_g N_A_193_47#_c_197_n 0.00319082f $X=0.89 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_N_M1019_g N_A_193_47#_c_204_n 6.32016e-19 $X=0.89 $Y=2.275 $X2=0
+ $Y2=0
cc_148 N_A_N_M1006_g N_A_27_47#_c_273_n 0.0154571f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_149 A_N N_A_27_47#_c_273_n 0.0252677f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_150 N_A_N_c_153_n N_A_27_47#_c_273_n 0.0018241f $X=0.725 $Y=1.255 $X2=0 $Y2=0
cc_151 N_A_N_M1019_g N_A_27_47#_c_282_n 0.0165818f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_152 A_N N_A_27_47#_c_282_n 0.0247117f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_153 N_A_N_c_153_n N_A_27_47#_c_282_n 0.00132492f $X=0.725 $Y=1.255 $X2=0
+ $Y2=0
cc_154 N_A_N_M1006_g N_A_27_47#_c_275_n 0.0202073f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_155 A_N N_A_27_47#_c_275_n 0.0384297f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_156 N_A_N_M1006_g N_A_27_47#_c_276_n 0.00537474f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_157 A_N N_A_27_47#_c_276_n 0.00814713f $X=0.61 $Y=1.445 $X2=0 $Y2=0
cc_158 N_A_N_M1019_g N_VPWR_c_481_n 0.00276606f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_159 N_A_N_M1019_g N_VPWR_c_491_n 0.00423478f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_160 N_A_N_M1019_g N_VPWR_c_480_n 0.00710834f $X=0.89 $Y=2.275 $X2=0 $Y2=0
cc_161 N_A_N_M1006_g N_VGND_c_660_n 0.00279634f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_N_M1006_g N_VGND_c_663_n 0.004224f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_N_M1006_g N_VGND_c_665_n 0.00717845f $X=0.89 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_193_47#_M1015_g N_A_27_47#_M1014_g 0.026121f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_165 N_A_193_47#_M1008_g N_A_27_47#_M1000_g 0.0299407f $X=2.46 $Y=1.985 $X2=0
+ $Y2=0
cc_166 N_A_193_47#_c_194_n N_A_27_47#_c_273_n 0.020379f $X=1.4 $Y=0.407 $X2=0
+ $Y2=0
cc_167 N_A_193_47#_c_195_n N_A_27_47#_c_273_n 0.014376f $X=1.49 $Y=0.805 $X2=0
+ $Y2=0
cc_168 N_A_193_47#_c_202_n N_A_27_47#_c_282_n 0.0210067f $X=1.4 $Y=2.307 $X2=0
+ $Y2=0
cc_169 N_A_193_47#_c_203_n N_A_27_47#_c_282_n 0.0165021f $X=1.487 $Y=2.15 $X2=0
+ $Y2=0
cc_170 N_A_193_47#_c_193_n N_A_27_47#_c_275_n 0.00248958f $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_A_193_47#_c_196_n N_A_27_47#_c_275_n 0.0645263f $X=1.495 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_A_193_47#_c_190_n N_A_27_47#_c_276_n 0.0104287f $X=2.46 $Y=1.025 $X2=0
+ $Y2=0
cc_173 N_A_193_47#_M1008_g N_A_27_47#_c_276_n 0.00114597f $X=2.46 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_193_47#_c_193_n N_A_27_47#_c_276_n 0.0243211f $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_175 N_A_193_47#_c_194_n N_A_27_47#_c_276_n 0.00681895f $X=1.4 $Y=0.407 $X2=0
+ $Y2=0
cc_176 N_A_193_47#_c_196_n N_A_27_47#_c_276_n 0.031219f $X=1.495 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_193_47#_c_190_n N_A_27_47#_c_277_n 8.41987e-19 $X=2.46 $Y=1.025 $X2=0
+ $Y2=0
cc_178 N_A_193_47#_c_190_n N_A_27_47#_c_278_n 0.0190966f $X=2.46 $Y=1.025 $X2=0
+ $Y2=0
cc_179 N_A_193_47#_M1005_g N_VPWR_c_482_n 0.0030732f $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_193_47#_c_193_n N_VPWR_c_482_n 0.00732098f $X=1.965 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_193_47#_c_202_n N_VPWR_c_482_n 0.0260524f $X=1.4 $Y=2.307 $X2=0 $Y2=0
cc_182 N_A_193_47#_c_203_n N_VPWR_c_482_n 0.0485182f $X=1.487 $Y=2.15 $X2=0
+ $Y2=0
cc_183 N_A_193_47#_M1005_g N_VPWR_c_483_n 0.00541359f $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_193_47#_M1008_g N_VPWR_c_483_n 0.0046653f $X=2.46 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_193_47#_M1005_g N_VPWR_c_484_n 7.17238e-19 $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_193_47#_M1008_g N_VPWR_c_484_n 0.0108434f $X=2.46 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_193_47#_c_202_n N_VPWR_c_491_n 0.0413283f $X=1.4 $Y=2.307 $X2=0 $Y2=0
cc_188 N_A_193_47#_M1019_d N_VPWR_c_480_n 0.00381519f $X=0.965 $Y=2.065 $X2=0
+ $Y2=0
cc_189 N_A_193_47#_M1005_g N_VPWR_c_480_n 0.0108276f $X=2.04 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_193_47#_M1008_g N_VPWR_c_480_n 0.00789179f $X=2.46 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_193_47#_c_202_n N_VPWR_c_480_n 0.0240801f $X=1.4 $Y=2.307 $X2=0 $Y2=0
cc_192 N_A_193_47#_c_189_n N_Y_c_576_n 0.00820509f $X=2.04 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_193_47#_M1005_g N_Y_c_576_n 0.00365567f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_193_47#_c_190_n N_Y_c_576_n 0.0225417f $X=2.46 $Y=1.025 $X2=0 $Y2=0
cc_195 N_A_193_47#_M1015_g N_Y_c_576_n 0.00854614f $X=2.46 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A_193_47#_M1008_g N_Y_c_576_n 0.00449457f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_197 N_A_193_47#_c_195_n N_Y_c_576_n 0.0185319f $X=1.49 $Y=0.805 $X2=0 $Y2=0
cc_198 N_A_193_47#_c_203_n N_Y_c_576_n 0.00111996f $X=1.487 $Y=2.15 $X2=0 $Y2=0
cc_199 N_A_193_47#_c_197_n N_Y_c_576_n 0.00195876f $X=1.49 $Y=0.715 $X2=0 $Y2=0
cc_200 N_A_193_47#_M1005_g N_Y_c_584_n 0.0101262f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_193_47#_M1008_g N_Y_c_569_n 0.0112739f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_193_47#_M1008_g N_Y_c_586_n 4.51827e-19 $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_193_47#_M1005_g N_Y_c_587_n 0.00454f $X=2.04 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_193_47#_M1008_g N_Y_c_587_n 0.00374603f $X=2.46 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_193_47#_c_203_n N_Y_c_587_n 0.00173948f $X=1.487 $Y=2.15 $X2=0 $Y2=0
cc_206 N_A_193_47#_c_189_n N_VGND_c_663_n 0.00357877f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_193_47#_M1015_g N_VGND_c_663_n 0.00357877f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_193_47#_c_194_n N_VGND_c_663_n 0.0413319f $X=1.4 $Y=0.407 $X2=0 $Y2=0
cc_209 N_A_193_47#_M1006_d N_VGND_c_665_n 0.00382322f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_210 N_A_193_47#_c_189_n N_VGND_c_665_n 0.00655123f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_193_47#_M1015_g N_VGND_c_665_n 0.00525237f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_212 N_A_193_47#_c_194_n N_VGND_c_665_n 0.0241431f $X=1.4 $Y=0.407 $X2=0 $Y2=0
cc_213 N_A_193_47#_c_189_n N_A_341_47#_c_728_n 0.010498f $X=2.04 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_193_47#_c_190_n N_A_341_47#_c_728_n 2.99382e-19 $X=2.46 $Y=1.025
+ $X2=0 $Y2=0
cc_215 N_A_193_47#_M1015_g N_A_341_47#_c_728_n 0.0104381f $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_216 N_A_193_47#_c_193_n N_A_341_47#_c_732_n 0.00522193f $X=1.965 $Y=1.16
+ $X2=0 $Y2=0
cc_217 N_A_193_47#_c_194_n N_A_341_47#_c_732_n 0.0271886f $X=1.4 $Y=0.407 $X2=0
+ $Y2=0
cc_218 N_A_193_47#_c_197_n N_A_341_47#_c_732_n 0.00175035f $X=1.49 $Y=0.715
+ $X2=0 $Y2=0
cc_219 N_A_193_47#_M1015_g N_A_591_47#_c_752_n 7.25252e-19 $X=2.46 $Y=0.56 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_278_n C 5.91111e-19 $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_278_n N_C_c_386_n 0.00700334f $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_282_n N_VPWR_c_481_n 0.0122859f $X=1.06 $Y=1.882 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_276_n N_VPWR_c_482_n 0.00840714f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1000_g N_VPWR_c_484_n 0.00151363f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_M1000_g N_VPWR_c_485_n 0.00541359f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_M1001_g N_VPWR_c_485_n 0.00541359f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1001_g N_VPWR_c_486_n 0.0158595f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_282_n N_VPWR_c_491_n 0.00231103f $X=1.06 $Y=1.882 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_281_n N_VPWR_c_493_n 0.0162479f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_282_n N_VPWR_c_493_n 0.00225651f $X=1.06 $Y=1.882 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1004_s N_VPWR_c_480_n 0.00223307f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1000_g N_VPWR_c_480_n 0.00952874f $X=2.88 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_M1001_g N_VPWR_c_480_n 0.0109543f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_281_n N_VPWR_c_480_n 0.0107554f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_282_n N_VPWR_c_480_n 0.00871932f $X=1.06 $Y=1.882 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_M1014_g N_Y_c_576_n 0.00132575f $X=2.88 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A_27_47#_M1000_g N_Y_c_576_n 7.70335e-19 $X=2.88 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_276_n N_Y_c_576_n 0.0416332f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_277_n N_Y_c_576_n 0.00595387f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_278_n N_Y_c_576_n 8.52883e-19 $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_27_47#_M1000_g N_Y_c_569_n 0.0119079f $X=2.88 $Y=1.985 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_276_n N_Y_c_569_n 0.0265173f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_277_n N_Y_c_569_n 0.0205629f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_278_n N_Y_c_569_n 0.00104437f $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_27_47#_M1000_g N_Y_c_586_n 0.0100736f $X=2.88 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_27_47#_M1001_g N_Y_c_586_n 0.0146918f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_27_47#_M1000_g N_Y_c_571_n 0.00152451f $X=2.88 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_27_47#_M1001_g N_Y_c_571_n 0.0153112f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_278_n N_Y_c_571_n 0.00181896f $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1000_g Y 8.95807e-19 $X=2.88 $Y=1.985 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1001_g Y 0.00686543f $X=3.3 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_276_n Y 0.00787629f $X=2.99 $Y=1.19 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_277_n Y 0.0123491f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_278_n Y 0.00996983f $X=3.3 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_273_n N_VGND_c_660_n 0.0155298f $X=1.06 $Y=0.815 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_272_n N_VGND_c_662_n 0.0179318f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_273_n N_VGND_c_662_n 0.00223864f $X=1.06 $Y=0.815 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1014_g N_VGND_c_663_n 0.00357877f $X=2.88 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1018_g N_VGND_c_663_n 0.00357877f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_273_n N_VGND_c_663_n 0.00233669f $X=1.06 $Y=0.815 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_M1017_s N_VGND_c_665_n 0.00234549f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_M1014_g N_VGND_c_665_n 0.00525237f $X=2.88 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A_27_47#_M1018_g N_VGND_c_665_n 0.00655123f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_272_n N_VGND_c_665_n 0.00992225f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_273_n N_VGND_c_665_n 0.00883861f $X=1.06 $Y=0.815 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1014_g N_A_341_47#_c_728_n 0.0107394f $X=2.88 $Y=0.56 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_M1018_g N_A_341_47#_c_728_n 0.00918728f $X=3.3 $Y=0.56 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_276_n N_A_341_47#_c_728_n 0.0190922f $X=2.99 $Y=1.19 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_277_n N_A_341_47#_c_728_n 0.00190279f $X=2.91 $Y=1.16 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_278_n N_A_341_47#_c_728_n 7.98699e-19 $X=3.3 $Y=1.16 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_276_n N_A_341_47#_c_732_n 0.00575495f $X=2.99 $Y=1.19 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1014_g N_A_591_47#_c_752_n 0.00533972f $X=2.88 $Y=0.56 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1018_g N_A_591_47#_c_752_n 0.0140594f $X=3.3 $Y=0.56 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_276_n N_A_591_47#_c_752_n 0.005333f $X=2.99 $Y=1.19 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_277_n N_A_591_47#_c_752_n 0.00963143f $X=2.91 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_278_n N_A_591_47#_c_752_n 0.00234906f $X=3.3 $Y=1.16 $X2=0
+ $Y2=0
cc_277 N_C_M1016_g N_D_M1003_g 0.0138954f $X=4.66 $Y=0.56 $X2=0 $Y2=0
cc_278 N_C_M1013_g N_D_M1002_g 0.0309046f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_279 C N_D_c_432_n 2.06311e-19 $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_280 N_C_c_387_n N_D_c_432_n 0.0192816f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_281 C D 0.00980712f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_282 N_C_c_387_n D 8.59565e-19 $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_283 N_C_M1011_g N_VPWR_c_486_n 0.0158595f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_284 N_C_M1011_g N_VPWR_c_487_n 0.00541359f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_285 N_C_M1013_g N_VPWR_c_487_n 0.00541359f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_286 N_C_M1013_g N_VPWR_c_488_n 0.00146448f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_287 N_C_M1011_g N_VPWR_c_480_n 0.0109543f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_288 N_C_M1013_g N_VPWR_c_480_n 0.00952874f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_289 N_C_M1011_g N_Y_c_570_n 0.0147646f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_290 C N_Y_c_570_n 0.0416536f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_291 N_C_c_386_n N_Y_c_570_n 0.00729564f $X=4.24 $Y=1.16 $X2=0 $Y2=0
cc_292 N_C_M1011_g N_Y_c_612_n 0.0145598f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_293 N_C_M1013_g N_Y_c_612_n 0.00975139f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_294 N_C_M1013_g N_Y_c_572_n 0.0157539f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_295 N_C_M1013_g N_Y_c_615_n 6.1949e-19 $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_296 N_C_M1011_g N_Y_c_574_n 0.00149073f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_297 N_C_M1013_g N_Y_c_574_n 0.00149073f $X=4.66 $Y=1.985 $X2=0 $Y2=0
cc_298 C N_Y_c_574_n 0.026643f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_299 N_C_c_387_n N_Y_c_574_n 0.00206439f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_300 N_C_M1011_g Y 0.00346355f $X=4.24 $Y=1.985 $X2=0 $Y2=0
cc_301 C Y 0.0169443f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_302 N_C_c_386_n Y 0.00107795f $X=4.24 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_M1010_g N_VGND_c_663_n 0.00357877f $X=4.24 $Y=0.56 $X2=0 $Y2=0
cc_304 N_C_M1016_g N_VGND_c_663_n 0.00357877f $X=4.66 $Y=0.56 $X2=0 $Y2=0
cc_305 N_C_M1010_g N_VGND_c_665_n 0.00655123f $X=4.24 $Y=0.56 $X2=0 $Y2=0
cc_306 N_C_M1016_g N_VGND_c_665_n 0.00525237f $X=4.66 $Y=0.56 $X2=0 $Y2=0
cc_307 N_C_M1010_g N_A_591_47#_c_752_n 0.0138053f $X=4.24 $Y=0.56 $X2=0 $Y2=0
cc_308 N_C_M1016_g N_A_591_47#_c_752_n 0.00362121f $X=4.66 $Y=0.56 $X2=0 $Y2=0
cc_309 C N_A_591_47#_c_752_n 0.0665138f $X=4.305 $Y=1.105 $X2=0 $Y2=0
cc_310 N_C_c_386_n N_A_591_47#_c_752_n 0.00758649f $X=4.24 $Y=1.16 $X2=0 $Y2=0
cc_311 N_C_c_387_n N_A_591_47#_c_752_n 0.00207461f $X=4.66 $Y=1.16 $X2=0 $Y2=0
cc_312 N_C_M1010_g N_A_781_47#_c_778_n 0.00918728f $X=4.24 $Y=0.56 $X2=0 $Y2=0
cc_313 N_C_M1016_g N_A_781_47#_c_778_n 0.0129875f $X=4.66 $Y=0.56 $X2=0 $Y2=0
cc_314 N_D_M1002_g N_VPWR_c_488_n 0.00146448f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_315 N_D_M1012_g N_VPWR_c_490_n 0.00411437f $X=5.5 $Y=1.985 $X2=0 $Y2=0
cc_316 D N_VPWR_c_490_n 0.020304f $X=5.685 $Y=1.105 $X2=0 $Y2=0
cc_317 N_D_c_434_n N_VPWR_c_490_n 0.00586305f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_318 N_D_M1002_g N_VPWR_c_494_n 0.00541359f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_319 N_D_M1012_g N_VPWR_c_494_n 0.00541359f $X=5.5 $Y=1.985 $X2=0 $Y2=0
cc_320 N_D_M1002_g N_VPWR_c_480_n 0.00952874f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_321 N_D_M1012_g N_VPWR_c_480_n 0.0104652f $X=5.5 $Y=1.985 $X2=0 $Y2=0
cc_322 N_D_M1002_g N_Y_c_612_n 6.1949e-19 $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_323 N_D_M1002_g N_Y_c_572_n 0.0119784f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_324 N_D_c_432_n N_Y_c_572_n 0.00133007f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_325 D N_Y_c_572_n 0.0127988f $X=5.685 $Y=1.105 $X2=0 $Y2=0
cc_326 N_D_M1002_g N_Y_c_573_n 0.00149073f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_327 N_D_M1012_g N_Y_c_573_n 0.00331821f $X=5.5 $Y=1.985 $X2=0 $Y2=0
cc_328 N_D_c_432_n N_Y_c_573_n 0.00206439f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_329 D N_Y_c_573_n 0.026643f $X=5.685 $Y=1.105 $X2=0 $Y2=0
cc_330 N_D_M1002_g N_Y_c_615_n 0.00975139f $X=5.08 $Y=1.985 $X2=0 $Y2=0
cc_331 N_D_M1012_g N_Y_c_615_n 0.00902485f $X=5.5 $Y=1.985 $X2=0 $Y2=0
cc_332 N_D_M1003_g N_VGND_c_661_n 0.00268723f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_333 N_D_M1007_g N_VGND_c_661_n 0.00268723f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_334 N_D_M1003_g N_VGND_c_663_n 0.00422898f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_335 N_D_M1007_g N_VGND_c_664_n 0.00424416f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_336 N_D_M1003_g N_VGND_c_665_n 0.00577235f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_337 N_D_M1007_g N_VGND_c_665_n 0.00669975f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_338 N_D_M1003_g N_A_781_47#_c_784_n 0.00265763f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_339 N_D_M1003_g N_A_781_47#_c_779_n 0.00482239f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_340 N_D_M1007_g N_A_781_47#_c_779_n 4.58193e-19 $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_341 N_D_c_432_n N_A_781_47#_c_779_n 0.00142286f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_342 D N_A_781_47#_c_779_n 0.00717595f $X=5.685 $Y=1.105 $X2=0 $Y2=0
cc_343 N_D_M1003_g N_A_781_47#_c_780_n 0.00850187f $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_344 N_D_M1007_g N_A_781_47#_c_780_n 0.00973154f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_345 N_D_c_432_n N_A_781_47#_c_780_n 0.00205431f $X=5.575 $Y=1.16 $X2=0 $Y2=0
cc_346 D N_A_781_47#_c_780_n 0.0625861f $X=5.685 $Y=1.105 $X2=0 $Y2=0
cc_347 N_D_c_434_n N_A_781_47#_c_780_n 0.00728275f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_348 N_D_M1003_g N_A_781_47#_c_781_n 5.24843e-19 $X=5.08 $Y=0.56 $X2=0 $Y2=0
cc_349 N_D_M1007_g N_A_781_47#_c_781_n 0.00641402f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_350 N_VPWR_c_480_n N_Y_M1005_s 0.0038878f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_351 N_VPWR_c_480_n N_Y_M1000_s 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_352 N_VPWR_c_480_n N_Y_M1011_s 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_353 N_VPWR_c_480_n N_Y_M1002_d 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_354 N_VPWR_c_483_n N_Y_c_584_n 0.0151499f $X=2.505 $Y=2.72 $X2=0 $Y2=0
cc_355 N_VPWR_c_480_n N_Y_c_584_n 0.00934584f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_356 N_VPWR_M1008_d N_Y_c_569_n 0.00167154f $X=2.535 $Y=1.485 $X2=0 $Y2=0
cc_357 N_VPWR_c_484_n N_Y_c_569_n 0.0146104f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_358 N_VPWR_c_485_n N_Y_c_586_n 0.0189039f $X=3.425 $Y=2.72 $X2=0 $Y2=0
cc_359 N_VPWR_c_480_n N_Y_c_586_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_360 N_VPWR_M1001_d N_Y_c_570_n 0.0102286f $X=3.375 $Y=1.485 $X2=0 $Y2=0
cc_361 N_VPWR_M1001_d N_Y_c_571_n 0.00126437f $X=3.375 $Y=1.485 $X2=0 $Y2=0
cc_362 N_VPWR_c_486_n N_Y_c_571_n 0.0559319f $X=3.95 $Y=2 $X2=0 $Y2=0
cc_363 N_VPWR_c_487_n N_Y_c_612_n 0.0189039f $X=4.785 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_480_n N_Y_c_612_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_M1013_d N_Y_c_572_n 0.00167154f $X=4.735 $Y=1.485 $X2=0 $Y2=0
cc_366 N_VPWR_c_488_n N_Y_c_572_n 0.0129161f $X=4.87 $Y=2 $X2=0 $Y2=0
cc_367 N_VPWR_c_490_n N_Y_c_573_n 0.010848f $X=5.71 $Y=1.66 $X2=0 $Y2=0
cc_368 N_VPWR_c_494_n N_Y_c_615_n 0.0189039f $X=5.625 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_c_480_n N_Y_c_615_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_490_n N_A_781_47#_c_780_n 7.91944e-19 $X=5.71 $Y=1.66 $X2=0
+ $Y2=0
cc_371 N_Y_M1009_d N_VGND_c_665_n 0.00216833f $X=2.115 $Y=0.235 $X2=0 $Y2=0
cc_372 N_Y_M1009_d N_A_341_47#_c_728_n 0.00303391f $X=2.115 $Y=0.235 $X2=0 $Y2=0
cc_373 N_Y_c_576_n N_A_341_47#_c_728_n 0.0161002f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_374 N_Y_c_576_n N_A_591_47#_c_752_n 0.00804581f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_375 N_Y_c_571_n N_A_591_47#_c_752_n 0.0106638f $X=3.55 $Y=1.555 $X2=0 $Y2=0
cc_376 Y N_A_591_47#_c_752_n 0.0239972f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_377 N_Y_c_572_n N_A_781_47#_c_779_n 0.00613486f $X=5.125 $Y=1.555 $X2=0 $Y2=0
cc_378 N_VGND_c_665_n N_A_341_47#_M1009_s 0.00348203f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_379 N_VGND_c_665_n N_A_341_47#_M1015_s 0.00215227f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_665_n N_A_341_47#_M1018_s 0.00209344f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_663_n N_A_341_47#_c_732_n 0.110485f $X=5.205 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_665_n N_A_341_47#_c_732_n 0.0693887f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_665_n N_A_591_47#_M1014_d 0.00216833f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_384 N_VGND_c_665_n N_A_591_47#_M1010_d 0.00216833f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_663_n N_A_591_47#_c_752_n 0.00342407f $X=5.205 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_665_n N_A_591_47#_c_752_n 0.00827928f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_665_n N_A_781_47#_M1010_s 0.00209344f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_388 N_VGND_c_665_n N_A_781_47#_M1016_s 0.00215206f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_665_n N_A_781_47#_M1007_d 0.00209319f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_663_n N_A_781_47#_c_778_n 0.0524263f $X=5.205 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_665_n N_A_781_47#_c_778_n 0.0329788f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_663_n N_A_781_47#_c_784_n 0.0152108f $X=5.205 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_665_n N_A_781_47#_c_784_n 0.00940698f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_M1003_s N_A_781_47#_c_780_n 0.00162006f $X=5.155 $Y=0.235 $X2=0
+ $Y2=0
cc_395 N_VGND_c_661_n N_A_781_47#_c_780_n 0.0122414f $X=5.29 $Y=0.4 $X2=0 $Y2=0
cc_396 N_VGND_c_663_n N_A_781_47#_c_780_n 0.00193763f $X=5.205 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_664_n N_A_781_47#_c_780_n 0.00193763f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_c_665_n N_A_781_47#_c_780_n 0.00825759f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_664_n N_A_781_47#_c_781_n 0.0224042f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_665_n N_A_781_47#_c_781_n 0.0131812f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_401 N_A_341_47#_c_728_n N_A_591_47#_M1014_d 0.00304247f $X=3.51 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_402 N_A_341_47#_M1018_s N_A_591_47#_c_752_n 0.00312742f $X=3.375 $Y=0.235
+ $X2=0 $Y2=0
cc_403 N_A_341_47#_c_728_n N_A_591_47#_c_752_n 0.0410128f $X=3.51 $Y=0.4 $X2=0
+ $Y2=0
cc_404 N_A_341_47#_c_728_n N_A_781_47#_c_778_n 0.0197363f $X=3.51 $Y=0.4 $X2=0
+ $Y2=0
cc_405 N_A_591_47#_c_752_n N_A_781_47#_M1010_s 0.00312742f $X=4.45 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_406 N_A_591_47#_M1010_d N_A_781_47#_c_778_n 0.0030596f $X=4.315 $Y=0.235
+ $X2=0 $Y2=0
cc_407 N_A_591_47#_c_752_n N_A_781_47#_c_778_n 0.0413036f $X=4.45 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_591_47#_c_752_n N_A_781_47#_c_779_n 0.00799569f $X=4.45 $Y=0.74 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__and2_1.spice
* Created: Thu Aug 27 14:06:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2_1.pex.spice"
.subckt sky130_fd_sc_hd__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_145_75# N_A_M1004_g N_A_59_75#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g A_145_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0877682 AS=0.0567 PD=0.816449 PS=0.69 NRD=34.284 NRS=22.848 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_59_75#_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.135832 PD=1.86 PS=1.26355 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_59_75#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_59_75#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0985225 AS=0.0567 PD=0.822254 PS=0.69 NRD=55.1009 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_59_75#_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1
+ AD=0.475 AS=0.234577 PD=2.95 PS=1.95775 NRD=18.715 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.4 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__and2_1.pxi.spice"
*
.ends
*
*

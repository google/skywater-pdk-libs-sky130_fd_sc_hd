* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_2.spice.pex
* Created: Thu Aug 27 14:23:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A 3 7 8 11 12 15
c34 11 0 6.88932e-20 $X=0.505 $Y=1.395
c35 3 0 5.879e-20 $X=0.475 $Y=0.445
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.065 $X2=0.53 $Y2=1.065
r37 12 16 6.88265 $w=3.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.605 $Y=0.85
+ $X2=0.605 $Y2=1.065
r38 10 15 30.6554 $w=3.2e-07 $l=1.7e-07 $layer=POLY_cond $X=0.505 $Y=1.235
+ $X2=0.505 $Y2=1.065
r39 10 11 38.8075 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=0.505 $Y=1.235
+ $X2=0.505 $Y2=1.395
r40 8 15 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.06
+ $X2=0.505 $Y2=1.065
r41 8 9 38.8075 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=0.505 $Y=1.06
+ $X2=0.505 $Y2=0.9
r42 7 11 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=1.985
+ $X2=0.475 $Y2=1.395
r43 3 9 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%A_27_47# 1 2 7 9 10 12 13 15 16
+ 18 20 23 25 29 30 35 37
c72 29 0 1.509e-19 $X=1.05 $Y=1.16
r73 32 35 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.42 $X2=0.26
+ $Y2=0.42
r74 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r75 27 29 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.09 $Y=1.41
+ $X2=1.09 $Y2=1.16
r76 26 37 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=1.495
+ $X2=0.22 $Y2=1.495
r77 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.965 $Y=1.495
+ $X2=1.09 $Y2=1.41
r78 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.965 $Y=1.495
+ $X2=0.355 $Y2=1.495
r79 21 37 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=1.58 $X2=0.22
+ $Y2=1.495
r80 21 23 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.22 $Y=1.58
+ $X2=0.22 $Y2=1.745
r81 20 37 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.17 $Y=1.41
+ $X2=0.22 $Y2=1.495
r82 19 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=0.42
r83 19 20 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.17 $Y2=1.41
r84 16 30 42.1856 $w=2.85e-07 $l=3.23381e-07 $layer=POLY_cond $X=1.37 $Y=1.395
+ $X2=1.16 $Y2=1.16
r85 16 18 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.37 $Y=1.395
+ $X2=1.37 $Y2=1.985
r86 13 30 72.6277 $w=2.85e-07 $l=5.09289e-07 $layer=POLY_cond $X=1.37 $Y=0.745
+ $X2=1.16 $Y2=1.16
r87 13 15 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.37 $Y=0.745 $X2=1.37
+ $Y2=0.445
r88 10 30 42.1856 $w=2.85e-07 $l=3.23381e-07 $layer=POLY_cond $X=0.95 $Y=1.395
+ $X2=1.16 $Y2=1.16
r89 10 12 189.587 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.95 $Y=1.395
+ $X2=0.95 $Y2=1.985
r90 7 30 72.6277 $w=2.85e-07 $l=2.1e-07 $layer=POLY_cond $X=0.95 $Y=1.16
+ $X2=1.16 $Y2=1.16
r91 7 9 96.4 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.95 $Y=1.16 $X2=0.95
+ $Y2=0.445
r92 2 23 300 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.745
r93 1 35 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%KAPWR 1 2 7 13 14 17 18 21 32
r35 18 32 0.00230263 $w=2e-07 $l=3e-09 $layer=MET1_cond $X=0.237 $Y=2.24
+ $X2=0.24 $Y2=2.24
r36 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.58 $Y=2.225
+ $X2=1.58 $Y2=2.225
r37 13 32 0.237939 $w=2e-07 $l=3.1e-07 $layer=MET1_cond $X=0.55 $Y=2.24 $X2=0.24
+ $Y2=2.24
r38 12 21 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.69 $Y=2.21
+ $X2=0.69 $Y2=1.94
r39 11 14 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.695 $Y=2.21
+ $X2=0.84 $Y2=2.21
r40 11 13 0.090534 $w=2.6e-07 $l=1.45e-07 $layer=MET1_cond $X=0.695 $Y=2.21
+ $X2=0.55 $Y2=2.21
r41 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=2.21
+ $X2=0.695 $Y2=2.21
r42 7 16 0.0777288 $w=2.51e-07 $l=1.59295e-07 $layer=MET1_cond $X=1.435 $Y=2.24
+ $X2=1.58 $Y2=2.21
r43 7 14 0.456689 $w=2e-07 $l=5.95e-07 $layer=MET1_cond $X=1.435 $Y=2.24
+ $X2=0.84 $Y2=2.24
r44 2 17 600 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.485 $X2=1.58 $Y2=2.295
r45 1 21 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.94
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%X 1 2 9 13 18 20 21 22 29
c43 20 0 5.879e-20 $X=1.525 $Y=0.765
r44 27 29 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=1.555 $Y=0.825
+ $X2=1.555 $Y2=0.85
r45 21 22 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.555 $Y=1.19
+ $X2=1.555 $Y2=1.53
r46 20 27 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=0.74
+ $X2=1.555 $Y2=0.74
r47 20 21 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=1.555 $Y=0.88
+ $X2=1.555 $Y2=1.19
r48 20 29 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=1.555 $Y=0.88
+ $X2=1.555 $Y2=0.85
r49 18 22 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=1.555 $Y=1.75
+ $X2=1.555 $Y2=1.53
r50 15 18 21.1107 $w=2.18e-07 $l=4.03e-07 $layer=LI1_cond $X=1.152 $Y=1.86
+ $X2=1.555 $Y2=1.86
r51 11 15 1.7811 $w=1.85e-07 $l=1.1e-07 $layer=LI1_cond $X=1.152 $Y=1.97
+ $X2=1.152 $Y2=1.86
r52 11 13 17.9853 $w=1.83e-07 $l=3e-07 $layer=LI1_cond $X=1.152 $Y=1.97
+ $X2=1.152 $Y2=2.27
r53 7 27 26.9444 $w=1.68e-07 $l=4.13e-07 $layer=LI1_cond $X=1.142 $Y=0.74
+ $X2=1.555 $Y2=0.74
r54 7 9 12.714 $w=2.03e-07 $l=2.35e-07 $layer=LI1_cond $X=1.142 $Y=0.655
+ $X2=1.142 $Y2=0.42
r55 2 13 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.485 $X2=1.16 $Y2=2.27
r56 1 9 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.16 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VGND 1 2 9 11 13 15 17 22 28 32
r30 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r31 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r32 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r33 26 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r34 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r35 23 28 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r36 23 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.15
+ $Y2=0
r37 22 31 4.8404 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.627
+ $Y2=0
r38 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.15
+ $Y2=0
r39 17 28 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r40 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.23
+ $Y2=0
r41 15 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r42 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r43 11 31 2.96817 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.582 $Y=0.085
+ $X2=1.627 $Y2=0
r44 11 13 10.8364 $w=3.33e-07 $l=3.15e-07 $layer=LI1_cond $X=1.582 $Y=0.085
+ $X2=1.582 $Y2=0.4
r45 7 28 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r46 7 9 13.2007 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.4
r47 2 13 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.4
r48 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_2%VPWR 1 8 9
r26 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72 $X2=1.61
+ $Y2=2.72
r27 4 8 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=1.61
+ $Y2=2.72
r28 1 9 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 1 4 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends


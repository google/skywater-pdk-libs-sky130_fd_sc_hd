* File: sky130_fd_sc_hd__o2111a_2.spice
* Created: Thu Aug 27 14:33:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2111a_2.pex.spice"
.subckt sky130_fd_sc_hd__o2111a_2  VNB VPB D1 C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1002 N_X_M1002_d N_A_80_21#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1002_d N_A_80_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 A_386_47# N_D1_M1008_g N_A_80_21#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1009 A_458_47# N_C1_M1009_g A_386_47# VNB NSHORT L=0.15 W=0.65 AD=0.12675
+ AS=0.06825 PD=1.04 PS=0.86 NRD=25.836 NRS=9.228 M=1 R=4.33333 SA=75000.5
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1013 N_A_566_47#_M1013_d N_B1_M1013_g A_458_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.12675 PD=1.04 PS=1.04 NRD=11.076 NRS=25.836 M=1 R=4.33333
+ SA=75001.1 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_566_47#_M1013_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.12675 PD=1.04 PS=1.04 NRD=7.38 NRS=9.228 M=1 R=4.33333
+ SA=75001.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_A_566_47#_M1005_d N_A1_M1005_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.12675 PD=1.83 PS=1.04 NRD=0 NRS=12.912 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_80_21#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1012 N_X_M1003_d N_A_80_21#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.365 PD=1.28 PS=1.73 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1010 N_A_80_21#_M1010_d N_D1_M1010_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.365 PD=1.28 PS=1.73 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_A_80_21#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.14 PD=1.39 PS=1.28 NRD=11.8003 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.8 A=0.15 P=2.3 MULT=1
MM1011 N_A_80_21#_M1011_d N_B1_M1011_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=11.8003 NRS=9.8303 M=1 R=6.66667
+ SA=75002.5 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1000 A_674_297# N_A2_M1000_g N_A_80_21#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=27.5603 NRS=9.8303 M=1 R=6.66667
+ SA=75003 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_674_297# VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.195 PD=2.53 PS=1.39 NRD=0 NRS=27.5603 M=1 R=6.66667 SA=75003.5 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_68 VPB 0 1.50018e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hd__o2111a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__a41oi_2.spice.pex
* Created: Thu Aug 27 14:06:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A41OI_2%B1 1 3 4 6 9 13 15 16 28 29
r42 27 29 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.39 $Y=1.16 $X2=1.5
+ $Y2=1.16
r43 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.16 $X2=1.39 $Y2=1.16
r44 25 27 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=1.08 $Y=1.16 $X2=1.39
+ $Y2=1.16
r45 24 25 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=0.98 $Y=1.16 $X2=1.08
+ $Y2=1.16
r46 22 24 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.71 $Y=1.16
+ $X2=0.98 $Y2=1.16
r47 19 22 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.56 $Y=1.16
+ $X2=0.71 $Y2=1.16
r48 16 28 12.9845 $w=2.03e-07 $l=2.4e-07 $layer=LI1_cond $X=1.15 $Y=1.177
+ $X2=1.39 $Y2=1.177
r49 15 16 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=1.177
+ $X2=1.15 $Y2=1.177
r50 15 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.16 $X2=0.71 $Y2=1.16
r51 11 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.325
+ $X2=1.5 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.5 $Y=1.325 $X2=1.5
+ $Y2=1.985
r53 7 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=1.325
+ $X2=1.08 $Y2=1.16
r54 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.08 $Y=1.325 $X2=1.08
+ $Y2=1.985
r55 4 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=0.995
+ $X2=0.98 $Y2=1.16
r56 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.98 $Y=0.995 $X2=0.98
+ $Y2=0.56
r57 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=0.995
+ $X2=0.56 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.56 $Y=0.995 $X2=0.56
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A1 1 3 6 8 10 13 15 20 21
c43 21 0 1.90366e-19 $X=2.34 $Y=1.16
c44 8 0 1.21078e-19 $X=2.34 $Y=0.995
c45 6 0 1.85225e-19 $X=1.92 $Y=1.985
r46 19 21 7.50779 $w=3.21e-07 $l=5e-08 $layer=POLY_cond $X=2.29 $Y=1.16 $X2=2.34
+ $Y2=1.16
r47 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.16 $X2=2.29 $Y2=1.16
r48 17 19 55.5576 $w=3.21e-07 $l=3.7e-07 $layer=POLY_cond $X=1.92 $Y=1.16
+ $X2=2.29 $Y2=1.16
r49 15 20 11.5244 $w=2.18e-07 $l=2.2e-07 $layer=LI1_cond $X=2.07 $Y=1.185
+ $X2=2.29 $Y2=1.185
r50 11 21 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.325
+ $X2=2.34 $Y2=1.16
r51 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.34 $Y=1.325
+ $X2=2.34 $Y2=1.985
r52 8 21 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=0.995
+ $X2=2.34 $Y2=1.16
r53 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.34 $Y=0.995
+ $X2=2.34 $Y2=0.56
r54 4 17 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.325
+ $X2=1.92 $Y2=1.16
r55 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.92 $Y=1.325 $X2=1.92
+ $Y2=1.985
r56 1 17 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=0.995
+ $X2=1.92 $Y2=1.16
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.92 $Y=0.995 $X2=1.92
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A2 3 7 11 15 17 23 24
r43 22 24 2.22174 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=3.17 $Y=1.16 $X2=3.18
+ $Y2=1.16
r44 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.16 $X2=3.17 $Y2=1.16
r45 19 22 91.0912 $w=2.7e-07 $l=4.1e-07 $layer=POLY_cond $X=2.76 $Y=1.16
+ $X2=3.17 $Y2=1.16
r46 17 23 0.512605 $w=6.98e-07 $l=3e-08 $layer=LI1_cond $X=3.015 $Y=1.19
+ $X2=3.015 $Y2=1.16
r47 13 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.295
+ $X2=3.18 $Y2=1.16
r48 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.18 $Y=1.295
+ $X2=3.18 $Y2=1.985
r49 9 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.18 $Y=1.025
+ $X2=3.18 $Y2=1.16
r50 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.18 $Y=1.025
+ $X2=3.18 $Y2=0.56
r51 5 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=1.295
+ $X2=2.76 $Y2=1.16
r52 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.76 $Y=1.295 $X2=2.76
+ $Y2=1.985
r53 1 19 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=1.025
+ $X2=2.76 $Y2=1.16
r54 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.76 $Y=1.025
+ $X2=2.76 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A3 3 7 11 15 17 18 19 22 30
r49 28 30 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=4.41 $Y=1.16
+ $X2=4.54 $Y2=1.16
r50 26 28 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=4.12 $Y=1.16
+ $X2=4.41 $Y2=1.16
r51 24 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.16 $X2=3.71 $Y2=1.16
r52 22 26 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.12 $Y2=1.16
r53 22 24 74.4282 $w=2.7e-07 $l=3.35e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.71 $Y2=1.16
r54 19 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.41
+ $Y=1.16 $X2=4.41 $Y2=1.16
r55 18 19 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=3.93 $Y=1.185
+ $X2=4.39 $Y2=1.185
r56 18 25 11.5244 $w=2.18e-07 $l=2.2e-07 $layer=LI1_cond $X=3.93 $Y=1.185
+ $X2=3.71 $Y2=1.185
r57 17 24 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=3.695 $Y=1.16
+ $X2=3.71 $Y2=1.16
r58 13 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.54 $Y=1.295
+ $X2=4.54 $Y2=1.16
r59 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.54 $Y=1.295
+ $X2=4.54 $Y2=1.985
r60 9 30 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.54 $Y=1.025
+ $X2=4.54 $Y2=1.16
r61 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.54 $Y=1.025
+ $X2=4.54 $Y2=0.56
r62 5 26 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.12 $Y=1.025
+ $X2=4.12 $Y2=1.16
r63 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.12 $Y=1.025
+ $X2=4.12 $Y2=0.56
r64 1 17 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.62 $Y=1.295
+ $X2=3.695 $Y2=1.16
r65 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.62 $Y=1.295 $X2=3.62
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A4 3 7 11 15 17 18 19 23 25
c39 23 0 1.90366e-19 $X=5.455 $Y=1.16
r40 30 32 61.5693 $w=2.74e-07 $l=3.5e-07 $layer=POLY_cond $X=5.03 $Y=1.16
+ $X2=5.38 $Y2=1.16
r41 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.03
+ $Y=1.16 $X2=5.03 $Y2=1.16
r42 23 32 12.6663 $w=2.9e-07 $l=7.5e-08 $layer=POLY_cond $X=5.455 $Y=1.16
+ $X2=5.38 $Y2=1.16
r43 23 25 52.7471 $w=2.9e-07 $l=2.55e-07 $layer=POLY_cond $X=5.455 $Y=1.16
+ $X2=5.71 $Y2=1.16
r44 19 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=1.16 $X2=5.71 $Y2=1.16
r45 18 19 22.0012 $w=2.18e-07 $l=4.2e-07 $layer=LI1_cond $X=5.29 $Y=1.185
+ $X2=5.71 $Y2=1.185
r46 18 31 13.6198 $w=2.18e-07 $l=2.6e-07 $layer=LI1_cond $X=5.29 $Y=1.185
+ $X2=5.03 $Y2=1.185
r47 17 31 9.42908 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=4.85 $Y=1.185
+ $X2=5.03 $Y2=1.185
r48 13 32 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.38 $Y=1.305
+ $X2=5.38 $Y2=1.16
r49 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.38 $Y=1.305
+ $X2=5.38 $Y2=1.985
r50 9 32 16.847 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.38 $Y=1.015
+ $X2=5.38 $Y2=1.16
r51 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.38 $Y=1.015
+ $X2=5.38 $Y2=0.56
r52 1 30 12.3139 $w=2.74e-07 $l=7e-08 $layer=POLY_cond $X=4.96 $Y=1.16 $X2=5.03
+ $Y2=1.16
r53 1 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.96 $Y=1.295 $X2=4.96
+ $Y2=1.985
r54 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.96 $Y=1.025
+ $X2=4.96 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A_149_297# 1 2 3 4 5 6 21 23 24 29 30 33 35
+ 39 41 45 47 51 54 55
c57 55 0 1.90366e-19 $X=4.75 $Y=1.62
c58 30 0 1.90366e-19 $X=1.795 $Y=1.62
r59 49 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.59 $Y=1.705
+ $X2=5.59 $Y2=1.96
r60 48 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=1.62
+ $X2=4.75 $Y2=1.62
r61 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.505 $Y=1.62
+ $X2=5.59 $Y2=1.705
r62 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.505 $Y=1.62
+ $X2=4.835 $Y2=1.62
r63 43 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=1.705
+ $X2=4.75 $Y2=1.62
r64 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.75 $Y=1.705
+ $X2=4.75 $Y2=1.96
r65 42 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=1.62
+ $X2=3.41 $Y2=1.62
r66 41 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=1.62
+ $X2=4.75 $Y2=1.62
r67 41 42 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.665 $Y=1.62
+ $X2=3.495 $Y2=1.62
r68 37 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.705
+ $X2=3.41 $Y2=1.62
r69 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.41 $Y=1.705
+ $X2=3.41 $Y2=1.96
r70 36 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=1.62
+ $X2=2.55 $Y2=1.62
r71 35 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.62
+ $X2=3.41 $Y2=1.62
r72 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.325 $Y=1.62
+ $X2=2.635 $Y2=1.62
r73 31 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=1.705
+ $X2=2.55 $Y2=1.62
r74 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.55 $Y=1.705
+ $X2=2.55 $Y2=1.96
r75 29 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=1.62
+ $X2=2.55 $Y2=1.62
r76 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.465 $Y=1.62
+ $X2=1.795 $Y2=1.62
r77 26 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.71 $Y=2.295
+ $X2=1.71 $Y2=1.96
r78 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.71 $Y=1.705
+ $X2=1.795 $Y2=1.62
r79 25 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.71 $Y=1.705
+ $X2=1.71 $Y2=1.96
r80 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.625 $Y=2.38
+ $X2=1.71 $Y2=2.295
r81 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.625 $Y=2.38
+ $X2=0.955 $Y2=2.38
r82 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.87 $Y=2.295
+ $X2=0.955 $Y2=2.38
r83 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.87 $Y=2.295
+ $X2=0.87 $Y2=1.96
r84 6 51 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.455
+ $Y=1.485 $X2=5.59 $Y2=1.96
r85 5 45 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.615
+ $Y=1.485 $X2=4.75 $Y2=1.96
r86 4 39 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=3.255
+ $Y=1.485 $X2=3.41 $Y2=1.96
r87 3 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.415
+ $Y=1.485 $X2=2.55 $Y2=1.96
r88 2 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.575
+ $Y=1.485 $X2=1.71 $Y2=1.96
r89 1 21 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.745
+ $Y=1.485 $X2=0.87 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%Y 1 2 3 12 16 20 22 23 24 25 26 27 35 36 38
c54 20 0 1.85225e-19 $X=1.29 $Y=1.7
r55 35 38 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.23 $Y=0.815
+ $X2=0.23 $Y2=0.85
r56 27 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=1.54 $X2=0.23
+ $Y2=1.455
r57 27 36 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.23 $Y=1.45 $X2=0.23
+ $Y2=1.455
r58 26 27 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.23 $Y2=1.45
r59 25 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=0.73 $X2=0.23
+ $Y2=0.815
r60 25 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.23 $Y=0.875
+ $X2=0.23 $Y2=1.19
r61 25 38 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=0.875
+ $X2=0.23 $Y2=0.85
r62 24 27 29.6808 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=1.125 $Y=1.54
+ $X2=0.315 $Y2=1.54
r63 22 25 20.0073 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.685 $Y=0.73
+ $X2=0.315 $Y2=0.73
r64 22 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.73
+ $X2=0.77 $Y2=0.73
r65 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.29 $Y=1.625
+ $X2=1.125 $Y2=1.54
r66 18 20 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.29 $Y=1.625
+ $X2=1.29 $Y2=1.7
r67 14 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.73
+ $X2=0.77 $Y2=0.73
r68 14 16 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=0.855 $Y=0.73
+ $X2=2.13 $Y2=0.73
r69 10 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.645
+ $X2=0.77 $Y2=0.73
r70 10 12 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.77 $Y=0.645
+ $X2=0.77 $Y2=0.42
r71 3 20 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=1.155
+ $Y=1.485 $X2=1.29 $Y2=1.7
r72 2 16 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.235 $X2=2.13 $Y2=0.73
r73 1 12 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.235 $X2=0.77 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%VPWR 1 2 3 4 15 19 23 27 30 31 32 34 42 47
+ 57 58 61 64 67
r76 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r78 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r79 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r80 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r81 55 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r82 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r83 52 67 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.09 $Y2=2.72
r84 52 54 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.425 $Y=2.72
+ $X2=4.83 $Y2=2.72
r85 51 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r86 51 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r87 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=2.97 $Y2=2.72
r89 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.45 $Y2=2.72
r90 47 67 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=4.09 $Y2=2.72
r91 47 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r92 46 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r93 46 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r94 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r95 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.13 $Y2=2.72
r96 43 45 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.53 $Y2=2.72
r97 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=2.97 $Y2=2.72
r98 42 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.805 $Y=2.72
+ $X2=2.53 $Y2=2.72
r99 41 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r101 36 40 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r102 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=2.72
+ $X2=2.13 $Y2=2.72
r103 34 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.965 $Y=2.72
+ $X2=1.61 $Y2=2.72
r104 32 41 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r105 32 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r106 30 54 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=4.83 $Y2=2.72
r107 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=5.17 $Y2=2.72
r108 29 57 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.335 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=2.72
+ $X2=5.17 $Y2=2.72
r110 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=2.635
+ $X2=5.17 $Y2=2.72
r111 25 27 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.17 $Y=2.635
+ $X2=5.17 $Y2=2
r112 21 67 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=2.635
+ $X2=4.09 $Y2=2.72
r113 21 23 11.336 $w=6.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.09 $Y=2.635
+ $X2=4.09 $Y2=2
r114 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.72
r115 17 19 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2
r116 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=2.635
+ $X2=2.13 $Y2=2.72
r117 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.13 $Y=2.635
+ $X2=2.13 $Y2=2
r118 4 27 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.035
+ $Y=1.485 $X2=5.17 $Y2=2
r119 3 23 150 $w=1.7e-07 $l=7.81153e-07 $layer=licon1_PDIFF $count=4 $X=3.695
+ $Y=1.485 $X2=4.26 $Y2=2
r120 2 19 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.835
+ $Y=1.485 $X2=2.97 $Y2=2
r121 1 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.13 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r79 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r80 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r81 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r82 37 38 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r83 35 38 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=4.83
+ $Y2=0
r84 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r85 34 37 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=4.83
+ $Y2=0
r86 34 35 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r87 32 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.2
+ $Y2=0
r88 32 34 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.61
+ $Y2=0
r89 31 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r90 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r91 28 44 4.59558 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.257
+ $Y2=0
r92 28 30 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.69
+ $Y2=0
r93 27 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.2
+ $Y2=0
r94 27 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.69
+ $Y2=0
r95 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r96 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r97 23 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=4.83
+ $Y2=0
r98 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.17
+ $Y2=0
r99 22 40 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.75
+ $Y2=0
r100 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.17
+ $Y2=0
r101 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0
r102 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.17 $Y=0.085
+ $X2=5.17 $Y2=0.38
r103 14 47 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r104 14 16 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.38
r105 10 44 3.17059 $w=3.3e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.257 $Y2=0
r106 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.35 $Y2=0.38
r107 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.035
+ $Y=0.235 $X2=5.17 $Y2=0.38
r108 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.235 $X2=1.19 $Y2=0.38
r109 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A_317_47# 1 2 3 10 18
r26 16 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.73
+ $X2=2.55 $Y2=0.73
r27 16 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.635 $Y=0.73
+ $X2=3.39 $Y2=0.73
r28 15 21 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.55 $Y=0.645
+ $X2=2.55 $Y2=0.73
r29 14 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.55 $Y=0.465
+ $X2=2.55 $Y2=0.645
r30 10 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=0.38
+ $X2=2.55 $Y2=0.465
r31 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.465 $Y=0.38
+ $X2=1.71 $Y2=0.38
r32 3 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.235 $X2=3.39 $Y2=0.73
r33 2 21 182 $w=1.7e-07 $l=4.77755e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.55 $Y2=0.65
r34 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A_567_47# 1 2 11
c19 11 0 1.21078e-19 $X=4.33 $Y=0.38
r20 8 11 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.97 $Y=0.38
+ $X2=4.33 $Y2=0.38
r21 2 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.195
+ $Y=0.235 $X2=4.33 $Y2=0.38
r22 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.235 $X2=2.97 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A41OI_2%A_757_47# 1 2 3 10 18
r25 16 18 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.59 $Y=0.645
+ $X2=5.59 $Y2=0.42
r26 12 15 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.91 $Y=0.73
+ $X2=4.75 $Y2=0.73
r27 10 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.505 $Y=0.73
+ $X2=5.59 $Y2=0.645
r28 10 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.505 $Y=0.73
+ $X2=4.75 $Y2=0.73
r29 3 18 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.455
+ $Y=0.235 $X2=5.59 $Y2=0.42
r30 2 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.235 $X2=4.75 $Y2=0.73
r31 1 12 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.235 $X2=3.91 $Y2=0.73
.ends


* File: sky130_fd_sc_hd__nand2b_4.pex.spice
* Created: Tue Sep  1 19:15:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NAND2B_4%A_N 3 7 9 15
c26 9 0 1.2849e-19 $X=0.235 $Y=1.19
r27 12 15 40.336 $w=2.9e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r28 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r29 5 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r30 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r31 1 15 18.1727 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r32 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 48 50 56 61 66 68 69 76
c121 69 0 1.2849e-19 $X=1.335 $Y=1.16
r122 75 76 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.67 $Y2=1.16
r123 72 73 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=1.41 $Y=1.16
+ $X2=1.83 $Y2=1.16
r124 69 72 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.16
+ $X2=1.41 $Y2=1.16
r125 57 75 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.04 $Y=1.16
+ $X2=2.25 $Y2=1.16
r126 57 73 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=2.04 $Y=1.16
+ $X2=1.83 $Y2=1.16
r127 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.16 $X2=2.04 $Y2=1.16
r128 54 69 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.16
+ $X2=1.335 $Y2=1.16
r129 53 56 48.2455 $w=1.98e-07 $l=8.7e-07 $layer=LI1_cond $X=1.17 $Y=1.175
+ $X2=2.04 $Y2=1.175
r130 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.16 $X2=1.17 $Y2=1.16
r131 51 68 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.175
+ $X2=0.695 $Y2=1.175
r132 51 53 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=0.78 $Y=1.175
+ $X2=1.17 $Y2=1.175
r133 50 66 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.695 $Y=1.445
+ $X2=0.695 $Y2=1.555
r134 49 68 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.275
+ $X2=0.695 $Y2=1.175
r135 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.695 $Y=1.275
+ $X2=0.695 $Y2=1.445
r136 48 68 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=1.175
r137 47 61 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.695 $Y=0.905
+ $X2=0.695 $Y2=0.81
r138 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.695 $Y=0.905
+ $X2=0.695 $Y2=1.075
r139 43 66 22.9441 $w=2.18e-07 $l=4.38e-07 $layer=LI1_cond $X=0.257 $Y=1.555
+ $X2=0.695 $Y2=1.555
r140 43 45 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.34
r141 39 61 25.5675 $w=1.88e-07 $l=4.38e-07 $layer=LI1_cond $X=0.257 $Y=0.81
+ $X2=0.695 $Y2=0.81
r142 39 41 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r143 35 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.16
r144 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.985
r145 31 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=1.16
r146 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.67 $Y=1.025
+ $X2=2.67 $Y2=0.56
r147 27 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.16
r148 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.985
r149 23 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=1.16
r150 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.25 $Y=1.025
+ $X2=2.25 $Y2=0.56
r151 19 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.16
r152 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.83 $Y=1.295
+ $X2=1.83 $Y2=1.985
r153 15 73 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=1.16
r154 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.83 $Y=1.025
+ $X2=1.83 $Y2=0.56
r155 11 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.16
r156 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.41 $Y=1.295
+ $X2=1.41 $Y2=1.985
r157 7 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.16
r158 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r159 2 43 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r160 2 45 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r161 1 41 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%B 3 7 11 15 19 23 27 31 33 34 35 36 41 43
c88 3 0 8.71462e-20 $X=3.105 $Y=0.56
r89 52 53 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.945 $Y=1.16
+ $X2=4.365 $Y2=1.16
r90 51 52 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=3.525 $Y=1.16
+ $X2=3.945 $Y2=1.16
r91 49 51 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=3.32 $Y=1.16
+ $X2=3.525 $Y2=1.16
r92 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r93 46 49 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=3.105 $Y=1.16
+ $X2=3.32 $Y2=1.16
r94 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.16 $X2=4.605 $Y2=1.16
r95 41 53 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.365 $Y2=1.16
r96 41 43 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=1.16
+ $X2=4.605 $Y2=1.16
r97 36 44 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=4.605 $Y2=1.175
r98 35 44 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.605 $Y2=1.175
r99 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.395 $Y2=1.175
r100 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.935 $Y2=1.175
r101 33 50 8.59545 $w=1.98e-07 $l=1.55e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.32 $Y2=1.175
r102 29 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.365 $Y=1.295
+ $X2=4.365 $Y2=1.16
r103 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.365 $Y=1.295
+ $X2=4.365 $Y2=1.985
r104 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.365 $Y=1.025
+ $X2=4.365 $Y2=1.16
r105 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.365 $Y=1.025
+ $X2=4.365 $Y2=0.56
r106 21 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.945 $Y=1.295
+ $X2=3.945 $Y2=1.16
r107 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.945 $Y=1.295
+ $X2=3.945 $Y2=1.985
r108 17 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.945 $Y=1.025
+ $X2=3.945 $Y2=1.16
r109 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.945 $Y=1.025
+ $X2=3.945 $Y2=0.56
r110 13 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.525 $Y=1.295
+ $X2=3.525 $Y2=1.16
r111 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.525 $Y=1.295
+ $X2=3.525 $Y2=1.985
r112 9 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.525 $Y=1.025
+ $X2=3.525 $Y2=1.16
r113 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.525 $Y=1.025
+ $X2=3.525 $Y2=0.56
r114 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.16
r115 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.985
r116 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.105 $Y=1.025
+ $X2=3.105 $Y2=1.16
r117 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.105 $Y=1.025
+ $X2=3.105 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%VPWR 1 2 3 4 5 6 22 25 29 33 37 39 41 46 49
+ 50 52 53 55 56 57 59 74 79 83
r81 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r82 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 77 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r84 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 74 82 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=4.52 $Y=2.72 $X2=4.79
+ $Y2=2.72
r86 74 76 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.52 $Y=2.72 $X2=4.37
+ $Y2=2.72
r87 73 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r88 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r90 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r91 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r92 67 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 64 79 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=0.94 $Y2=2.72
r95 64 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.61 $Y2=2.72
r96 59 79 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.94 $Y2=2.72
r97 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r98 57 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r99 57 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r100 55 72 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.65 $Y=2.72 $X2=3.45
+ $Y2=2.72
r101 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=2.72
+ $X2=3.735 $Y2=2.72
r102 54 76 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.735 $Y2=2.72
r104 52 69 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.895 $Y2=2.72
r106 51 72 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.72
+ $X2=2.895 $Y2=2.72
r108 49 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.04 $Y2=2.72
r110 48 69 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.53 $Y2=2.72
r111 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=2.72
+ $X2=2.04 $Y2=2.72
r112 46 47 6.43014 $w=6.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=2 $X2=0.94
+ $Y2=1.835
r113 41 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.685 $Y=1.66
+ $X2=4.685 $Y2=2.34
r114 39 82 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.685 $Y=2.635
+ $X2=4.79 $Y2=2.72
r115 39 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.685 $Y=2.635
+ $X2=4.685 $Y2=2.34
r116 35 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=2.635
+ $X2=3.735 $Y2=2.72
r117 35 37 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=2.635
+ $X2=3.735 $Y2=2
r118 31 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.635
+ $X2=2.895 $Y2=2.72
r119 31 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.895 $Y=2.635
+ $X2=2.895 $Y2=2
r120 27 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2.72
r121 27 29 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.04 $Y=2.635
+ $X2=2.04 $Y2=2
r122 25 47 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=1.127 $Y=1.66
+ $X2=1.127 $Y2=1.835
r123 20 79 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.72
r124 20 22 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.94 $Y=2.635
+ $X2=0.94 $Y2=2.34
r125 19 46 3.1202 $w=6.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.94 $Y=2.18
+ $X2=0.94 $Y2=2
r126 19 22 2.77352 $w=6.88e-07 $l=1.6e-07 $layer=LI1_cond $X=0.94 $Y=2.18
+ $X2=0.94 $Y2=2.34
r127 6 44 400 $w=1.7e-07 $l=9.69794e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.485 $X2=4.685 $Y2=2.34
r128 6 41 400 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.485 $X2=4.685 $Y2=1.66
r129 5 37 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.6
+ $Y=1.485 $X2=3.735 $Y2=2
r130 4 33 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.895 $Y2=2
r131 3 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=2
r132 2 25 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.66
r133 2 22 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=2.34
r134 1 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%Y 1 2 3 4 5 6 19 23 25 27 31 35 37 39 41 45
+ 47 50 51 52 59
c95 59 0 8.71462e-20 $X=2.507 $Y=0.905
c96 47 0 1.4834e-19 $X=3.315 $Y=1.66
r97 51 52 8.50329 $w=4.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.507 $Y=1.19
+ $X2=2.507 $Y2=1.445
r98 50 59 3.44693 $w=2.65e-07 $l=1.35e-07 $layer=LI1_cond $X=2.507 $Y=0.77
+ $X2=2.507 $Y2=0.905
r99 50 51 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=2.507 $Y=0.92
+ $X2=2.507 $Y2=1.19
r100 50 59 0.652326 $w=2.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.507 $Y=0.92
+ $X2=2.507 $Y2=0.905
r101 45 52 16.3436 $w=3.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.15 $Y=1.555
+ $X2=2.64 $Y2=1.555
r102 45 47 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=1.555
+ $X2=3.315 $Y2=1.555
r103 39 49 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.155 $Y=1.665
+ $X2=4.155 $Y2=1.555
r104 39 41 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.155 $Y=1.665
+ $X2=4.155 $Y2=2.34
r105 38 47 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=1.555
+ $X2=3.315 $Y2=1.555
r106 37 49 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=1.555
+ $X2=4.155 $Y2=1.555
r107 37 38 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=3.99 $Y=1.555
+ $X2=3.48 $Y2=1.555
r108 33 47 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.315 $Y=1.665
+ $X2=3.315 $Y2=1.555
r109 33 35 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.315 $Y=1.665
+ $X2=3.315 $Y2=2.34
r110 29 52 2.11712 $w=3.45e-07 $l=1.1e-07 $layer=LI1_cond $X=2.467 $Y=1.665
+ $X2=2.467 $Y2=1.555
r111 29 31 22.5478 $w=3.43e-07 $l=6.75e-07 $layer=LI1_cond $X=2.467 $Y=1.665
+ $X2=2.467 $Y2=2.34
r112 28 44 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=1.555
+ $X2=1.62 $Y2=1.555
r113 27 52 4.10039 $w=2.2e-07 $l=1.72e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=2.467 $Y2=1.555
r114 27 28 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=2.295 $Y=1.555
+ $X2=1.785 $Y2=1.555
r115 23 44 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.555
r116 23 25 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2.34
r117 19 50 3.37033 $w=2.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.375 $Y=0.77
+ $X2=2.507 $Y2=0.77
r118 19 21 32.2257 $w=2.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.375 $Y=0.77
+ $X2=1.62 $Y2=0.77
r119 6 49 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.485 $X2=4.155 $Y2=1.66
r120 6 41 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.485 $X2=4.155 $Y2=2.34
r121 5 47 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.315 $Y2=1.66
r122 5 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.485 $X2=3.315 $Y2=2.34
r123 4 52 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=1.66
r124 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.485 $X2=2.46 $Y2=2.34
r125 3 44 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=1.66
r126 3 25 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.485 $X2=1.62 $Y2=2.34
r127 2 50 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.46 $Y2=0.72
r128 1 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.62 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r73 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r74 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r75 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r76 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r77 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r78 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r79 38 41 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r80 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r81 37 40 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r82 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r83 35 50 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.692
+ $Y2=0
r84 35 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=1.15
+ $Y2=0
r85 30 50 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.692
+ $Y2=0
r86 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r87 28 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r88 28 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r89 26 43 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.91
+ $Y2=0
r90 26 27 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.19
+ $Y2=0
r91 25 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.83
+ $Y2=0
r92 25 27 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.31 $Y=0 $X2=4.19
+ $Y2=0
r93 23 40 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.23 $Y=0 $X2=2.99
+ $Y2=0
r94 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.315
+ $Y2=0
r95 22 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.91
+ $Y2=0
r96 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.315
+ $Y2=0
r97 18 27 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0
r98 18 20 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0.38
r99 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r100 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.38
r101 10 50 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r102 10 12 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.38
r103 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.155 $Y2=0.38
r104 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.18
+ $Y=0.235 $X2=3.315 $Y2=0.38
r105 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__NAND2B_4%A_215_47# 1 2 3 4 5 16 18 20 24 25 26 30 32
+ 36 44
c78 26 0 1.4834e-19 $X=3.57 $Y=0.81
r79 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.685 $Y=0.715
+ $X2=4.685 $Y2=0.38
r80 33 44 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=0.81
+ $X2=3.735 $Y2=0.81
r81 32 34 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.52 $Y=0.81
+ $X2=4.685 $Y2=0.715
r82 32 33 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=4.52 $Y=0.81 $X2=3.9
+ $Y2=0.81
r83 28 44 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.735 $Y=0.715
+ $X2=3.735 $Y2=0.81
r84 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.735 $Y=0.715
+ $X2=3.735 $Y2=0.38
r85 27 43 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=0.81
+ $X2=2.935 $Y2=0.81
r86 26 44 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.57 $Y=0.81
+ $X2=3.735 $Y2=0.81
r87 26 27 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.57 $Y=0.81
+ $X2=3.06 $Y2=0.81
r88 25 43 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.935 $Y=0.715
+ $X2=2.935 $Y2=0.81
r89 24 41 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.935 $Y=0.465
+ $X2=2.935 $Y2=0.36
r90 24 25 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.935 $Y=0.465
+ $X2=2.935 $Y2=0.715
r91 21 39 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=1.16 $Y2=0.36
r92 21 23 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=2.04 $Y2=0.36
r93 20 41 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.81 $Y=0.36
+ $X2=2.935 $Y2=0.36
r94 20 23 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=2.81 $Y=0.36
+ $X2=2.04 $Y2=0.36
r95 16 39 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.36
r96 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.72
r97 5 36 91 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.235 $X2=4.685 $Y2=0.38
r98 4 30 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.6
+ $Y=0.235 $X2=3.735 $Y2=0.38
r99 3 43 182 $w=1.7e-07 $l=5.54955e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.895 $Y2=0.72
r100 3 41 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.895 $Y2=0.38
r101 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.38
r102 1 39 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.38
r103 1 18 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.72
.ends


* File: sky130_fd_sc_hd__einvp_1.pxi.spice
* Created: Tue Sep  1 19:08:14 2020
* 
x_PM_SKY130_FD_SC_HD__EINVP_1%TE N_TE_M1004_g N_TE_M1003_g N_TE_c_42_n
+ N_TE_c_43_n N_TE_c_44_n N_TE_M1005_g TE TE PM_SKY130_FD_SC_HD__EINVP_1%TE
x_PM_SKY130_FD_SC_HD__EINVP_1%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1003_s
+ N_A_27_47#_M1002_g N_A_27_47#_c_79_n N_A_27_47#_c_85_n N_A_27_47#_c_80_n
+ N_A_27_47#_c_81_n N_A_27_47#_c_86_n N_A_27_47#_c_87_n N_A_27_47#_c_82_n
+ N_A_27_47#_c_83_n PM_SKY130_FD_SC_HD__EINVP_1%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVP_1%A N_A_c_145_n N_A_M1000_g N_A_M1001_g A A A
+ N_A_c_147_n PM_SKY130_FD_SC_HD__EINVP_1%A
x_PM_SKY130_FD_SC_HD__EINVP_1%VPWR N_VPWR_M1003_d N_VPWR_c_175_n N_VPWR_c_176_n
+ N_VPWR_c_177_n N_VPWR_c_178_n VPWR N_VPWR_c_179_n N_VPWR_c_174_n
+ PM_SKY130_FD_SC_HD__EINVP_1%VPWR
x_PM_SKY130_FD_SC_HD__EINVP_1%Z N_Z_M1000_d N_Z_M1001_d N_Z_c_208_n Z Z
+ N_Z_c_209_n PM_SKY130_FD_SC_HD__EINVP_1%Z
x_PM_SKY130_FD_SC_HD__EINVP_1%VGND N_VGND_M1004_d VGND N_VGND_c_242_n
+ N_VGND_c_243_n N_VGND_c_244_n N_VGND_c_245_n PM_SKY130_FD_SC_HD__EINVP_1%VGND
cc_1 VNB N_TE_M1004_g 0.0344171f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_c_42_n 0.0306674f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.035
cc_3 VNB N_TE_c_43_n 0.0391157f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.035
cc_4 VNB N_TE_c_44_n 0.0163246f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.96
cc_5 VNB TE 0.0149293f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_27_47#_c_79_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_7 VNB N_A_27_47#_c_80_n 0.00414379f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_8 VNB N_A_27_47#_c_81_n 0.00940848f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_9 VNB N_A_27_47#_c_82_n 0.00295656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_83_n 0.0290413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_145_n 0.0254248f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_12 VNB A 0.0141773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_c_147_n 0.0355645f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_174_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Z_c_208_n 0.00265178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_Z_c_209_n 0.0237445f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB N_VGND_c_242_n 0.0234438f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_18 VNB N_VGND_c_243_n 0.142377f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_19 VNB N_VGND_c_244_n 0.0143174f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.132
cc_20 VNB N_VGND_c_245_n 0.0174669f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.53
cc_21 VPB N_TE_M1003_g 0.0726954f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_22 VPB N_TE_c_43_n 0.00815016f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_23 VPB TE 0.020344f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_24 VPB N_A_27_47#_M1002_g 0.0203531f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.035
cc_25 VPB N_A_27_47#_c_85_n 0.0155207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_86_n 0.00421245f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.132
cc_27 VPB N_A_27_47#_c_87_n 0.00974254f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_28 VPB N_A_27_47#_c_82_n 0.00432875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_83_n 0.00597707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_M1001_g 0.0223055f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_31 VPB A 0.0254958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_c_147_n 0.0121578f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_175_n 0.00489839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_176_n 0.0143174f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_35 VPB N_VPWR_c_177_n 0.0076689f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_178_n 0.00572156f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.035
cc_37 VPB N_VPWR_c_179_n 0.0228069f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_38 VPB N_VPWR_c_174_n 0.0433952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Z_c_208_n 0.00111361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB Z 0.0149768f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_41 N_TE_M1003_g N_A_27_47#_M1002_g 0.0074303f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_42 N_TE_M1004_g N_A_27_47#_c_80_n 0.0133028f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_43 N_TE_c_42_n N_A_27_47#_c_80_n 0.0028268f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_44 N_TE_c_43_n N_A_27_47#_c_80_n 3.31368e-19 $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_45 N_TE_c_44_n N_A_27_47#_c_80_n 0.0105602f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_46 TE N_A_27_47#_c_80_n 0.0155346f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_47 N_TE_c_43_n N_A_27_47#_c_81_n 0.00172695f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_48 TE N_A_27_47#_c_81_n 0.0239473f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_49 N_TE_M1003_g N_A_27_47#_c_86_n 0.014462f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_50 TE N_A_27_47#_c_86_n 0.0155353f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_51 N_TE_c_43_n N_A_27_47#_c_87_n 7.77994e-19 $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_52 TE N_A_27_47#_c_87_n 0.0239512f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_53 N_TE_M1004_g N_A_27_47#_c_82_n 0.00374902f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_54 N_TE_c_42_n N_A_27_47#_c_82_n 0.0182646f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_55 N_TE_c_43_n N_A_27_47#_c_82_n 0.0118596f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_56 N_TE_c_44_n N_A_27_47#_c_82_n 0.00591461f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_57 TE N_A_27_47#_c_82_n 0.0617392f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_TE_c_42_n N_A_27_47#_c_83_n 0.00748335f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_59 N_TE_c_43_n N_A_27_47#_c_83_n 0.0074303f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_60 TE N_A_27_47#_c_83_n 4.42301e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_61 N_TE_M1003_g N_VPWR_c_175_n 0.00981763f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_62 N_TE_M1003_g N_VPWR_c_176_n 0.00341689f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_63 N_TE_M1003_g N_VPWR_c_174_n 0.00500115f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_64 N_TE_c_42_n N_Z_c_208_n 5.4457e-19 $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_65 N_TE_c_44_n N_Z_c_209_n 0.00568018f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_66 N_TE_M1004_g N_VGND_c_243_n 0.00500115f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_67 N_TE_M1004_g N_VGND_c_244_n 0.00341689f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_68 N_TE_M1004_g N_VGND_c_245_n 0.00891715f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_69 N_TE_c_42_n N_VGND_c_245_n 4.05591e-19 $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_70 N_TE_c_44_n N_VGND_c_245_n 0.0202143f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_80_n N_A_c_145_n 0.00101466f $X=0.715 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_27_47#_c_82_n N_A_c_145_n 9.97532e-19 $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_27_47#_M1002_g N_A_M1001_g 0.0405843f $X=1.305 $Y=1.985 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_86_n N_A_M1001_g 5.41511e-19 $X=0.715 $Y=1.98 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_82_n N_A_M1001_g 0.00181599f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_82_n N_A_c_147_n 3.03521e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_83_n N_A_c_147_n 0.0165902f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_86_n N_VPWR_M1003_d 0.0125059f $X=0.715 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_27_47#_c_82_n N_VPWR_M1003_d 0.0117838f $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_47#_c_86_n N_VPWR_c_175_n 0.0640151f $X=0.715 $Y=1.98 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_85_n N_VPWR_c_176_n 0.0177719f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_86_n N_VPWR_c_176_n 0.00273399f $X=0.715 $Y=1.98 $X2=0 $Y2=0
cc_83 N_A_27_47#_M1002_g N_VPWR_c_178_n 0.020663f $X=1.305 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_27_47#_M1003_s N_VPWR_c_174_n 0.00229009f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_85 N_A_27_47#_c_85_n N_VPWR_c_174_n 0.00989054f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_86_n N_VPWR_c_174_n 0.00849566f $X=0.715 $Y=1.98 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_86_n A_276_297# 0.00168179f $X=0.715 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_27_47#_c_82_n A_276_297# 0.00374691f $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_27_47#_M1002_g N_Z_c_208_n 0.00331884f $X=1.305 $Y=1.985 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_86_n N_Z_c_208_n 0.0138578f $X=0.715 $Y=1.98 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_82_n N_Z_c_208_n 0.0871139f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_83_n N_Z_c_208_n 0.00204072f $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1002_g Z 0.0035637f $X=1.305 $Y=1.985 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_80_n N_Z_c_209_n 0.0149229f $X=0.715 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_80_n N_VGND_M1004_d 0.00348575f $X=0.715 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_27_47#_c_82_n N_VGND_M1004_d 8.09036e-19 $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_27_47#_M1004_s N_VGND_c_243_n 0.00229009f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_79_n N_VGND_c_243_n 0.00989054f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_80_n N_VGND_c_243_n 0.00850693f $X=0.715 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_79_n N_VGND_c_244_n 0.0177719f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_80_n N_VGND_c_244_n 0.00273399f $X=0.715 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_80_n N_VGND_c_245_n 0.0642171f $X=0.715 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_83_n N_VGND_c_245_n 8.21139e-19 $X=1.365 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_80_n A_204_47# 0.00776184f $X=0.715 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_27_47#_c_82_n A_204_47# 5.40508e-19 $X=1.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A_M1001_g N_VPWR_c_178_n 0.0032157f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_M1001_g N_VPWR_c_179_n 0.00357877f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1001_g N_VPWR_c_174_n 0.00644121f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_109 A N_Z_M1001_d 0.0106786f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A_c_145_n N_Z_c_208_n 0.0105861f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_Z_c_208_n 0.0223753f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_112 A N_Z_c_208_n 0.0671443f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_113 N_A_c_147_n N_Z_c_208_n 0.00813133f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_M1001_g Z 0.0138808f $X=1.82 $Y=1.985 $X2=0 $Y2=0
cc_115 A Z 0.0197866f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_116 N_A_c_145_n N_Z_c_209_n 0.0232454f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_117 A N_Z_c_209_n 0.0216291f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_c_147_n N_Z_c_209_n 0.00374057f $X=2.06 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_145_n N_VGND_c_242_n 0.00357668f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_145_n N_VGND_c_243_n 0.00756576f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_c_145_n N_VGND_c_245_n 0.0051216f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_122 N_VPWR_c_178_n A_276_297# 0.00253851f $X=1.45 $Y=2.52 $X2=-0.19 $Y2=-0.24
cc_123 N_VPWR_c_174_n A_276_297# 0.00826258f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_124 N_VPWR_c_174_n N_Z_M1001_d 0.00217543f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_125 N_VPWR_c_178_n Z 0.020355f $X=1.45 $Y=2.52 $X2=0 $Y2=0
cc_126 N_VPWR_c_179_n Z 0.0356567f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_174_n Z 0.0217421f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_128 A_276_297# N_Z_c_208_n 0.0059103f $X=1.38 $Y=1.485 $X2=1.305 $Y2=1.985
cc_129 A_276_297# Z 0.0044287f $X=1.38 $Y=1.485 $X2=0 $Y2=0
cc_130 N_Z_c_209_n N_VGND_c_242_n 0.0370535f $X=2.03 $Y=0.38 $X2=0 $Y2=0
cc_131 N_Z_M1000_d N_VGND_c_243_n 0.00217517f $X=1.895 $Y=0.235 $X2=0 $Y2=0
cc_132 N_Z_c_209_n N_VGND_c_243_n 0.0219912f $X=2.03 $Y=0.38 $X2=0 $Y2=0
cc_133 N_Z_c_209_n N_VGND_c_245_n 0.0203492f $X=2.03 $Y=0.38 $X2=0 $Y2=0
cc_134 N_Z_c_208_n A_204_47# 7.70016e-19 $X=1.707 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_135 N_Z_c_209_n A_204_47# 0.00781851f $X=2.03 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_136 N_VGND_c_243_n A_204_47# 0.0083052f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
cc_137 N_VGND_c_245_n A_204_47# 0.00969276f $X=1.45 $Y=0.2 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__a32oi_2.spice.SKY130_FD_SC_HD__A32OI_2.pxi
* Created: Thu Aug 27 14:05:45 2020
* 
x_PM_SKY130_FD_SC_HD__A32OI_2%B2 N_B2_c_82_n N_B2_M1006_g N_B2_M1002_g
+ N_B2_c_83_n N_B2_M1016_g N_B2_M1010_g B2 B2 B2 N_B2_c_85_n N_B2_c_86_n
+ PM_SKY130_FD_SC_HD__A32OI_2%B2
x_PM_SKY130_FD_SC_HD__A32OI_2%B1 N_B1_c_132_n N_B1_M1008_g N_B1_M1000_g
+ N_B1_c_134_n N_B1_M1009_g N_B1_M1015_g B1 B1 N_B1_c_137_n
+ PM_SKY130_FD_SC_HD__A32OI_2%B1
x_PM_SKY130_FD_SC_HD__A32OI_2%A1 N_A1_M1011_g N_A1_c_176_n N_A1_c_177_n
+ N_A1_M1012_g N_A1_M1013_g N_A1_M1019_g A1 A1 N_A1_c_181_n N_A1_c_182_n
+ PM_SKY130_FD_SC_HD__A32OI_2%A1
x_PM_SKY130_FD_SC_HD__A32OI_2%A2 N_A2_M1003_g N_A2_M1001_g N_A2_M1005_g
+ N_A2_M1017_g A2 A2 N_A2_c_232_n PM_SKY130_FD_SC_HD__A32OI_2%A2
x_PM_SKY130_FD_SC_HD__A32OI_2%A3 N_A3_M1007_g N_A3_M1004_g N_A3_M1014_g
+ N_A3_M1018_g N_A3_c_278_n A3 A3 A3 N_A3_c_280_n N_A3_c_281_n
+ PM_SKY130_FD_SC_HD__A32OI_2%A3
x_PM_SKY130_FD_SC_HD__A32OI_2%A_27_297# N_A_27_297#_M1002_d N_A_27_297#_M1010_d
+ N_A_27_297#_M1015_s N_A_27_297#_M1013_d N_A_27_297#_M1017_d
+ N_A_27_297#_M1018_d N_A_27_297#_c_322_n N_A_27_297#_c_325_n
+ N_A_27_297#_c_374_p N_A_27_297#_c_352_p N_A_27_297#_c_327_n
+ N_A_27_297#_c_357_p N_A_27_297#_c_376_p N_A_27_297#_c_330_n
+ N_A_27_297#_c_378_p N_A_27_297#_c_336_n N_A_27_297#_c_380_p
+ N_A_27_297#_c_342_n N_A_27_297#_c_346_n N_A_27_297#_c_366_p
+ N_A_27_297#_c_383_p N_A_27_297#_c_334_n N_A_27_297#_c_340_n
+ PM_SKY130_FD_SC_HD__A32OI_2%A_27_297#
x_PM_SKY130_FD_SC_HD__A32OI_2%Y N_Y_M1008_s N_Y_M1012_d N_Y_M1002_s N_Y_M1000_d
+ N_Y_c_403_n N_Y_c_404_n N_Y_c_420_n N_Y_c_448_n N_Y_c_405_n N_Y_c_400_n
+ N_Y_c_414_n N_Y_c_406_n Y Y Y N_Y_c_435_n Y PM_SKY130_FD_SC_HD__A32OI_2%Y
x_PM_SKY130_FD_SC_HD__A32OI_2%VPWR N_VPWR_M1011_s N_VPWR_M1003_s N_VPWR_M1007_s
+ VPWR N_VPWR_c_477_n N_VPWR_c_476_n N_VPWR_c_479_n N_VPWR_c_480_n
+ N_VPWR_c_481_n N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n
+ PM_SKY130_FD_SC_HD__A32OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A32OI_2%A_27_47# N_A_27_47#_M1006_d N_A_27_47#_M1016_d
+ N_A_27_47#_M1009_d N_A_27_47#_c_557_n N_A_27_47#_c_564_n N_A_27_47#_c_568_n
+ N_A_27_47#_c_558_n N_A_27_47#_c_559_n N_A_27_47#_c_560_n
+ PM_SKY130_FD_SC_HD__A32OI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__A32OI_2%VGND N_VGND_M1006_s N_VGND_M1004_s N_VGND_M1014_s
+ N_VGND_c_600_n N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n
+ N_VGND_c_605_n VGND N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n
+ N_VGND_c_609_n PM_SKY130_FD_SC_HD__A32OI_2%VGND
x_PM_SKY130_FD_SC_HD__A32OI_2%A_478_47# N_A_478_47#_M1012_s N_A_478_47#_M1019_s
+ N_A_478_47#_M1005_d N_A_478_47#_c_673_n PM_SKY130_FD_SC_HD__A32OI_2%A_478_47#
x_PM_SKY130_FD_SC_HD__A32OI_2%A_730_47# N_A_730_47#_M1001_s N_A_730_47#_M1004_d
+ N_A_730_47#_c_693_n N_A_730_47#_c_703_n PM_SKY130_FD_SC_HD__A32OI_2%A_730_47#
cc_1 VNB N_B2_c_82_n 0.0219013f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B2_c_83_n 0.0161517f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB B2 6.57328e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_4 VNB N_B2_c_85_n 0.0507873f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_5 VNB N_B2_c_86_n 0.00861916f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.285
cc_6 VNB N_B1_c_132_n 0.0152125f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_7 VNB N_B1_M1000_g 4.65621e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_8 VNB N_B1_c_134_n 0.0181628f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_B1_M1015_g 4.63504e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_10 VNB B1 0.00381609f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_11 VNB N_B1_c_137_n 0.039394f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_12 VNB N_A1_M1011_g 4.62694e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A1_c_176_n 0.032483f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_14 VNB N_A1_c_177_n 0.0119447f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A1_M1012_g 0.0216798f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_16 VNB N_A1_M1013_g 5.28479e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_17 VNB N_A1_M1019_g 0.0179079f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_18 VNB N_A1_c_181_n 0.00220275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_182_n 0.0312744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_M1003_g 5.64201e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_A2_M1001_g 0.0179079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A2_M1005_g 0.0243831f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_23 VNB N_A2_M1017_g 4.63448e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB A2 0.00257508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A2_c_232_n 0.0628616f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.53
cc_26 VNB N_A3_M1007_g 5.21805e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_27 VNB N_A3_M1004_g 0.0254286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A3_M1014_g 0.0236726f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_29 VNB N_A3_c_278_n 0.0315294f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_30 VNB A3 0.00932659f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_31 VNB N_A3_c_280_n 0.0231563f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.18
cc_32 VNB N_A3_c_281_n 0.0298227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_400_n 0.00592398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB Y 0.00204788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB Y 0.00611398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_476_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_557_n 0.00100766f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_38 VNB N_A_27_47#_c_558_n 0.00164082f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_39 VNB N_A_27_47#_c_559_n 0.00248458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_560_n 0.00821998f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_41 VNB N_VGND_c_600_n 0.00464042f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_42 VNB N_VGND_c_601_n 0.0079466f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_43 VNB N_VGND_c_602_n 0.0102695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_603_n 0.0300854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_604_n 0.0902898f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_46 VNB N_VGND_c_605_n 0.00641049f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_47 VNB N_VGND_c_606_n 0.0175798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_607_n 0.0164642f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_49 VNB N_VGND_c_608_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_609_n 0.301036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_478_47#_c_673_n 0.00439769f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_52 VNB N_A_730_47#_c_693_n 0.0102706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_B2_M1002_g 0.0218837f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_54 VPB N_B2_M1010_g 0.0184996f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_55 VPB B2 0.00761713f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_56 VPB N_B2_c_85_n 0.0128453f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_57 VPB N_B1_M1000_g 0.0195714f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_58 VPB N_B1_M1015_g 0.0195344f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_59 VPB N_A1_M1011_g 0.0225271f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_60 VPB N_A1_M1013_g 0.0239754f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_61 VPB N_A1_c_181_n 0.00305119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A2_M1003_g 0.0230808f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_63 VPB N_A2_M1017_g 0.0208864f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_64 VPB A2 0.00293746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A3_M1007_g 0.0223658f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_66 VPB N_A3_M1018_g 0.0266701f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_67 VPB A3 0.0137789f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.16
cc_68 VPB N_A3_c_281_n 0.00786419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_403_n 0.00368711f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_70 VPB N_Y_c_404_n 0.00152513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_Y_c_405_n 0.00277361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Y_c_406_n 0.00127988f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_73 VPB Y 0.00146229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_477_n 0.0170088f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.53
cc_75 VPB N_VPWR_c_476_n 0.0472033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_479_n 0.0553924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_480_n 0.0198069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_481_n 0.0139376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_482_n 0.0120907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_483_n 0.012158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_484_n 0.0169846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 N_B2_c_83_n N_B1_c_132_n 0.0114813f $X=0.89 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_83 N_B2_c_85_n N_B1_M1000_g 0.0294963f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_84 B2 B1 0.0149648f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_85 N_B2_c_85_n B1 0.00190115f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B2_c_83_n N_B1_c_137_n 0.0227063f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_87 B2 N_A_27_297#_M1002_d 0.0108712f $X=0.15 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_88 B2 N_A_27_297#_c_322_n 0.0131226f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_89 B2 N_A_27_297#_c_322_n 5.14459e-19 $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_90 N_B2_c_85_n N_A_27_297#_c_322_n 9.81971e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B2_M1002_g N_A_27_297#_c_325_n 0.0112878f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_92 N_B2_M1010_g N_A_27_297#_c_325_n 0.00940156f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_93 N_B2_M1010_g N_Y_c_403_n 0.0125535f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_94 B2 N_Y_c_403_n 0.00428436f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B2_M1002_g N_Y_c_404_n 3.78062e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_96 B2 N_Y_c_404_n 0.00546013f $X=0.15 $Y=1.445 $X2=0 $Y2=0
cc_97 B2 N_Y_c_404_n 0.013891f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B2_c_85_n N_Y_c_404_n 0.00219557f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B2_M1002_g N_Y_c_414_n 0.00305424f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B2_M1010_g N_Y_c_414_n 0.00266265f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_101 B2 N_Y_c_414_n 0.00118262f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_102 N_B2_M1002_g N_VPWR_c_476_n 0.00617937f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B2_M1010_g N_VPWR_c_476_n 0.00525237f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B2_M1002_g N_VPWR_c_479_n 0.00357877f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B2_M1010_g N_VPWR_c_479_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_106 B2 N_A_27_47#_c_557_n 0.00113678f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B2_c_85_n N_A_27_47#_c_557_n 0.00426518f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B2_c_86_n N_A_27_47#_c_557_n 0.0117085f $X=0.235 $Y=1.285 $X2=0 $Y2=0
cc_109 N_B2_c_82_n N_A_27_47#_c_564_n 0.00991871f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B2_c_83_n N_A_27_47#_c_564_n 0.0115876f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_111 B2 N_A_27_47#_c_564_n 0.0255175f $X=0.61 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B2_c_85_n N_A_27_47#_c_564_n 0.00218981f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B2_c_83_n N_A_27_47#_c_568_n 0.0025227f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B2_c_82_n N_A_27_47#_c_560_n 0.00248939f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B2_c_85_n N_A_27_47#_c_560_n 3.49353e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B2_c_86_n N_A_27_47#_c_560_n 8.89165e-19 $X=0.235 $Y=1.285 $X2=0 $Y2=0
cc_117 N_B2_c_82_n N_VGND_c_600_n 0.00268723f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B2_c_83_n N_VGND_c_600_n 0.00268723f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B2_c_83_n N_VGND_c_604_n 0.00422371f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B2_c_82_n N_VGND_c_606_n 0.00422842f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B2_c_82_n N_VGND_c_609_n 0.00666796f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B2_c_83_n N_VGND_c_609_n 0.00573566f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B1_M1015_g N_A1_M1011_g 0.0205666f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_c_137_n N_A1_c_177_n 0.0205666f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_125 N_B1_M1000_g N_A_27_297#_c_327_n 0.00984328f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_126 N_B1_M1015_g N_A_27_297#_c_327_n 0.00988743f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B1_M1000_g N_Y_c_403_n 0.0125959f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_128 B1 N_Y_c_403_n 0.0283661f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B1_c_137_n N_Y_c_403_n 0.00135177f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_130 N_B1_c_132_n N_Y_c_420_n 0.00265203f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_131 N_B1_c_134_n N_Y_c_420_n 0.0119086f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_132 B1 N_Y_c_420_n 0.0161131f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B1_c_137_n N_Y_c_420_n 0.00214152f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_134 N_B1_M1015_g N_Y_c_405_n 0.0137013f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 B1 N_Y_c_405_n 0.00844795f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_136 B1 N_Y_c_406_n 0.0139492f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_137 N_B1_c_137_n N_Y_c_406_n 0.00210302f $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_138 N_B1_c_134_n Y 0.0139125f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_139 B1 Y 0.0130281f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_140 N_B1_M1000_g N_VPWR_c_476_n 0.00525237f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B1_M1015_g N_VPWR_c_476_n 0.00525237f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B1_M1000_g N_VPWR_c_479_n 0.00357877f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B1_M1015_g N_VPWR_c_479_n 0.00357877f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_144 B1 N_A_27_47#_c_558_n 0.0102352f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_145 N_B1_c_137_n N_A_27_47#_c_558_n 2.30684e-19 $X=1.73 $Y=1.135 $X2=0 $Y2=0
cc_146 N_B1_c_132_n N_A_27_47#_c_559_n 0.00956005f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_147 N_B1_c_134_n N_A_27_47#_c_559_n 0.00801257f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_148 B1 N_A_27_47#_c_559_n 0.00347347f $X=1.53 $Y=1.105 $X2=0 $Y2=0
cc_149 N_B1_c_132_n N_VGND_c_604_n 0.00366111f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_150 N_B1_c_134_n N_VGND_c_604_n 0.00366111f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_151 N_B1_c_132_n N_VGND_c_609_n 0.00526729f $X=1.31 $Y=0.975 $X2=0 $Y2=0
cc_152 N_B1_c_134_n N_VGND_c_609_n 0.00656615f $X=1.73 $Y=0.975 $X2=0 $Y2=0
cc_153 N_A1_M1013_g N_A2_M1003_g 0.025021f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A1_c_181_n N_A2_M1003_g 0.00350407f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A1_M1019_g N_A2_M1001_g 0.014117f $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A1_c_181_n A2 0.0213892f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_181_n N_A2_c_232_n 0.00104004f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A1_c_182_n N_A2_c_232_n 0.0322132f $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A1_c_181_n N_A_27_297#_M1013_d 0.00231502f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_M1011_g N_A_27_297#_c_330_n 0.0136819f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A1_c_176_n N_A_27_297#_c_330_n 0.00394077f $X=2.65 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_M1013_g N_A_27_297#_c_330_n 0.0124955f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_c_181_n N_A_27_297#_c_330_n 0.0345657f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A1_c_181_n N_A_27_297#_c_334_n 0.0029123f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_c_177_n N_Y_c_400_n 0.0138351f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_M1012_g N_Y_c_400_n 0.0110467f $X=2.725 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A1_M1019_g N_Y_c_400_n 0.00391909f $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A1_c_181_n N_Y_c_400_n 0.0339521f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A1_c_182_n N_Y_c_400_n 0.00237042f $X=3.145 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A1_M1011_g N_Y_c_435_n 0.00694622f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_c_181_n N_Y_c_435_n 0.0115461f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_M1011_g Y 0.00376314f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A1_c_177_n Y 0.0123986f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A1_M1012_g Y 0.00510972f $X=2.725 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A1_c_181_n Y 0.0233162f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A1_c_181_n N_VPWR_M1011_s 0.0115227f $X=3.055 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A1_M1011_g N_VPWR_c_476_n 0.00710026f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_178 N_A1_M1013_g N_VPWR_c_476_n 0.00715993f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A1_M1011_g N_VPWR_c_479_n 0.00425094f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_180 N_A1_M1011_g N_VPWR_c_480_n 0.00927673f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A1_M1013_g N_VPWR_c_480_n 0.00779316f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_182 N_A1_M1013_g N_VPWR_c_481_n 0.00396755f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A1_M1013_g N_VPWR_c_482_n 5.53705e-19 $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A1_M1012_g N_VGND_c_604_n 0.00366111f $X=2.725 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A1_M1019_g N_VGND_c_604_n 0.00366111f $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A1_M1012_g N_VGND_c_609_n 0.00656615f $X=2.725 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A1_M1019_g N_VGND_c_609_n 0.0052918f $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A1_M1012_g N_A_478_47#_c_673_n 0.00801257f $X=2.725 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A1_M1019_g N_A_478_47#_c_673_n 0.00956283f $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A1_c_181_n N_A_478_47#_c_673_n 0.00308926f $X=3.055 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A1_M1019_g N_A_730_47#_c_693_n 5.33998e-19 $X=3.145 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A2_M1017_g N_A3_M1007_g 0.027506f $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_193 A2 N_A3_c_278_n 0.00446129f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_194 N_A2_c_232_n N_A3_c_278_n 0.0177431f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A2_M1017_g A3 2.92151e-19 $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_196 A2 A3 0.0379773f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A2_c_232_n A3 2.01765e-19 $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_198 A2 N_A_27_297#_M1017_d 0.00227451f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A2_M1003_g N_A_27_297#_c_336_n 0.0152317f $X=3.505 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A2_M1017_g N_A_27_297#_c_336_n 0.0113632f $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_201 A2 N_A_27_297#_c_336_n 0.0291917f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A2_c_232_n N_A_27_297#_c_336_n 0.00272599f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_203 A2 N_A_27_297#_c_340_n 0.00732487f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A2_M1001_g N_Y_c_400_n 5.33998e-19 $X=3.575 $Y=0.56 $X2=0 $Y2=0
cc_205 A2 N_VPWR_M1003_s 0.00985749f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_206 N_A2_M1003_g N_VPWR_c_476_n 0.00402785f $X=3.505 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1017_g N_VPWR_c_476_n 0.00396795f $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_M1003_g N_VPWR_c_481_n 0.00198377f $X=3.505 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A2_M1003_g N_VPWR_c_482_n 0.00815414f $X=3.505 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1017_g N_VPWR_c_482_n 0.00785119f $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_M1017_g N_VPWR_c_483_n 0.00198377f $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A2_M1017_g N_VPWR_c_484_n 4.2177e-19 $X=4.265 $Y=1.985 $X2=0 $Y2=0
cc_213 N_A2_M1005_g N_VGND_c_601_n 0.00296976f $X=3.995 $Y=0.56 $X2=0 $Y2=0
cc_214 N_A2_M1001_g N_VGND_c_604_n 0.00366111f $X=3.575 $Y=0.56 $X2=0 $Y2=0
cc_215 N_A2_M1005_g N_VGND_c_604_n 0.00366111f $X=3.995 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A2_M1001_g N_VGND_c_609_n 0.0052918f $X=3.575 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A2_M1005_g N_VGND_c_609_n 0.00656615f $X=3.995 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A2_M1001_g N_A_478_47#_c_673_n 0.0115259f $X=3.575 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A2_M1005_g N_A_478_47#_c_673_n 0.00789149f $X=3.995 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A2_c_232_n N_A_478_47#_c_673_n 0.00126404f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_M1001_g N_A_730_47#_c_693_n 0.0046906f $X=3.575 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A2_M1005_g N_A_730_47#_c_693_n 0.0110355f $X=3.995 $Y=0.56 $X2=0 $Y2=0
cc_223 A2 N_A_730_47#_c_693_n 0.0379447f $X=4.29 $Y=1.105 $X2=0 $Y2=0
cc_224 N_A2_c_232_n N_A_730_47#_c_693_n 0.00978572f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_225 A3 N_A_27_297#_M1018_d 0.00417024f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_226 N_A3_M1007_g N_A_27_297#_c_342_n 0.0143549f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A3_M1018_g N_A_27_297#_c_342_n 0.0119845f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A3_c_278_n N_A_27_297#_c_342_n 0.00169285f $X=5.065 $Y=1.16 $X2=0 $Y2=0
cc_229 A3 N_A_27_297#_c_342_n 0.0395745f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_230 A3 N_A_27_297#_c_346_n 0.0143851f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_231 N_A3_c_281_n N_A_27_297#_c_346_n 6.66445e-19 $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_232 A3 N_VPWR_M1007_s 0.0102386f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A3_M1018_g N_VPWR_c_477_n 0.00424386f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A3_M1007_g N_VPWR_c_476_n 0.00481068f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A3_M1018_g N_VPWR_c_476_n 0.00572537f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A3_M1007_g N_VPWR_c_482_n 5.35972e-19 $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A3_M1007_g N_VPWR_c_483_n 0.00283396f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_238 N_A3_M1007_g N_VPWR_c_484_n 0.00238518f $X=4.69 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A3_M1018_g N_VPWR_c_484_n 0.00408381f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A3_M1004_g N_VGND_c_601_n 0.00342139f $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_241 N_A3_M1004_g N_VGND_c_603_n 4.59439e-19 $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A3_M1014_g N_VGND_c_603_n 0.0131032f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_243 A3 N_VGND_c_603_n 0.0210599f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_244 N_A3_c_281_n N_VGND_c_603_n 0.00644411f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A3_M1004_g N_VGND_c_607_n 0.00424476f $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A3_M1014_g N_VGND_c_607_n 0.00486043f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_247 N_A3_M1004_g N_VGND_c_609_n 0.00712125f $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A3_M1014_g N_VGND_c_609_n 0.00852643f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A3_M1004_g N_A_730_47#_c_693_n 0.0122117f $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A3_c_278_n N_A_730_47#_c_693_n 0.00867145f $X=5.065 $Y=1.16 $X2=0 $Y2=0
cc_251 A3 N_A_730_47#_c_693_n 0.0339639f $X=5.67 $Y=1.105 $X2=0 $Y2=0
cc_252 N_A3_c_280_n N_A_730_47#_c_693_n 0.00423012f $X=5.435 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A3_M1004_g N_A_730_47#_c_703_n 0.00881054f $X=4.99 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_27_297#_c_325_n N_Y_M1002_s 0.00312348f $X=1.015 $Y=2.38 $X2=0.47
+ $Y2=0.56
cc_255 N_A_27_297#_c_327_n N_Y_M1000_d 0.00312348f $X=1.855 $Y=2.38 $X2=0.47
+ $Y2=1.325
cc_256 N_A_27_297#_M1010_d N_Y_c_403_n 0.00165831f $X=0.965 $Y=1.485 $X2=0.61
+ $Y2=1.105
cc_257 N_A_27_297#_c_325_n N_Y_c_403_n 0.00259534f $X=1.015 $Y=2.38 $X2=0.61
+ $Y2=1.105
cc_258 N_A_27_297#_c_352_p N_Y_c_403_n 0.0126766f $X=1.1 $Y=1.96 $X2=0.61
+ $Y2=1.105
cc_259 N_A_27_297#_c_327_n N_Y_c_403_n 0.00321995f $X=1.855 $Y=2.38 $X2=0.61
+ $Y2=1.105
cc_260 N_A_27_297#_c_327_n N_Y_c_448_n 0.0118729f $X=1.855 $Y=2.38 $X2=0.66
+ $Y2=1.16
cc_261 N_A_27_297#_M1015_s N_Y_c_405_n 0.00108428f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_262 N_A_27_297#_c_327_n N_Y_c_405_n 0.00321995f $X=1.855 $Y=2.38 $X2=0 $Y2=0
cc_263 N_A_27_297#_c_357_p N_Y_c_405_n 0.00833331f $X=1.94 $Y=2.085 $X2=0 $Y2=0
cc_264 N_A_27_297#_c_325_n N_Y_c_414_n 0.0155384f $X=1.015 $Y=2.38 $X2=0 $Y2=0
cc_265 N_A_27_297#_M1015_s N_Y_c_435_n 5.86511e-19 $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_357_p N_Y_c_435_n 0.00477333f $X=1.94 $Y=2.085 $X2=0 $Y2=0
cc_267 N_A_27_297#_c_330_n N_Y_c_435_n 0.00515916f $X=3.18 $Y=2 $X2=0 $Y2=0
cc_268 N_A_27_297#_c_330_n N_VPWR_M1011_s 0.0195044f $X=3.18 $Y=2 $X2=0.47
+ $Y2=0.995
cc_269 N_A_27_297#_c_336_n N_VPWR_M1003_s 0.0146717f $X=4.39 $Y=2 $X2=0.47
+ $Y2=0.56
cc_270 N_A_27_297#_c_342_n N_VPWR_M1007_s 0.0155134f $X=5.635 $Y=2 $X2=0.47
+ $Y2=0.56
cc_271 N_A_27_297#_c_342_n N_VPWR_c_477_n 0.00292742f $X=5.635 $Y=2 $X2=0.235
+ $Y2=1.53
cc_272 N_A_27_297#_c_366_p N_VPWR_c_477_n 0.0115924f $X=5.72 $Y=2.3 $X2=0.235
+ $Y2=1.53
cc_273 N_A_27_297#_M1002_d N_VPWR_c_476_n 0.00348186f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_M1010_d N_VPWR_c_476_n 0.0021521f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_M1015_s N_VPWR_c_476_n 0.00233082f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_M1013_d N_VPWR_c_476_n 0.00284382f $X=3.13 $Y=1.485 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_M1017_d N_VPWR_c_476_n 0.00255187f $X=4.34 $Y=1.485 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_M1018_d N_VPWR_c_476_n 0.00368727f $X=5.585 $Y=1.485 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_c_325_n N_VPWR_c_476_n 0.0234424f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_374_p N_VPWR_c_476_n 0.00654447f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_c_327_n N_VPWR_c_476_n 0.0234424f $X=1.855 $Y=2.38 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_376_p N_VPWR_c_476_n 0.00654444f $X=1.94 $Y=2.295 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_c_330_n N_VPWR_c_476_n 0.0158571f $X=3.18 $Y=2 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_378_p N_VPWR_c_476_n 0.00646745f $X=3.265 $Y=2.3 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_336_n N_VPWR_c_476_n 0.013349f $X=4.39 $Y=2 $X2=0 $Y2=0
cc_286 N_A_27_297#_c_380_p N_VPWR_c_476_n 0.00646224f $X=4.475 $Y=2.3 $X2=0
+ $Y2=0
cc_287 N_A_27_297#_c_342_n N_VPWR_c_476_n 0.0135005f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_366_p N_VPWR_c_476_n 0.00646745f $X=5.72 $Y=2.3 $X2=0 $Y2=0
cc_289 N_A_27_297#_c_383_p N_VPWR_c_476_n 0.00654447f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_290 N_A_27_297#_c_325_n N_VPWR_c_479_n 0.0358391f $X=1.015 $Y=2.38 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_c_374_p N_VPWR_c_479_n 0.0116982f $X=0.345 $Y=2.38 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_c_327_n N_VPWR_c_479_n 0.0358391f $X=1.855 $Y=2.38 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_c_376_p N_VPWR_c_479_n 0.0114548f $X=1.94 $Y=2.295 $X2=0
+ $Y2=0
cc_294 N_A_27_297#_c_330_n N_VPWR_c_479_n 0.00336774f $X=3.18 $Y=2 $X2=0 $Y2=0
cc_295 N_A_27_297#_c_383_p N_VPWR_c_479_n 0.0114548f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_296 N_A_27_297#_c_330_n N_VPWR_c_480_n 0.0486454f $X=3.18 $Y=2 $X2=0 $Y2=0
cc_297 N_A_27_297#_c_330_n N_VPWR_c_481_n 0.00277357f $X=3.18 $Y=2 $X2=0 $Y2=0
cc_298 N_A_27_297#_c_378_p N_VPWR_c_481_n 0.0115924f $X=3.265 $Y=2.3 $X2=0 $Y2=0
cc_299 N_A_27_297#_c_336_n N_VPWR_c_481_n 0.0021306f $X=4.39 $Y=2 $X2=0 $Y2=0
cc_300 N_A_27_297#_c_378_p N_VPWR_c_482_n 0.01446f $X=3.265 $Y=2.3 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_336_n N_VPWR_c_482_n 0.0418204f $X=4.39 $Y=2 $X2=0 $Y2=0
cc_302 N_A_27_297#_c_336_n N_VPWR_c_483_n 0.00162812f $X=4.39 $Y=2 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_380_p N_VPWR_c_483_n 0.0115577f $X=4.475 $Y=2.3 $X2=0 $Y2=0
cc_304 N_A_27_297#_c_342_n N_VPWR_c_483_n 0.00216795f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_305 N_A_27_297#_c_342_n N_VPWR_c_484_n 0.0421947f $X=5.635 $Y=2 $X2=0 $Y2=0
cc_306 N_Y_M1002_s N_VPWR_c_476_n 0.00216833f $X=0.545 $Y=1.485 $X2=0 $Y2=0
cc_307 N_Y_M1000_d N_VPWR_c_476_n 0.00216833f $X=1.385 $Y=1.485 $X2=0 $Y2=0
cc_308 N_Y_c_420_n N_A_27_47#_M1009_d 0.0030652f $X=1.965 $Y=0.74 $X2=0 $Y2=0
cc_309 Y N_A_27_47#_M1009_d 0.00187356f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_310 Y N_A_27_47#_M1009_d 7.83609e-19 $X=2.075 $Y=0.85 $X2=0 $Y2=0
cc_311 N_Y_c_403_n N_A_27_47#_c_564_n 0.00430475f $X=1.435 $Y=1.54 $X2=0 $Y2=0
cc_312 N_Y_c_403_n N_A_27_47#_c_558_n 8.97464e-19 $X=1.435 $Y=1.54 $X2=0 $Y2=0
cc_313 N_Y_M1008_s N_A_27_47#_c_559_n 0.00322663f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_314 N_Y_c_420_n N_A_27_47#_c_559_n 0.026632f $X=1.965 $Y=0.74 $X2=0 $Y2=0
cc_315 Y N_A_27_47#_c_559_n 0.0106311f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_316 N_Y_c_400_n N_VGND_c_604_n 0.00297094f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_317 Y N_VGND_c_604_n 0.00126693f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_318 N_Y_M1008_s N_VGND_c_609_n 0.00219239f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_319 N_Y_M1012_d N_VGND_c_609_n 0.00219239f $X=2.8 $Y=0.235 $X2=0 $Y2=0
cc_320 N_Y_c_400_n N_VGND_c_609_n 0.00622316f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_321 Y N_VGND_c_609_n 0.00233732f $X=1.99 $Y=0.765 $X2=0 $Y2=0
cc_322 N_Y_c_400_n N_A_478_47#_M1012_s 0.00498049f $X=2.935 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_323 N_Y_M1012_d N_A_478_47#_c_673_n 0.00324009f $X=2.8 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_c_400_n N_A_478_47#_c_673_n 0.0355575f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_325 N_Y_c_400_n N_A_730_47#_c_693_n 0.00499003f $X=2.935 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_564_n N_VGND_M1006_s 0.00312505f $X=1.015 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_327 N_A_27_47#_c_564_n N_VGND_c_600_n 0.012179f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_328 N_A_27_47#_c_564_n N_VGND_c_604_n 0.00203142f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_329 N_A_27_47#_c_568_n N_VGND_c_604_n 0.0119274f $X=1.1 $Y=0.465 $X2=0 $Y2=0
cc_330 N_A_27_47#_c_559_n N_VGND_c_604_n 0.0416716f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_331 N_A_27_47#_c_564_n N_VGND_c_606_n 0.0020451f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_560_n N_VGND_c_606_n 0.0161209f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_333 N_A_27_47#_M1006_d N_VGND_c_609_n 0.00211564f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_M1016_d N_VGND_c_609_n 0.00217541f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_27_47#_M1009_d N_VGND_c_609_n 0.00211652f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_564_n N_VGND_c_609_n 0.00878868f $X=1.015 $Y=0.8 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_568_n N_VGND_c_609_n 0.00909294f $X=1.1 $Y=0.465 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_559_n N_VGND_c_609_n 0.0322604f $X=1.94 $Y=0.38 $X2=0 $Y2=0
cc_339 N_A_27_47#_c_560_n N_VGND_c_609_n 0.0119347f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_559_n N_A_478_47#_c_673_n 0.0125258f $X=1.94 $Y=0.38 $X2=0
+ $Y2=0
cc_341 N_VGND_c_609_n N_A_478_47#_M1012_s 0.00211652f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_342 N_VGND_c_609_n N_A_478_47#_M1019_s 0.00225735f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_609_n N_A_478_47#_M1005_d 0.00211652f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_601_n N_A_478_47#_c_673_n 0.0140123f $X=4.725 $Y=0.38 $X2=0
+ $Y2=0
cc_345 N_VGND_c_604_n N_A_478_47#_c_673_n 0.0911064f $X=4.555 $Y=0 $X2=0 $Y2=0
cc_346 N_VGND_c_609_n N_A_478_47#_c_673_n 0.0703441f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_609_n N_A_730_47#_M1001_s 0.00219239f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_348 N_VGND_c_609_n N_A_730_47#_M1004_d 0.00457f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_M1004_s N_A_730_47#_c_693_n 0.00713746f $X=4.6 $Y=0.235 $X2=0
+ $Y2=0
cc_350 N_VGND_c_601_n N_A_730_47#_c_693_n 0.023169f $X=4.725 $Y=0.38 $X2=0 $Y2=0
cc_351 N_VGND_c_604_n N_A_730_47#_c_693_n 0.00337127f $X=4.555 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_607_n N_A_730_47#_c_693_n 0.00260098f $X=5.56 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_609_n N_A_730_47#_c_693_n 0.0121901f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_607_n N_A_730_47#_c_703_n 0.0180353f $X=5.56 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_609_n N_A_730_47#_c_703_n 0.0123348f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_356 N_A_478_47#_c_673_n N_A_730_47#_M1001_s 0.0031669f $X=4.205 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_357 N_A_478_47#_M1005_d N_A_730_47#_c_693_n 0.0049097f $X=4.07 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_A_478_47#_c_673_n N_A_730_47#_c_693_n 0.0390874f $X=4.205 $Y=0.38 $X2=0
+ $Y2=0

* NGSPICE file created from sky130_fd_sc_hd__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_193_47# a_27_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.664e+11p pd=1.8e+06u as=1.2548e+12p ps=1.26e+07u
M1001 a_644_413# a_193_47# a_560_47# VPB phighvt w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_560_47# a_27_47# a_465_369# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.915e+11p ps=1.93e+06u
M1003 VGND D a_299_47# VNB nshort w=420000u l=150000u
+  ad=7.0325e+11p pd=7.85e+06u as=1.092e+11p ps=1.36e+06u
M1004 Q a_711_307# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1005 VGND a_711_307# a_657_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.32e+11p ps=1.49e+06u
M1006 a_711_307# a_560_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
M1007 a_465_47# a_299_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.32e+11p pd=1.49e+06u as=0p ps=0u
M1008 VGND a_711_307# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Q a_711_307# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.05e+11p pd=2.61e+06u as=0p ps=0u
M1010 VPWR GATE a_27_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1011 VPWR a_711_307# a_644_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_193_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1013 a_465_369# a_299_47# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_711_307# Q VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND RESET_B a_940_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1016 VPWR D a_299_47# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.664e+11p ps=1.8e+06u
M1017 a_560_47# a_193_47# a_465_47# VNB nshort w=360000u l=150000u
+  ad=1.206e+11p pd=1.39e+06u as=0p ps=0u
M1018 a_657_47# a_27_47# a_560_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_940_47# a_560_47# a_711_307# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1020 VGND GATE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1021 VPWR RESET_B a_711_307# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_hd__inv_16.pxi.spice
* Created: Tue Sep  1 19:09:49 2020
* 
x_PM_SKY130_FD_SC_HD__INV_16%A N_A_c_106_n N_A_M1005_g N_A_M1000_g N_A_c_107_n
+ N_A_M1007_g N_A_M1001_g N_A_c_108_n N_A_M1008_g N_A_M1002_g N_A_c_109_n
+ N_A_M1011_g N_A_M1003_g N_A_c_110_n N_A_M1012_g N_A_M1004_g N_A_c_111_n
+ N_A_M1013_g N_A_M1006_g N_A_c_112_n N_A_M1016_g N_A_M1009_g N_A_c_113_n
+ N_A_M1018_g N_A_M1010_g N_A_c_114_n N_A_M1019_g N_A_M1014_g N_A_c_115_n
+ N_A_M1022_g N_A_M1015_g N_A_c_116_n N_A_M1023_g N_A_M1017_g N_A_c_117_n
+ N_A_M1024_g N_A_M1020_g N_A_c_118_n N_A_M1026_g N_A_M1021_g N_A_c_119_n
+ N_A_M1027_g N_A_M1025_g N_A_c_120_n N_A_M1028_g N_A_M1030_g N_A_c_121_n
+ N_A_M1029_g N_A_M1031_g A A A A A A N_A_c_122_n N_A_c_123_n
+ PM_SKY130_FD_SC_HD__INV_16%A
x_PM_SKY130_FD_SC_HD__INV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_M1025_d
+ N_VPWR_M1031_d N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n
+ N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n VPWR
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_419_n
+ PM_SKY130_FD_SC_HD__INV_16%VPWR
x_PM_SKY130_FD_SC_HD__INV_16%Y N_Y_M1005_d N_Y_M1008_d N_Y_M1012_d N_Y_M1016_d
+ N_Y_M1019_d N_Y_M1023_d N_Y_M1026_d N_Y_M1028_d N_Y_M1000_s N_Y_M1002_s
+ N_Y_M1004_s N_Y_M1009_s N_Y_M1014_s N_Y_M1017_s N_Y_M1021_s N_Y_M1030_s
+ N_Y_c_549_n N_Y_c_552_n N_Y_c_556_n N_Y_c_535_n N_Y_c_536_n N_Y_c_567_n
+ N_Y_c_571_n N_Y_c_575_n N_Y_c_537_n N_Y_c_583_n N_Y_c_587_n N_Y_c_591_n
+ N_Y_c_538_n N_Y_c_599_n N_Y_c_603_n N_Y_c_607_n N_Y_c_539_n N_Y_c_615_n
+ N_Y_c_619_n N_Y_c_623_n N_Y_c_540_n N_Y_c_631_n N_Y_c_635_n N_Y_c_639_n
+ N_Y_c_541_n N_Y_c_647_n N_Y_c_651_n N_Y_c_655_n N_Y_c_542_n N_Y_c_662_n
+ N_Y_c_665_n N_Y_c_668_n N_Y_c_543_n N_Y_c_675_n N_Y_c_544_n N_Y_c_683_n
+ N_Y_c_545_n N_Y_c_691_n N_Y_c_546_n N_Y_c_699_n N_Y_c_547_n N_Y_c_707_n
+ N_Y_c_548_n N_Y_c_714_n N_Y_c_717_n Y Y PM_SKY130_FD_SC_HD__INV_16%Y
x_PM_SKY130_FD_SC_HD__INV_16%VGND N_VGND_M1005_s N_VGND_M1007_s N_VGND_M1011_s
+ N_VGND_M1013_s N_VGND_M1018_s N_VGND_M1022_s N_VGND_M1024_s N_VGND_M1027_s
+ N_VGND_M1029_s N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n VGND
+ N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n
+ PM_SKY130_FD_SC_HD__INV_16%VGND
cc_1 VNB N_A_c_106_n 0.0218814f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=0.995
cc_2 VNB N_A_c_107_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_A_c_108_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.375 $Y2=0.995
cc_4 VNB N_A_c_109_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=0.995
cc_5 VNB N_A_c_110_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=0.995
cc_6 VNB N_A_c_111_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.995
cc_7 VNB N_A_c_112_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.055 $Y2=0.995
cc_8 VNB N_A_c_113_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.475 $Y2=0.995
cc_9 VNB N_A_c_114_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_10 VNB N_A_c_115_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=4.315 $Y2=0.995
cc_11 VNB N_A_c_116_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=4.735 $Y2=0.995
cc_12 VNB N_A_c_117_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=5.155 $Y2=0.995
cc_13 VNB N_A_c_118_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=5.575 $Y2=0.995
cc_14 VNB N_A_c_119_n 0.0157766f $X=-0.19 $Y=-0.24 $X2=5.995 $Y2=0.995
cc_15 VNB N_A_c_120_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=6.415 $Y2=0.995
cc_16 VNB N_A_c_121_n 0.0214956f $X=-0.19 $Y=-0.24 $X2=6.835 $Y2=0.995
cc_17 VNB N_A_c_122_n 0.0109395f $X=-0.19 $Y=-0.24 $X2=5.36 $Y2=1.16
cc_18 VNB N_A_c_123_n 0.293671f $X=-0.19 $Y=-0.24 $X2=6.835 $Y2=1.16
cc_19 VNB N_VPWR_c_419_n 0.30769f $X=-0.19 $Y=-0.24 $X2=4.285 $Y2=1.105
cc_20 VNB N_Y_c_535_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_21 VNB N_Y_c_536_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.56
cc_22 VNB N_Y_c_537_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=4.315 $Y2=1.985
cc_23 VNB N_Y_c_538_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=5.155 $Y2=1.325
cc_24 VNB N_Y_c_539_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=5.995 $Y2=0.56
cc_25 VNB N_Y_c_540_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_541_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=3.825 $Y2=1.105
cc_27 VNB N_Y_c_542_n 0.00325491f $X=-0.19 $Y=-0.24 $X2=0.535 $Y2=1.16
cc_28 VNB N_Y_c_543_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=5.36 $Y2=1.16
cc_29 VNB N_Y_c_544_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=6.415 $Y2=1.16
cc_30 VNB N_Y_c_545_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.195
cc_31 VNB N_Y_c_546_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.195
cc_32 VNB N_Y_c_547_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.195
cc_33 VNB N_Y_c_548_n 0.0032479f $X=-0.19 $Y=-0.24 $X2=4.37 $Y2=1.195
cc_34 VNB N_VGND_c_823_n 0.0123634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_824_n 0.0293904f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=0.56
cc_36 VNB N_VGND_c_825_n 0.017296f $X=-0.19 $Y=-0.24 $X2=2.215 $Y2=1.325
cc_37 VNB N_VGND_c_826_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=0.995
cc_38 VNB N_VGND_c_827_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.635 $Y2=1.985
cc_39 VNB N_VGND_c_828_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.055 $Y2=0.56
cc_40 VNB N_VGND_c_829_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.055 $Y2=1.985
cc_41 VNB N_VGND_c_830_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.475 $Y2=0.56
cc_42 VNB N_VGND_c_831_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.475 $Y2=1.985
cc_43 VNB N_VGND_c_832_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.56
cc_44 VNB N_VGND_c_833_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=1.985
cc_45 VNB N_VGND_c_834_n 0.0122977f $X=-0.19 $Y=-0.24 $X2=4.315 $Y2=0.995
cc_46 VNB N_VGND_c_835_n 0.0126159f $X=-0.19 $Y=-0.24 $X2=4.315 $Y2=0.56
cc_47 VNB N_VGND_c_836_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=4.315 $Y2=1.985
cc_48 VNB N_VGND_c_837_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_838_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=4.735 $Y2=0.56
cc_50 VNB N_VGND_c_839_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=4.735 $Y2=0.56
cc_51 VNB N_VGND_c_840_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=4.735 $Y2=1.985
cc_52 VNB N_VGND_c_841_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=4.735 $Y2=1.985
cc_53 VNB N_VGND_c_842_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_843_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=5.155 $Y2=0.995
cc_55 VNB N_VGND_c_844_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=5.155 $Y2=0.56
cc_56 VNB N_VGND_c_845_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=5.155 $Y2=1.325
cc_57 VNB N_VGND_c_846_n 0.017296f $X=-0.19 $Y=-0.24 $X2=6.415 $Y2=0.56
cc_58 VNB N_VGND_c_847_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=6.835 $Y2=1.325
cc_59 VNB N_VGND_c_848_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_849_n 0.358694f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_61 VPB N_A_M1000_g 0.0259842f $X=-0.19 $Y=1.305 $X2=0.535 $Y2=1.985
cc_62 VPB N_A_M1001_g 0.0185065f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_63 VPB N_A_M1002_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.375 $Y2=1.985
cc_64 VPB N_A_M1003_g 0.0185065f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.985
cc_65 VPB N_A_M1004_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.215 $Y2=1.985
cc_66 VPB N_A_M1006_g 0.0185065f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=1.985
cc_67 VPB N_A_M1009_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.055 $Y2=1.985
cc_68 VPB N_A_M1010_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.475 $Y2=1.985
cc_69 VPB N_A_M1014_g 0.0185065f $X=-0.19 $Y=1.305 $X2=3.895 $Y2=1.985
cc_70 VPB N_A_M1015_g 0.0185065f $X=-0.19 $Y=1.305 $X2=4.315 $Y2=1.985
cc_71 VPB N_A_M1017_g 0.0185065f $X=-0.19 $Y=1.305 $X2=4.735 $Y2=1.985
cc_72 VPB N_A_M1020_g 0.0185065f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=1.985
cc_73 VPB N_A_M1021_g 0.0185065f $X=-0.19 $Y=1.305 $X2=5.575 $Y2=1.985
cc_74 VPB N_A_M1025_g 0.0184947f $X=-0.19 $Y=1.305 $X2=5.995 $Y2=1.985
cc_75 VPB N_A_M1030_g 0.0178241f $X=-0.19 $Y=1.305 $X2=6.415 $Y2=1.985
cc_76 VPB N_A_M1031_g 0.0253019f $X=-0.19 $Y=1.305 $X2=6.835 $Y2=1.985
cc_77 VPB N_A_c_122_n 0.00197941f $X=-0.19 $Y=1.305 $X2=5.36 $Y2=1.16
cc_78 VPB N_A_c_123_n 0.0605983f $X=-0.19 $Y=1.305 $X2=6.835 $Y2=1.16
cc_79 VPB N_VPWR_c_420_n 0.0125908f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_421_n 0.00562374f $X=-0.19 $Y=1.305 $X2=2.215 $Y2=0.56
cc_81 VPB N_VPWR_c_422_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.215 $Y2=1.985
cc_82 VPB N_VPWR_c_423_n 0.00358901f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=0.56
cc_83 VPB N_VPWR_c_424_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_425_n 0.00358901f $X=-0.19 $Y=1.305 $X2=3.055 $Y2=1.325
cc_85 VPB N_VPWR_c_426_n 0.00358901f $X=-0.19 $Y=1.305 $X2=3.475 $Y2=0.995
cc_86 VPB N_VPWR_c_427_n 0.00358901f $X=-0.19 $Y=1.305 $X2=3.475 $Y2=1.985
cc_87 VPB N_VPWR_c_428_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_429_n 0.00358901f $X=-0.19 $Y=1.305 $X2=3.895 $Y2=1.325
cc_89 VPB N_VPWR_c_430_n 0.00358901f $X=-0.19 $Y=1.305 $X2=4.315 $Y2=0.995
cc_90 VPB N_VPWR_c_431_n 0.0122718f $X=-0.19 $Y=1.305 $X2=4.315 $Y2=0.56
cc_91 VPB N_VPWR_c_432_n 0.00438892f $X=-0.19 $Y=1.305 $X2=4.315 $Y2=1.985
cc_92 VPB N_VPWR_c_433_n 0.017949f $X=-0.19 $Y=1.305 $X2=4.735 $Y2=0.995
cc_93 VPB N_VPWR_c_434_n 0.00323736f $X=-0.19 $Y=1.305 $X2=4.735 $Y2=0.56
cc_94 VPB N_VPWR_c_435_n 0.017949f $X=-0.19 $Y=1.305 $X2=4.735 $Y2=1.325
cc_95 VPB N_VPWR_c_436_n 0.00323736f $X=-0.19 $Y=1.305 $X2=4.735 $Y2=1.985
cc_96 VPB N_VPWR_c_437_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_438_n 0.00323736f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=0.995
cc_98 VPB N_VPWR_c_439_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=0.56
cc_99 VPB N_VPWR_c_440_n 0.00323736f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=0.56
cc_100 VPB N_VPWR_c_441_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=1.985
cc_101 VPB N_VPWR_c_442_n 0.00323736f $X=-0.19 $Y=1.305 $X2=5.155 $Y2=1.985
cc_102 VPB N_VPWR_c_443_n 0.017949f $X=-0.19 $Y=1.305 $X2=6.415 $Y2=1.985
cc_103 VPB N_VPWR_c_444_n 0.00323736f $X=-0.19 $Y=1.305 $X2=6.835 $Y2=1.985
cc_104 VPB N_VPWR_c_445_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_105 VPB N_VPWR_c_419_n 0.0517919f $X=-0.19 $Y=1.305 $X2=4.285 $Y2=1.105
cc_106 N_A_M1000_g N_VPWR_c_421_n 0.0031902f $X=0.535 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_c_122_n N_VPWR_c_421_n 0.0165339f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_c_123_n N_VPWR_c_421_n 0.00488545f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VPWR_c_422_n 0.00541359f $X=0.535 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_VPWR_c_422_n 0.00541359f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_VPWR_c_423_n 0.00146448f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1002_g N_VPWR_c_423_n 0.00146448f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_M1003_g N_VPWR_c_424_n 0.00146448f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_M1004_g N_VPWR_c_424_n 0.00146448f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_M1006_g N_VPWR_c_425_n 0.00146448f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_M1009_g N_VPWR_c_425_n 0.00146448f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_M1010_g N_VPWR_c_426_n 0.00146448f $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_M1014_g N_VPWR_c_426_n 0.00146448f $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_119 N_A_M1015_g N_VPWR_c_427_n 0.00146448f $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A_M1017_g N_VPWR_c_427_n 0.00146448f $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A_M1017_g N_VPWR_c_428_n 0.00541359f $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_M1020_g N_VPWR_c_428_n 0.00541359f $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A_M1020_g N_VPWR_c_429_n 0.00146448f $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_M1021_g N_VPWR_c_429_n 0.00146448f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_125 N_A_M1025_g N_VPWR_c_430_n 0.00146448f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_126 N_A_M1030_g N_VPWR_c_430_n 0.00146448f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A_M1031_g N_VPWR_c_432_n 0.0031902f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_M1002_g N_VPWR_c_433_n 0.00541359f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_M1003_g N_VPWR_c_433_n 0.00541359f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_130 N_A_M1004_g N_VPWR_c_435_n 0.00541359f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_M1006_g N_VPWR_c_435_n 0.00541359f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_M1009_g N_VPWR_c_437_n 0.00541359f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_133 N_A_M1010_g N_VPWR_c_437_n 0.00541359f $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A_M1014_g N_VPWR_c_439_n 0.00541359f $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_M1015_g N_VPWR_c_439_n 0.00541359f $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A_M1021_g N_VPWR_c_441_n 0.00541359f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A_M1025_g N_VPWR_c_441_n 0.00541359f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_138 N_A_M1030_g N_VPWR_c_443_n 0.00541359f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_139 N_A_M1031_g N_VPWR_c_443_n 0.00541359f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VPWR_c_419_n 0.0105125f $X=0.535 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VPWR_c_419_n 0.00950154f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VPWR_c_419_n 0.00950154f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_M1003_g N_VPWR_c_419_n 0.00950154f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_VPWR_c_419_n 0.00950154f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_M1006_g N_VPWR_c_419_n 0.00950154f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_M1009_g N_VPWR_c_419_n 0.00950154f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A_M1010_g N_VPWR_c_419_n 0.00950154f $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1014_g N_VPWR_c_419_n 0.00950154f $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_M1015_g N_VPWR_c_419_n 0.00950154f $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_M1017_g N_VPWR_c_419_n 0.00950154f $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_M1020_g N_VPWR_c_419_n 0.00950154f $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A_M1021_g N_VPWR_c_419_n 0.00950154f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_153 N_A_M1025_g N_VPWR_c_419_n 0.00950154f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_M1030_g N_VPWR_c_419_n 0.00950154f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1031_g N_VPWR_c_419_n 0.0105045f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_c_106_n N_Y_c_549_n 0.00528656f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_107_n N_Y_c_549_n 0.00620543f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_108_n N_Y_c_549_n 5.19281e-19 $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_M1000_g N_Y_c_552_n 0.00230941f $X=0.535 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1001_g N_Y_c_552_n 8.97266e-19 $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_c_122_n N_Y_c_552_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_c_123_n N_Y_c_552_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_M1000_g N_Y_c_556_n 0.00902485f $X=0.535 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1001_g N_Y_c_556_n 0.00975139f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_M1002_g N_Y_c_556_n 6.1949e-19 $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_c_107_n N_Y_c_535_n 0.00890471f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_108_n N_Y_c_535_n 0.00890471f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_122_n N_Y_c_535_n 0.0367667f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_c_123_n N_Y_c_535_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_106_n N_Y_c_536_n 0.00346724f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_c_107_n N_Y_c_536_n 0.00116017f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_122_n N_Y_c_536_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_123_n N_Y_c_536_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_M1001_g N_Y_c_567_n 0.0107675f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_M1002_g N_Y_c_567_n 0.0107675f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_176 N_A_c_122_n N_Y_c_567_n 0.0305424f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_c_123_n N_Y_c_567_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_107_n N_Y_c_571_n 5.19281e-19 $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_108_n N_Y_c_571_n 0.00620543f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_109_n N_Y_c_571_n 0.00620543f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_110_n N_Y_c_571_n 5.19281e-19 $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_M1001_g N_Y_c_575_n 6.1949e-19 $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A_M1002_g N_Y_c_575_n 0.00975139f $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_M1003_g N_Y_c_575_n 0.00975139f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A_M1004_g N_Y_c_575_n 6.1949e-19 $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_c_109_n N_Y_c_537_n 0.00890471f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_110_n N_Y_c_537_n 0.00890471f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_122_n N_Y_c_537_n 0.0367667f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_c_123_n N_Y_c_537_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_M1003_g N_Y_c_583_n 0.0107675f $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_M1004_g N_Y_c_583_n 0.0107675f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A_c_122_n N_Y_c_583_n 0.0305424f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_123_n N_Y_c_583_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_c_109_n N_Y_c_587_n 5.19281e-19 $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_110_n N_Y_c_587_n 0.00620543f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_111_n N_Y_c_587_n 0.00620543f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_112_n N_Y_c_587_n 5.19281e-19 $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_M1003_g N_Y_c_591_n 6.1949e-19 $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A_M1004_g N_Y_c_591_n 0.00975139f $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A_M1006_g N_Y_c_591_n 0.00975139f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_Y_c_591_n 6.1949e-19 $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_c_111_n N_Y_c_538_n 0.00890471f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_c_112_n N_Y_c_538_n 0.00890471f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_122_n N_Y_c_538_n 0.0367667f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_c_123_n N_Y_c_538_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_M1006_g N_Y_c_599_n 0.0107675f $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A_M1009_g N_Y_c_599_n 0.0107675f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_c_122_n N_Y_c_599_n 0.0305424f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_c_123_n N_Y_c_599_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_c_111_n N_Y_c_603_n 5.19281e-19 $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_c_112_n N_Y_c_603_n 0.00620543f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_c_113_n N_Y_c_603_n 0.00620543f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_114_n N_Y_c_603_n 5.19281e-19 $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_M1006_g N_Y_c_607_n 6.1949e-19 $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_M1009_g N_Y_c_607_n 0.00975139f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_M1010_g N_Y_c_607_n 0.00975139f $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_M1014_g N_Y_c_607_n 6.1949e-19 $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_c_113_n N_Y_c_539_n 0.00890471f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_114_n N_Y_c_539_n 0.00890471f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_c_122_n N_Y_c_539_n 0.0367667f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_c_123_n N_Y_c_539_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_M1010_g N_Y_c_615_n 0.0107675f $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_M1014_g N_Y_c_615_n 0.0107675f $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_c_122_n N_Y_c_615_n 0.0305424f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_c_123_n N_Y_c_615_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_c_113_n N_Y_c_619_n 5.19281e-19 $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_114_n N_Y_c_619_n 0.00620543f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_115_n N_Y_c_619_n 0.00620543f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_c_116_n N_Y_c_619_n 5.19281e-19 $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_M1010_g N_Y_c_623_n 6.1949e-19 $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A_M1014_g N_Y_c_623_n 0.00975139f $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_M1015_g N_Y_c_623_n 0.00975139f $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_233 N_A_M1017_g N_Y_c_623_n 6.1949e-19 $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_c_115_n N_Y_c_540_n 0.00890471f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_116_n N_Y_c_540_n 0.00890471f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_122_n N_Y_c_540_n 0.0367667f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_c_123_n N_Y_c_540_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_M1015_g N_Y_c_631_n 0.0107675f $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_M1017_g N_Y_c_631_n 0.0107675f $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_c_122_n N_Y_c_631_n 0.0305424f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_c_123_n N_Y_c_631_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_c_115_n N_Y_c_635_n 5.19281e-19 $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_116_n N_Y_c_635_n 0.00620543f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_117_n N_Y_c_635_n 0.00620543f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_118_n N_Y_c_635_n 5.19281e-19 $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_M1015_g N_Y_c_639_n 6.1949e-19 $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_M1017_g N_Y_c_639_n 0.00975139f $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_M1020_g N_Y_c_639_n 0.00975139f $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_249 N_A_M1021_g N_Y_c_639_n 6.1949e-19 $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_c_117_n N_Y_c_541_n 0.00890471f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_118_n N_Y_c_541_n 0.0100977f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_122_n N_Y_c_541_n 0.0301313f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_c_123_n N_Y_c_541_n 0.00222429f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_M1020_g N_Y_c_647_n 0.0107675f $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_M1021_g N_Y_c_647_n 0.0119284f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_c_122_n N_Y_c_647_n 0.0242567f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_c_123_n N_Y_c_647_n 0.00202853f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_c_117_n N_Y_c_651_n 5.19281e-19 $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_c_118_n N_Y_c_651_n 0.00620543f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_119_n N_Y_c_651_n 0.00620543f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_c_120_n N_Y_c_651_n 5.19281e-19 $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_M1020_g N_Y_c_655_n 6.1949e-19 $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_M1021_g N_Y_c_655_n 0.00975139f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A_M1025_g N_Y_c_655_n 0.00975139f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A_M1030_g N_Y_c_655_n 6.1949e-19 $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_c_119_n N_Y_c_542_n 0.010415f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_120_n N_Y_c_542_n 0.010415f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_c_123_n N_Y_c_542_n 0.00267852f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_M1025_g N_Y_c_662_n 0.0122371f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_M1030_g N_Y_c_662_n 0.0122371f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_c_123_n N_Y_c_662_n 0.0024013f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_c_119_n N_Y_c_665_n 5.19281e-19 $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_c_120_n N_Y_c_665_n 0.00620543f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_c_121_n N_Y_c_665_n 0.00528656f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_M1025_g N_Y_c_668_n 6.1949e-19 $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_M1030_g N_Y_c_668_n 0.00975139f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_M1031_g N_Y_c_668_n 0.0145598f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_c_108_n N_Y_c_543_n 0.00116017f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_109_n N_Y_c_543_n 0.00116017f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A_c_122_n N_Y_c_543_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_281 N_A_c_123_n N_Y_c_543_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_M1002_g N_Y_c_675_n 8.97266e-19 $X=1.375 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_M1003_g N_Y_c_675_n 8.97266e-19 $X=1.795 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_c_122_n N_Y_c_675_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_c_123_n N_Y_c_675_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_286 N_A_c_110_n N_Y_c_544_n 0.00116017f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_c_111_n N_Y_c_544_n 0.00116017f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_c_122_n N_Y_c_544_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_c_123_n N_Y_c_544_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_M1004_g N_Y_c_683_n 8.97266e-19 $X=2.215 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_M1006_g N_Y_c_683_n 8.97266e-19 $X=2.635 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A_c_122_n N_Y_c_683_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A_c_123_n N_Y_c_683_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_c_112_n N_Y_c_545_n 0.00116017f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_c_113_n N_Y_c_545_n 0.00116017f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_c_122_n N_Y_c_545_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_c_123_n N_Y_c_545_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_M1009_g N_Y_c_691_n 8.97266e-19 $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_M1010_g N_Y_c_691_n 8.97266e-19 $X=3.475 $Y=1.985 $X2=0 $Y2=0
cc_300 N_A_c_122_n N_Y_c_691_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_c_123_n N_Y_c_691_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_c_114_n N_Y_c_546_n 0.00116017f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A_c_115_n N_Y_c_546_n 0.00116017f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_c_122_n N_Y_c_546_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_c_123_n N_Y_c_546_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_M1014_g N_Y_c_699_n 8.97266e-19 $X=3.895 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_M1015_g N_Y_c_699_n 8.97266e-19 $X=4.315 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_c_122_n N_Y_c_699_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A_c_123_n N_Y_c_699_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_c_116_n N_Y_c_547_n 0.00116017f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A_c_117_n N_Y_c_547_n 0.00116017f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_c_122_n N_Y_c_547_n 0.0268677f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_c_123_n N_Y_c_547_n 0.00230339f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_M1017_g N_Y_c_707_n 8.97266e-19 $X=4.735 $Y=1.985 $X2=0 $Y2=0
cc_315 N_A_M1020_g N_Y_c_707_n 8.97266e-19 $X=5.155 $Y=1.985 $X2=0 $Y2=0
cc_316 N_A_c_122_n N_Y_c_707_n 0.020356f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_c_123_n N_Y_c_707_n 0.00211153f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_c_118_n N_Y_c_548_n 0.00150603f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_119_n N_Y_c_548_n 0.00150603f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_123_n N_Y_c_548_n 0.00290662f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_M1021_g N_Y_c_714_n 0.00122966f $X=5.575 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_M1025_g N_Y_c_714_n 0.00122966f $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_c_123_n N_Y_c_714_n 0.00263133f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_M1030_g N_Y_c_717_n 4.64231e-19 $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_325 N_A_M1031_g N_Y_c_717_n 0.00807109f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_c_119_n Y 4.37161e-19 $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_M1025_g Y 8.32629e-19 $X=5.995 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_c_120_n Y 0.0033952f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_M1030_g Y 0.0049513f $X=6.415 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_c_121_n Y 0.00792396f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_M1031_g Y 0.0091927f $X=6.835 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_c_123_n Y 0.0439472f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_c_106_n N_VGND_c_824_n 0.00320188f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_c_122_n N_VGND_c_824_n 0.0166874f $X=5.36 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_c_123_n N_VGND_c_824_n 0.00577382f $X=6.835 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_c_106_n N_VGND_c_825_n 0.00541359f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A_c_107_n N_VGND_c_825_n 0.00422241f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_c_107_n N_VGND_c_826_n 0.00146448f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_c_108_n N_VGND_c_826_n 0.00146448f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_c_109_n N_VGND_c_827_n 0.00146448f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A_c_110_n N_VGND_c_827_n 0.00146448f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A_c_111_n N_VGND_c_828_n 0.00146448f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A_c_112_n N_VGND_c_828_n 0.00146448f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A_c_113_n N_VGND_c_829_n 0.00146448f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A_c_114_n N_VGND_c_829_n 0.00146448f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A_c_115_n N_VGND_c_830_n 0.00146448f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A_c_116_n N_VGND_c_830_n 0.00146448f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A_c_116_n N_VGND_c_831_n 0.00422241f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A_c_117_n N_VGND_c_831_n 0.00422241f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A_c_117_n N_VGND_c_832_n 0.00146448f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A_c_118_n N_VGND_c_832_n 0.00146448f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A_c_119_n N_VGND_c_833_n 0.00146448f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A_c_120_n N_VGND_c_833_n 0.00146448f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_354 N_A_c_121_n N_VGND_c_835_n 0.0031902f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A_c_108_n N_VGND_c_836_n 0.00422241f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A_c_109_n N_VGND_c_836_n 0.00422241f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A_c_110_n N_VGND_c_838_n 0.00422241f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A_c_111_n N_VGND_c_838_n 0.00422241f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A_c_112_n N_VGND_c_840_n 0.00422241f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A_c_113_n N_VGND_c_840_n 0.00422241f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A_c_114_n N_VGND_c_842_n 0.00422241f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A_c_115_n N_VGND_c_842_n 0.00422241f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A_c_118_n N_VGND_c_844_n 0.00422241f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_c_119_n N_VGND_c_844_n 0.00422241f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A_c_120_n N_VGND_c_846_n 0.00422241f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A_c_121_n N_VGND_c_846_n 0.00541359f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A_c_106_n N_VGND_c_849_n 0.0105125f $X=0.535 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A_c_107_n N_VGND_c_849_n 0.00569656f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A_c_108_n N_VGND_c_849_n 0.00569656f $X=1.375 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A_c_109_n N_VGND_c_849_n 0.00569656f $X=1.795 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_c_110_n N_VGND_c_849_n 0.00569656f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A_c_111_n N_VGND_c_849_n 0.00569656f $X=2.635 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A_c_112_n N_VGND_c_849_n 0.00569656f $X=3.055 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A_c_113_n N_VGND_c_849_n 0.00569656f $X=3.475 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A_c_114_n N_VGND_c_849_n 0.00569656f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A_c_115_n N_VGND_c_849_n 0.00569656f $X=4.315 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A_c_116_n N_VGND_c_849_n 0.00569656f $X=4.735 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A_c_117_n N_VGND_c_849_n 0.00569656f $X=5.155 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A_c_118_n N_VGND_c_849_n 0.00569656f $X=5.575 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_c_119_n N_VGND_c_849_n 0.00569656f $X=5.995 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_c_120_n N_VGND_c_849_n 0.00569656f $X=6.415 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A_c_121_n N_VGND_c_849_n 0.0105045f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_383 N_VPWR_c_419_n N_Y_M1000_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_419_n N_Y_M1002_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_419_n N_Y_M1004_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_419_n N_Y_M1009_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_419_n N_Y_M1014_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_419_n N_Y_M1017_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_c_419_n N_Y_M1021_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_419_n N_Y_M1030_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_391 N_VPWR_c_422_n N_Y_c_556_n 0.0189039f $X=1.08 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_419_n N_Y_c_556_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_M1001_d N_Y_c_567_n 0.00314828f $X=1.03 $Y=1.485 $X2=0 $Y2=0
cc_394 N_VPWR_c_423_n N_Y_c_567_n 0.0126919f $X=1.165 $Y=2 $X2=0 $Y2=0
cc_395 N_VPWR_c_433_n N_Y_c_575_n 0.0189039f $X=1.92 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_419_n N_Y_c_575_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_M1003_d N_Y_c_583_n 0.00314828f $X=1.87 $Y=1.485 $X2=0 $Y2=0
cc_398 N_VPWR_c_424_n N_Y_c_583_n 0.0126919f $X=2.005 $Y=2 $X2=0 $Y2=0
cc_399 N_VPWR_c_435_n N_Y_c_591_n 0.0189039f $X=2.76 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_419_n N_Y_c_591_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_M1006_d N_Y_c_599_n 0.00314828f $X=2.71 $Y=1.485 $X2=0 $Y2=0
cc_402 N_VPWR_c_425_n N_Y_c_599_n 0.0126919f $X=2.845 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_437_n N_Y_c_607_n 0.0189039f $X=3.6 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_419_n N_Y_c_607_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1010_d N_Y_c_615_n 0.00314828f $X=3.55 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_c_426_n N_Y_c_615_n 0.0126919f $X=3.685 $Y=2 $X2=0 $Y2=0
cc_407 N_VPWR_c_439_n N_Y_c_623_n 0.0189039f $X=4.44 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_419_n N_Y_c_623_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_M1015_d N_Y_c_631_n 0.00314828f $X=4.39 $Y=1.485 $X2=0 $Y2=0
cc_410 N_VPWR_c_427_n N_Y_c_631_n 0.0126919f $X=4.525 $Y=2 $X2=0 $Y2=0
cc_411 N_VPWR_c_428_n N_Y_c_639_n 0.0189039f $X=5.28 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_419_n N_Y_c_639_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_M1020_d N_Y_c_647_n 0.00314828f $X=5.23 $Y=1.485 $X2=0 $Y2=0
cc_414 N_VPWR_c_429_n N_Y_c_647_n 0.0126919f $X=5.365 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_441_n N_Y_c_655_n 0.0189039f $X=6.12 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_419_n N_Y_c_655_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_M1025_d N_Y_c_662_n 0.00406737f $X=6.07 $Y=1.485 $X2=0 $Y2=0
cc_418 N_VPWR_c_430_n N_Y_c_662_n 0.0126919f $X=6.205 $Y=2 $X2=0 $Y2=0
cc_419 N_VPWR_c_443_n N_Y_c_668_n 0.0189039f $X=6.96 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_419_n N_Y_c_668_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_421 N_Y_c_535_n N_VGND_M1007_s 0.00162148f $X=1.42 $Y=0.81 $X2=0 $Y2=0
cc_422 N_Y_c_537_n N_VGND_M1011_s 0.00162148f $X=2.26 $Y=0.81 $X2=0 $Y2=0
cc_423 N_Y_c_538_n N_VGND_M1013_s 0.00162148f $X=3.1 $Y=0.81 $X2=0 $Y2=0
cc_424 N_Y_c_539_n N_VGND_M1018_s 0.00162148f $X=3.94 $Y=0.81 $X2=0 $Y2=0
cc_425 N_Y_c_540_n N_VGND_M1022_s 0.00162148f $X=4.78 $Y=0.81 $X2=0 $Y2=0
cc_426 N_Y_c_541_n N_VGND_M1024_s 0.00162148f $X=5.62 $Y=0.81 $X2=0 $Y2=0
cc_427 N_Y_c_542_n N_VGND_M1027_s 0.00162148f $X=6.46 $Y=0.81 $X2=0 $Y2=0
cc_428 N_Y_c_549_n N_VGND_c_825_n 0.0188551f $X=0.745 $Y=0.38 $X2=0 $Y2=0
cc_429 N_Y_c_535_n N_VGND_c_825_n 0.00203746f $X=1.42 $Y=0.81 $X2=0 $Y2=0
cc_430 N_Y_c_535_n N_VGND_c_826_n 0.0122675f $X=1.42 $Y=0.81 $X2=0 $Y2=0
cc_431 N_Y_c_537_n N_VGND_c_827_n 0.0122675f $X=2.26 $Y=0.81 $X2=0 $Y2=0
cc_432 N_Y_c_538_n N_VGND_c_828_n 0.0122675f $X=3.1 $Y=0.81 $X2=0 $Y2=0
cc_433 N_Y_c_539_n N_VGND_c_829_n 0.0122675f $X=3.94 $Y=0.81 $X2=0 $Y2=0
cc_434 N_Y_c_540_n N_VGND_c_830_n 0.0122675f $X=4.78 $Y=0.81 $X2=0 $Y2=0
cc_435 N_Y_c_540_n N_VGND_c_831_n 0.00203746f $X=4.78 $Y=0.81 $X2=0 $Y2=0
cc_436 N_Y_c_635_n N_VGND_c_831_n 0.0188551f $X=4.945 $Y=0.38 $X2=0 $Y2=0
cc_437 N_Y_c_541_n N_VGND_c_831_n 0.00203746f $X=5.62 $Y=0.81 $X2=0 $Y2=0
cc_438 N_Y_c_541_n N_VGND_c_832_n 0.0122675f $X=5.62 $Y=0.81 $X2=0 $Y2=0
cc_439 N_Y_c_542_n N_VGND_c_833_n 0.0122675f $X=6.46 $Y=0.81 $X2=0 $Y2=0
cc_440 N_Y_c_535_n N_VGND_c_836_n 0.00203746f $X=1.42 $Y=0.81 $X2=0 $Y2=0
cc_441 N_Y_c_571_n N_VGND_c_836_n 0.0188551f $X=1.585 $Y=0.38 $X2=0 $Y2=0
cc_442 N_Y_c_537_n N_VGND_c_836_n 0.00203746f $X=2.26 $Y=0.81 $X2=0 $Y2=0
cc_443 N_Y_c_537_n N_VGND_c_838_n 0.00203746f $X=2.26 $Y=0.81 $X2=0 $Y2=0
cc_444 N_Y_c_587_n N_VGND_c_838_n 0.0188551f $X=2.425 $Y=0.38 $X2=0 $Y2=0
cc_445 N_Y_c_538_n N_VGND_c_838_n 0.00203746f $X=3.1 $Y=0.81 $X2=0 $Y2=0
cc_446 N_Y_c_538_n N_VGND_c_840_n 0.00203746f $X=3.1 $Y=0.81 $X2=0 $Y2=0
cc_447 N_Y_c_603_n N_VGND_c_840_n 0.0188551f $X=3.265 $Y=0.38 $X2=0 $Y2=0
cc_448 N_Y_c_539_n N_VGND_c_840_n 0.00203746f $X=3.94 $Y=0.81 $X2=0 $Y2=0
cc_449 N_Y_c_539_n N_VGND_c_842_n 0.00203746f $X=3.94 $Y=0.81 $X2=0 $Y2=0
cc_450 N_Y_c_619_n N_VGND_c_842_n 0.0188551f $X=4.105 $Y=0.38 $X2=0 $Y2=0
cc_451 N_Y_c_540_n N_VGND_c_842_n 0.00203746f $X=4.78 $Y=0.81 $X2=0 $Y2=0
cc_452 N_Y_c_541_n N_VGND_c_844_n 0.00203746f $X=5.62 $Y=0.81 $X2=0 $Y2=0
cc_453 N_Y_c_651_n N_VGND_c_844_n 0.0188551f $X=5.785 $Y=0.38 $X2=0 $Y2=0
cc_454 N_Y_c_542_n N_VGND_c_844_n 0.00203746f $X=6.46 $Y=0.81 $X2=0 $Y2=0
cc_455 N_Y_c_542_n N_VGND_c_846_n 0.00203746f $X=6.46 $Y=0.81 $X2=0 $Y2=0
cc_456 N_Y_c_665_n N_VGND_c_846_n 0.0189039f $X=6.625 $Y=0.38 $X2=0 $Y2=0
cc_457 N_Y_M1005_d N_VGND_c_849_n 0.00215201f $X=0.61 $Y=0.235 $X2=0 $Y2=0
cc_458 N_Y_M1008_d N_VGND_c_849_n 0.00215201f $X=1.45 $Y=0.235 $X2=0 $Y2=0
cc_459 N_Y_M1012_d N_VGND_c_849_n 0.00215201f $X=2.29 $Y=0.235 $X2=0 $Y2=0
cc_460 N_Y_M1016_d N_VGND_c_849_n 0.00215201f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_461 N_Y_M1019_d N_VGND_c_849_n 0.00215201f $X=3.97 $Y=0.235 $X2=0 $Y2=0
cc_462 N_Y_M1023_d N_VGND_c_849_n 0.00215201f $X=4.81 $Y=0.235 $X2=0 $Y2=0
cc_463 N_Y_M1026_d N_VGND_c_849_n 0.00215201f $X=5.65 $Y=0.235 $X2=0 $Y2=0
cc_464 N_Y_M1028_d N_VGND_c_849_n 0.00215201f $X=6.49 $Y=0.235 $X2=0 $Y2=0
cc_465 N_Y_c_549_n N_VGND_c_849_n 0.0122069f $X=0.745 $Y=0.38 $X2=0 $Y2=0
cc_466 N_Y_c_535_n N_VGND_c_849_n 0.00845923f $X=1.42 $Y=0.81 $X2=0 $Y2=0
cc_467 N_Y_c_571_n N_VGND_c_849_n 0.0122069f $X=1.585 $Y=0.38 $X2=0 $Y2=0
cc_468 N_Y_c_537_n N_VGND_c_849_n 0.00845923f $X=2.26 $Y=0.81 $X2=0 $Y2=0
cc_469 N_Y_c_587_n N_VGND_c_849_n 0.0122069f $X=2.425 $Y=0.38 $X2=0 $Y2=0
cc_470 N_Y_c_538_n N_VGND_c_849_n 0.00845923f $X=3.1 $Y=0.81 $X2=0 $Y2=0
cc_471 N_Y_c_603_n N_VGND_c_849_n 0.0122069f $X=3.265 $Y=0.38 $X2=0 $Y2=0
cc_472 N_Y_c_539_n N_VGND_c_849_n 0.00845923f $X=3.94 $Y=0.81 $X2=0 $Y2=0
cc_473 N_Y_c_619_n N_VGND_c_849_n 0.0122069f $X=4.105 $Y=0.38 $X2=0 $Y2=0
cc_474 N_Y_c_540_n N_VGND_c_849_n 0.00845923f $X=4.78 $Y=0.81 $X2=0 $Y2=0
cc_475 N_Y_c_635_n N_VGND_c_849_n 0.0122069f $X=4.945 $Y=0.38 $X2=0 $Y2=0
cc_476 N_Y_c_541_n N_VGND_c_849_n 0.00845923f $X=5.62 $Y=0.81 $X2=0 $Y2=0
cc_477 N_Y_c_651_n N_VGND_c_849_n 0.0122069f $X=5.785 $Y=0.38 $X2=0 $Y2=0
cc_478 N_Y_c_542_n N_VGND_c_849_n 0.00845923f $X=6.46 $Y=0.81 $X2=0 $Y2=0
cc_479 N_Y_c_665_n N_VGND_c_849_n 0.0122217f $X=6.625 $Y=0.38 $X2=0 $Y2=0

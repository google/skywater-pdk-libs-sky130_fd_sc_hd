* File: sky130_fd_sc_hd__a2111o_1.pex.spice
* Created: Tue Sep  1 18:50:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2111O_1%A_85_193# 1 2 3 12 14 16 20 22 23 24 25 30
+ 32 36 39 40 42
r82 41 42 5.08707 $w=3.79e-07 $l=4e-08 $layer=POLY_cond $X=0.5 $Y=1.15 $X2=0.54
+ $Y2=1.15
r83 34 36 8.38581 $w=2.03e-07 $l=1.55e-07 $layer=LI1_cond $X=2.702 $Y=0.655
+ $X2=2.702 $Y2=0.5
r84 33 40 8.52281 $w=1.72e-07 $l=1.66493e-07 $layer=LI1_cond $X=1.915 $Y=0.74
+ $X2=1.75 $Y2=0.737
r85 32 34 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=2.6 $Y=0.74
+ $X2=2.702 $Y2=0.655
r86 32 33 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.6 $Y=0.74
+ $X2=1.915 $Y2=0.74
r87 28 40 0.850971 $w=3.3e-07 $l=8.7e-08 $layer=LI1_cond $X=1.75 $Y=0.65
+ $X2=1.75 $Y2=0.737
r88 28 30 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.75 $Y=0.65
+ $X2=1.75 $Y2=0.39
r89 24 39 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=1.135 $Y=1.555
+ $X2=1.24 $Y2=1.555
r90 24 25 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=1.135 $Y=1.555
+ $X2=0.915 $Y2=1.555
r91 22 40 8.52281 $w=1.72e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0.737
+ $X2=1.75 $Y2=0.737
r92 22 23 42.4623 $w=1.73e-07 $l=6.7e-07 $layer=LI1_cond $X=1.585 $Y=0.737
+ $X2=0.915 $Y2=0.737
r93 21 42 33.7018 $w=3.79e-07 $l=2.65e-07 $layer=POLY_cond $X=0.805 $Y=1.15
+ $X2=0.54 $Y2=1.15
r94 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.16 $X2=0.805 $Y2=1.16
r95 18 25 6.90553 $w=1.8e-07 $l=1.48324e-07 $layer=LI1_cond $X=0.805 $Y=1.465
+ $X2=0.915 $Y2=1.555
r96 18 20 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=0.805 $Y=1.465
+ $X2=0.805 $Y2=1.16
r97 17 23 6.93219 $w=1.75e-07 $l=1.4758e-07 $layer=LI1_cond $X=0.805 $Y=0.825
+ $X2=0.915 $Y2=0.737
r98 17 20 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=0.805 $Y=0.825
+ $X2=0.805 $Y2=1.16
r99 14 42 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.54 $Y=0.96
+ $X2=0.54 $Y2=1.15
r100 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.54 $Y=0.96 $X2=0.54
+ $Y2=0.56
r101 10 41 24.5487 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.5 $Y=1.34 $X2=0.5
+ $Y2=1.15
r102 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.5 $Y=1.34
+ $X2=0.5 $Y2=1.985
r103 3 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.485 $X2=1.26 $Y2=1.63
r104 2 36 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=2.58
+ $Y=0.235 $X2=2.72 $Y2=0.5
r105 1 30 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=1.61
+ $Y=0.235 $X2=1.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%D1 3 6 8 9 10 11 17 19 32
r44 21 32 1.68648 $w=2.05e-07 $l=1.2e-07 $layer=LI1_cond $X=1.617 $Y=1.29
+ $X2=1.617 $Y2=1.17
r45 17 20 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.495 $Y2=1.325
r46 17 19 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.495 $Y2=0.995
r47 10 11 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.617 $Y=1.87
+ $X2=1.617 $Y2=2.21
r48 9 10 18.3947 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.617 $Y=1.53
+ $X2=1.617 $Y2=1.87
r49 9 21 12.9845 $w=2.03e-07 $l=2.4e-07 $layer=LI1_cond $X=1.617 $Y=1.53
+ $X2=1.617 $Y2=1.29
r50 8 32 4.17761 $w=2.38e-07 $l=8.7e-08 $layer=LI1_cond $X=1.53 $Y=1.17
+ $X2=1.617 $Y2=1.17
r51 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.53
+ $Y=1.16 $X2=1.53 $Y2=1.16
r52 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.595 $Y=1.985
+ $X2=1.595 $Y2=1.325
r53 3 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.535 $Y=0.56
+ $X2=1.535 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%C1 3 6 7 8 9 10 16 18 19
r33 16 19 58.9771 $w=3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.07 $Y=1.16 $X2=2.07
+ $Y2=1.38
r34 16 18 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.16 $X2=2.07
+ $Y2=0.995
r35 9 10 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.055 $Y=1.87
+ $X2=2.055 $Y2=2.21
r36 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.055 $Y=1.53
+ $X2=2.055 $Y2=1.87
r37 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.055 $Y=1.16
+ $X2=2.055 $Y2=1.53
r38 7 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=1.16 $X2=2.055 $Y2=1.16
r39 6 19 194.407 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=1.995 $Y=1.985
+ $X2=1.995 $Y2=1.38
r40 3 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.995 $Y=0.56
+ $X2=1.995 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%B1 3 6 8 9 10 11 17 19
c37 17 0 1.21878e-19 $X=2.595 $Y=1.16
r38 17 20 47.0858 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.595 $Y2=1.33
r39 17 19 52.3316 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.595 $Y=1.16
+ $X2=2.595 $Y2=0.96
r40 10 11 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.54 $Y=1.87 $X2=2.54
+ $Y2=2.21
r41 9 10 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.54 $Y=1.53 $X2=2.54
+ $Y2=1.87
r42 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.54 $Y=1.16 $X2=2.54
+ $Y2=1.53
r43 8 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.595
+ $Y=1.16 $X2=2.595 $Y2=1.16
r44 6 20 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.505 $Y=1.985
+ $X2=2.505 $Y2=1.33
r45 3 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.505 $Y=0.56 $X2=2.505
+ $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%A1 1 3 5 7 8 9
c40 5 0 1.21878e-19 $X=3.225 $Y=0.965
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.145
+ $Y=1.16 $X2=3.145 $Y2=1.16
r42 9 14 17.0538 $w=4.65e-07 $l=6.5e-07 $layer=LI1_cond $X=3.222 $Y=0.51
+ $X2=3.222 $Y2=1.16
r43 8 14 0.787097 $w=4.65e-07 $l=3e-08 $layer=LI1_cond $X=3.222 $Y=1.19
+ $X2=3.222 $Y2=1.16
r44 5 13 42.9359 $w=3.39e-07 $l=2.31571e-07 $layer=POLY_cond $X=3.225 $Y=0.965
+ $X2=3.145 $Y2=1.16
r45 5 7 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.225 $Y=0.965
+ $X2=3.225 $Y2=0.56
r46 1 13 39.3813 $w=3.39e-07 $l=2.0199e-07 $layer=POLY_cond $X=3.215 $Y=1.33
+ $X2=3.145 $Y2=1.16
r47 1 3 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.215 $Y=1.33
+ $X2=3.215 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%A2 3 6 8 11 13
r24 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=1.16
+ $X2=3.725 $Y2=1.325
r25 11 13 51.398 $w=3.4e-07 $l=1.95e-07 $layer=POLY_cond $X=3.725 $Y=1.16
+ $X2=3.725 $Y2=0.965
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.16 $X2=3.71 $Y2=1.16
r27 8 12 8.69768 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=3.91 $Y=1.157 $X2=3.71
+ $Y2=1.157
r28 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.635 $Y=1.985
+ $X2=3.635 $Y2=1.325
r29 3 13 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.63 $Y=0.56 $X2=3.63
+ $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%X 1 2 7 8 9 10 11 12 22 39
r16 20 39 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.3 $Y=1.455 $X2=0.3
+ $Y2=1.53
r17 11 12 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.262 $Y=1.87
+ $X2=0.262 $Y2=2.21
r18 11 42 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=0.262 $Y=1.87
+ $X2=0.262 $Y2=1.62
r19 10 42 3.5937 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.3 $Y=1.535 $X2=0.3
+ $Y2=1.62
r20 10 39 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.3 $Y=1.535 $X2=0.3
+ $Y2=1.53
r21 10 20 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.3 $Y=1.45 $X2=0.3
+ $Y2=1.455
r22 9 10 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.3 $Y=1.19 $X2=0.3
+ $Y2=1.45
r23 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.3 $Y=0.85 $X2=0.3
+ $Y2=1.19
r24 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.3 $Y=0.51 $X2=0.3
+ $Y2=0.85
r25 7 22 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.3 $Y=0.51 $X2=0.3
+ $Y2=0.4
r26 2 10 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.61
r27 2 12 400 $w=1.7e-07 $l=8.79517e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.295
r28 1 22 91 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.3 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%VPWR 1 2 9 13 15 17 22 32 33 36 39
r51 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r54 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 30 39 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.54 $Y=2.72
+ $X2=3.432 $Y2=2.72
r56 30 32 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.54 $Y=2.72 $X2=3.91
+ $Y2=2.72
r57 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 26 29 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 25 28 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.73 $Y2=2.72
r64 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 22 39 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.432 $Y2=2.72
r66 22 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.73 $Y2=2.72
r68 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 11 39 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.432 $Y=2.635
+ $X2=3.432 $Y2=2.72
r72 11 13 33.7693 $w=2.13e-07 $l=6.3e-07 $layer=LI1_cond $X=3.432 $Y=2.635
+ $X2=3.432 $Y2=2.005
r73 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r74 7 9 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=1.98
r75 2 13 300 $w=1.7e-07 $l=5.83609e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=1.485 $X2=3.425 $Y2=2.005
r76 1 9 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=1.485 $X2=0.715 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%A_516_297# 1 2 9 11 12 15
r23 13 15 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=1.665
+ $X2=3.855 $Y2=1.89
r24 11 13 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.72 $Y=1.58
+ $X2=3.855 $Y2=1.665
r25 11 12 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.72 $Y=1.58
+ $X2=3.145 $Y2=1.58
r26 7 12 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.002 $Y=1.665
+ $X2=3.145 $Y2=1.58
r27 7 9 3.03274 $w=2.83e-07 $l=7.5e-08 $layer=LI1_cond $X=3.002 $Y=1.665
+ $X2=3.002 $Y2=1.74
r28 2 15 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=3.71
+ $Y=1.485 $X2=3.855 $Y2=1.89
r29 1 9 300 $w=1.7e-07 $l=5.37587e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.485 $X2=3.005 $Y2=1.74
.ends

.subckt PM_SKY130_FD_SC_HD__A2111O_1%VGND 1 2 3 14 16 18 21 22 23 29 37 45 48
r55 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r56 43 45 9.75637 $w=5.53e-07 $l=1.6e-07 $layer=LI1_cond $X=1.15 $Y=0.192
+ $X2=1.31 $Y2=0.192
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 41 43 0.107755 $w=5.53e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=0.192
+ $X2=1.15 $Y2=0.192
r59 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r60 37 41 9.80569 $w=5.53e-07 $l=4.55e-07 $layer=LI1_cond $X=0.69 $Y=0.192
+ $X2=1.145 $Y2=0.192
r61 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r62 35 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r63 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r64 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r65 31 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r66 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r67 29 47 3.8575 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.927
+ $Y2=0
r68 29 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.45
+ $Y2=0
r69 28 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r70 28 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r71 27 45 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.31
+ $Y2=0
r72 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 23 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r74 21 27 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.07
+ $Y2=0
r75 21 22 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.257
+ $Y2=0
r76 20 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.53
+ $Y2=0
r77 20 22 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.257
+ $Y2=0
r78 16 47 3.22065 $w=2.4e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.927 $Y2=0
r79 16 18 18.7272 $w=2.38e-07 $l=3.9e-07 $layer=LI1_cond $X=3.835 $Y=0.085
+ $X2=3.835 $Y2=0.475
r80 12 22 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.257 $Y=0.085
+ $X2=2.257 $Y2=0
r81 12 14 10.5223 $w=3.43e-07 $l=3.15e-07 $layer=LI1_cond $X=2.257 $Y=0.085
+ $X2=2.257 $Y2=0.4
r82 3 18 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.845 $Y2=0.475
r83 2 14 182 $w=1.7e-07 $l=2.49199e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.25 $Y2=0.4
r84 1 41 91 $w=1.7e-07 $l=5.89194e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=0.235 $X2=1.145 $Y2=0.36
.ends


* File: sky130_fd_sc_hd__buf_1.spice.pex
* Created: Thu Aug 27 14:09:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__BUF_1%A 1 3 5 8 9 10 11
c34 11 0 6.72902e-20 $X=0.23 $Y=1.19
c35 10 0 1.55858e-19 $X=0.455 $Y=1.62
r36 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r37 9 10 46.6452 $w=1.8e-07 $l=1.2e-07 $layer=POLY_cond $X=0.455 $Y=1.5
+ $X2=0.455 $Y2=1.62
r38 8 10 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.47 $Y=2.09 $X2=0.47
+ $Y2=1.62
r39 3 14 64.1867 $w=3.1e-07 $l=3.89615e-07 $layer=POLY_cond $X=0.47 $Y=0.83
+ $X2=0.34 $Y2=1.16
r40 3 5 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.47 $Y=0.83 $X2=0.47
+ $Y2=0.495
r41 1 14 38.5318 $w=3.1e-07 $l=2.09105e-07 $layer=POLY_cond $X=0.44 $Y=1.325
+ $X2=0.34 $Y2=1.16
r42 1 9 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.44 $Y=1.325 $X2=0.44
+ $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_1%A_27_47# 1 2 9 13 17 21 23 24 25 26 30 32 33
+ 34
c67 23 0 1.55858e-19 $X=0.67 $Y=0.72
c68 9 0 6.72902e-20 $X=0.91 $Y=0.495
r69 33 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.86 $Y=1.225
+ $X2=0.86 $Y2=1.39
r70 33 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.86 $Y=1.225
+ $X2=0.86 $Y2=1.06
r71 32 35 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.807 $Y=1.225
+ $X2=0.807 $Y2=1.39
r72 32 34 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.807 $Y=1.225
+ $X2=0.807 $Y2=1.06
r73 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.86
+ $Y=1.225 $X2=0.86 $Y2=1.225
r74 30 35 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.755 $Y=1.535
+ $X2=0.755 $Y2=1.39
r75 27 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.755 $Y=0.805
+ $X2=0.755 $Y2=1.06
r76 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.67 $Y=1.62
+ $X2=0.755 $Y2=1.535
r77 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.67 $Y=1.62
+ $X2=0.345 $Y2=1.62
r78 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.67 $Y=0.72
+ $X2=0.755 $Y2=0.805
r79 23 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.67 $Y=0.72
+ $X2=0.345 $Y2=0.72
r80 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r81 19 21 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.445
r82 15 26 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.255 $Y=1.705
+ $X2=0.345 $Y2=1.62
r83 15 17 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.255 $Y=1.705
+ $X2=0.255 $Y2=1.96
r84 13 38 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.91 $Y=2.09 $X2=0.91
+ $Y2=1.39
r85 9 37 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.91 $Y=0.495
+ $X2=0.91 $Y2=1.06
r86 2 17 300 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.695 $X2=0.26 $Y2=1.96
r87 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_1%VPWR 1 6 8 10 12 20 21 24
r22 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r23 21 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r24 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r26 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r27 12 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r28 10 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r29 8 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.525 $Y2=2.72
r30 8 10 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r31 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.72
r32 4 6 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=1.96
r33 1 6 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.695 $X2=0.69 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_1%X 1 2 9 10 12 13 14 15
r24 14 15 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.16 $Y=1.87
+ $X2=1.16 $Y2=2.21
r25 11 13 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=1.165 $Y=0.63
+ $X2=1.165 $Y2=0.51
r26 11 12 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.165 $Y=0.63
+ $X2=1.165 $Y2=0.76
r27 10 12 49.2929 $w=1.78e-07 $l=8e-07 $layer=LI1_cond $X=1.205 $Y=1.56
+ $X2=1.205 $Y2=0.76
r28 9 14 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.16 $Y=1.695
+ $X2=1.16 $Y2=1.87
r29 9 10 7.04571 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.16 $Y=1.695
+ $X2=1.16 $Y2=1.56
r30 2 14 300 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.695 $X2=1.12 $Y2=1.895
r31 1 13 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HD__BUF_1%VGND 1 6 8 10 12 17 21 22 25
r23 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r24 22 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r26 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r27 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.15
+ $Y2=0
r28 12 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r29 10 26 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r30 10 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r31 8 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.525
+ $Y2=0
r32 8 17 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.23
+ $Y2=0
r33 4 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r34 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r35 1 6 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o311ai_0.spice.SKY130_FD_SC_HD__O311AI_0.pxi
* Created: Thu Aug 27 14:39:17 2020
* 
x_PM_SKY130_FD_SC_HD__O311AI_0%A1 N_A1_M1005_g N_A1_M1008_g A1 A1 A1 N_A1_c_56_n
+ PM_SKY130_FD_SC_HD__O311AI_0%A1
x_PM_SKY130_FD_SC_HD__O311AI_0%A2 N_A2_M1000_g N_A2_M1001_g A2 A2 A2 A2
+ N_A2_c_82_n N_A2_c_83_n PM_SKY130_FD_SC_HD__O311AI_0%A2
x_PM_SKY130_FD_SC_HD__O311AI_0%A3 N_A3_M1004_g N_A3_M1009_g A3 N_A3_c_122_n
+ PM_SKY130_FD_SC_HD__O311AI_0%A3
x_PM_SKY130_FD_SC_HD__O311AI_0%B1 N_B1_M1002_g N_B1_M1007_g B1 N_B1_c_153_n
+ PM_SKY130_FD_SC_HD__O311AI_0%B1
x_PM_SKY130_FD_SC_HD__O311AI_0%C1 N_C1_M1006_g N_C1_M1003_g C1 C1 N_C1_c_189_n
+ PM_SKY130_FD_SC_HD__O311AI_0%C1
x_PM_SKY130_FD_SC_HD__O311AI_0%VPWR N_VPWR_M1008_s N_VPWR_M1002_d N_VPWR_c_214_n
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_218_n VPWR
+ N_VPWR_c_219_n N_VPWR_c_213_n PM_SKY130_FD_SC_HD__O311AI_0%VPWR
x_PM_SKY130_FD_SC_HD__O311AI_0%Y N_Y_M1006_d N_Y_M1009_d N_Y_M1003_d N_Y_c_256_n
+ Y Y Y Y Y Y Y Y Y PM_SKY130_FD_SC_HD__O311AI_0%Y
x_PM_SKY130_FD_SC_HD__O311AI_0%VGND N_VGND_M1005_s N_VGND_M1000_d N_VGND_c_301_n
+ N_VGND_c_302_n N_VGND_c_303_n N_VGND_c_304_n VGND N_VGND_c_305_n
+ N_VGND_c_306_n N_VGND_c_307_n PM_SKY130_FD_SC_HD__O311AI_0%VGND
x_PM_SKY130_FD_SC_HD__O311AI_0%A_138_47# N_A_138_47#_M1005_d N_A_138_47#_M1004_d
+ N_A_138_47#_c_362_n N_A_138_47#_c_344_n N_A_138_47#_c_345_n
+ N_A_138_47#_c_358_n PM_SKY130_FD_SC_HD__O311AI_0%A_138_47#
cc_1 VNB N_A1_M1005_g 0.035863f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_2 VNB A1 0.0304822f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_3 VNB N_A1_c_56_n 0.0335467f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.16
cc_4 VNB N_A2_M1000_g 0.0265096f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_5 VNB N_A2_c_82_n 0.0203352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A2_c_83_n 0.00331904f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_7 VNB N_A3_M1004_g 0.0311601f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_8 VNB A3 0.00405923f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_9 VNB N_A3_c_122_n 0.0215997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B1_M1007_g 0.0301025f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=2.165
cc_11 VNB B1 0.00346447f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_12 VNB N_B1_c_153_n 0.0265549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_C1_M1006_g 0.0314816f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=0.445
cc_14 VNB C1 0.0245479f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_15 VNB N_C1_c_189_n 0.04148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_213_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.0103443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.0194347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_301_n 0.0129726f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=2.165
cc_20 VNB N_VGND_c_302_n 0.0214654f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_21 VNB N_VGND_c_303_n 0.0117571f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_22 VNB N_VGND_c_304_n 3.95446e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_305_n 0.0476884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_306_n 0.181389f $X=-0.19 $Y=-0.24 $X2=0.432 $Y2=0.85
cc_25 VNB N_VGND_c_307_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0.432 $Y2=1.53
cc_26 VNB N_A_138_47#_c_344_n 0.0124928f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_27 VNB N_A_138_47#_c_345_n 0.00695153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_A1_M1008_g 0.0455848f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=2.165
cc_29 VPB A1 0.0213783f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_30 VPB N_A1_c_56_n 0.00938528f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.16
cc_31 VPB N_A2_M1001_g 0.0323189f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=2.165
cc_32 VPB N_A2_c_82_n 0.00567115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A2_c_83_n 0.00800646f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_34 VPB N_A3_M1009_g 0.0401533f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=2.165
cc_35 VPB A3 0.00132946f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_36 VPB N_A3_c_122_n 0.00409058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B1_M1002_g 0.0425324f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=0.445
cc_38 VPB N_B1_c_153_n 0.00555769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_C1_M1003_g 0.0451627f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=2.165
cc_40 VPB C1 0.0035685f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_41 VPB N_C1_c_189_n 0.01258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_214_n 0.0157691f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=2.165
cc_43 VPB N_VPWR_c_215_n 0.0428336f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_44 VPB N_VPWR_c_216_n 0.00850771f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_217_n 0.0346637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_218_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_219_n 0.0211349f $X=-0.19 $Y=1.305 $X2=0.432 $Y2=1.19
cc_48 VPB N_VPWR_c_213_n 0.0441037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_Y_c_256_n 0.0106449f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_50 VPB Y 0.0021058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB Y 0.00798423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB Y 0.0240089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB Y 0.0399824f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_54 N_A1_M1005_g N_A2_M1000_g 0.0231681f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_55 A1 N_A2_M1000_g 8.78978e-19 $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_56 N_A1_M1008_g N_A2_M1001_g 0.0603937f $X=0.615 $Y=2.165 $X2=0 $Y2=0
cc_57 A1 N_A2_M1001_g 0.00116229f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_58 A1 N_A2_c_82_n 0.00217873f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_59 N_A1_c_56_n N_A2_c_82_n 0.0202229f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A1_M1008_g N_A2_c_83_n 0.0049256f $X=0.615 $Y=2.165 $X2=0 $Y2=0
cc_61 A1 N_A2_c_83_n 0.054218f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_62 N_A1_c_56_n N_A2_c_83_n 3.16536e-19 $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A1_M1008_g N_VPWR_c_215_n 0.0248986f $X=0.615 $Y=2.165 $X2=0 $Y2=0
cc_64 A1 N_VPWR_c_215_n 0.0634689f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_65 N_A1_c_56_n N_VPWR_c_215_n 0.00111848f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A1_M1005_g N_VGND_c_302_n 0.00971354f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_67 A1 N_VGND_c_302_n 0.0404739f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_68 N_A1_c_56_n N_VGND_c_302_n 0.00115443f $X=0.615 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A1_M1005_g N_VGND_c_303_n 0.0046653f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A1_M1005_g N_VGND_c_304_n 5.43479e-19 $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A1_M1005_g N_VGND_c_306_n 0.00799591f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_72 A1 N_VGND_c_306_n 0.00194633f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_73 N_A1_M1005_g N_A_138_47#_c_345_n 0.00394031f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_74 A1 N_A_138_47#_c_345_n 0.00889989f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_75 N_A2_M1000_g N_A3_M1004_g 0.0273838f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A2_M1001_g N_A3_M1009_g 0.0559319f $X=1.035 $Y=2.165 $X2=0 $Y2=0
cc_77 N_A2_c_82_n A3 3.17145e-19 $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A2_c_83_n A3 0.0260652f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A2_c_82_n N_A3_c_122_n 0.0201765f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A2_c_83_n N_A3_c_122_n 0.012364f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_M1001_g N_VPWR_c_215_n 0.00549662f $X=1.035 $Y=2.165 $X2=0 $Y2=0
cc_82 N_A2_c_83_n N_VPWR_c_215_n 0.0321307f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A2_M1001_g N_VPWR_c_217_n 0.00357668f $X=1.035 $Y=2.165 $X2=0 $Y2=0
cc_84 N_A2_c_83_n N_VPWR_c_217_n 0.0190383f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A2_M1001_g N_VPWR_c_213_n 0.00532039f $X=1.035 $Y=2.165 $X2=0 $Y2=0
cc_86 N_A2_c_83_n N_VPWR_c_213_n 0.0111757f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A2_c_83_n A_222_369# 0.00610622f $X=1.035 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_88 N_A2_c_83_n N_Y_c_256_n 0.0141978f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A2_M1001_g Y 7.31762e-19 $X=1.035 $Y=2.165 $X2=0 $Y2=0
cc_90 N_A2_c_83_n Y 0.0644682f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A2_M1000_g N_VGND_c_302_n 5.83631e-19 $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A2_M1000_g N_VGND_c_303_n 0.00341689f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A2_M1000_g N_VGND_c_304_n 0.00681952f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A2_M1000_g N_VGND_c_306_n 0.00405445f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A2_M1000_g N_A_138_47#_c_344_n 0.0109948f $X=1.035 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A2_c_82_n N_A_138_47#_c_344_n 0.00200929f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A2_c_83_n N_A_138_47#_c_344_n 0.0244575f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A2_c_82_n N_A_138_47#_c_345_n 4.33113e-19 $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A3_M1009_g N_B1_M1002_g 0.0297906f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_100 N_A3_M1004_g N_B1_M1007_g 0.00999806f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A3_M1004_g B1 0.00415172f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_102 A3 B1 0.0221833f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A3_c_122_n B1 3.42843e-19 $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_104 A3 N_B1_c_153_n 0.00235967f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_105 N_A3_c_122_n N_B1_c_153_n 0.0113895f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A3_M1009_g N_VPWR_c_217_n 0.00435091f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_107 N_A3_M1009_g N_VPWR_c_213_n 0.00760094f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_108 N_A3_M1009_g N_Y_c_256_n 0.0068437f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_109 A3 N_Y_c_256_n 0.0296025f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_110 N_A3_c_122_n N_Y_c_256_n 0.00279548f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A3_M1009_g Y 0.0255298f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_112 N_A3_M1004_g N_VGND_c_304_n 0.00853411f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A3_M1004_g N_VGND_c_305_n 0.00341689f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A3_M1004_g N_VGND_c_306_n 0.00470573f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A3_M1004_g N_A_138_47#_c_344_n 0.0135051f $X=1.455 $Y=0.445 $X2=0 $Y2=0
cc_116 A3 N_A_138_47#_c_344_n 0.0254058f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A3_c_122_n N_A_138_47#_c_344_n 0.00273862f $X=1.515 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B1_M1007_g N_C1_M1006_g 0.0371457f $X=2.215 $Y=0.445 $X2=0 $Y2=0
cc_119 B1 N_C1_M1006_g 0.00107472f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_M1002_g N_C1_M1003_g 0.0201331f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_121 N_B1_c_153_n N_C1_c_189_n 0.0371457f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B1_M1002_g N_VPWR_c_216_n 0.00329424f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_VPWR_c_217_n 0.00585385f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_124 N_B1_M1002_g N_VPWR_c_213_n 0.0112137f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_125 N_B1_M1002_g N_Y_c_256_n 0.00280657f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_126 N_B1_M1002_g Y 0.00783906f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_127 N_B1_M1002_g Y 0.0032004f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_128 N_B1_M1007_g Y 0.00432365f $X=2.215 $Y=0.445 $X2=0 $Y2=0
cc_129 B1 Y 0.0394281f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_130 N_B1_M1002_g Y 0.0133675f $X=2.055 $Y=2.165 $X2=0 $Y2=0
cc_131 B1 Y 0.0165624f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B1_c_153_n Y 0.00554139f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B1_M1007_g N_VGND_c_305_n 0.004948f $X=2.215 $Y=0.445 $X2=0 $Y2=0
cc_134 B1 N_VGND_c_305_n 0.0125248f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_135 N_B1_M1007_g N_VGND_c_306_n 0.00913796f $X=2.215 $Y=0.445 $X2=0 $Y2=0
cc_136 B1 N_VGND_c_306_n 0.00798122f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_137 B1 N_A_138_47#_M1004_d 0.00518979f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_138 N_B1_M1007_g N_A_138_47#_c_344_n 6.18624e-19 $X=2.215 $Y=0.445 $X2=0
+ $Y2=0
cc_139 B1 N_A_138_47#_c_344_n 0.0116664f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_140 N_B1_M1007_g N_A_138_47#_c_358_n 0.0012399f $X=2.215 $Y=0.445 $X2=0 $Y2=0
cc_141 B1 N_A_138_47#_c_358_n 0.0229979f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_142 N_C1_M1003_g N_VPWR_c_216_n 0.00329424f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_143 N_C1_M1003_g N_VPWR_c_219_n 0.00585385f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_144 N_C1_M1003_g N_VPWR_c_213_n 0.0118001f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_145 N_C1_M1006_g Y 0.00706187f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_146 N_C1_M1006_g Y 0.0117356f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_147 N_C1_M1003_g Y 0.0058315f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_148 C1 Y 0.0422619f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_149 N_C1_c_189_n Y 0.010919f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_150 N_C1_M1003_g Y 0.0164585f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_151 C1 Y 0.0270124f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_152 N_C1_c_189_n Y 0.00933279f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_153 C1 Y 0.0254259f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_154 N_C1_c_189_n Y 0.00565168f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_155 N_C1_M1003_g Y 0.00578802f $X=2.575 $Y=2.165 $X2=0 $Y2=0
cc_156 N_C1_M1006_g N_VGND_c_305_n 0.00357668f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_157 N_C1_M1006_g N_VGND_c_306_n 0.00625597f $X=2.575 $Y=0.445 $X2=0 $Y2=0
cc_158 N_VPWR_c_215_n A_138_369# 0.0057299f $X=0.405 $Y=1.995 $X2=-0.19
+ $Y2=-0.24
cc_159 N_VPWR_c_213_n A_138_369# 0.00742451f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_160 N_VPWR_c_213_n A_222_369# 0.00636867f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_161 N_VPWR_c_213_n N_Y_M1009_d 0.00362055f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_c_213_n N_Y_M1003_d 0.00250309f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_216_n Y 7.78914e-19 $X=2.315 $Y=1.995 $X2=0 $Y2=0
cc_164 N_VPWR_c_217_n Y 0.0343869f $X=2.15 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_c_213_n Y 0.0206517f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_166 N_VPWR_c_216_n Y 0.0279323f $X=2.315 $Y=1.995 $X2=0 $Y2=0
cc_167 N_VPWR_c_216_n Y 0.0281112f $X=2.315 $Y=1.995 $X2=0 $Y2=0
cc_168 N_VPWR_c_219_n Y 0.032253f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_c_213_n Y 0.0186012f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_170 Y N_VGND_c_305_n 0.0125006f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_171 Y N_VGND_c_305_n 0.0303492f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_172 N_Y_M1006_d N_VGND_c_306_n 0.00226544f $X=2.65 $Y=0.235 $X2=0 $Y2=0
cc_173 Y N_VGND_c_306_n 0.0075842f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_174 Y N_VGND_c_306_n 0.0179634f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_175 N_VGND_c_306_n N_A_138_47#_M1005_d 0.00412745f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_176 N_VGND_c_306_n N_A_138_47#_M1004_d 0.0133231f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_177 N_VGND_c_303_n N_A_138_47#_c_362_n 0.0112554f $X=1.08 $Y=0 $X2=0 $Y2=0
cc_178 N_VGND_c_306_n N_A_138_47#_c_362_n 0.00644035f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_179 N_VGND_c_303_n N_A_138_47#_c_344_n 0.00273399f $X=1.08 $Y=0 $X2=0 $Y2=0
cc_180 N_VGND_c_304_n N_A_138_47#_c_344_n 0.020154f $X=1.245 $Y=0.36 $X2=0 $Y2=0
cc_181 N_VGND_c_305_n N_A_138_47#_c_344_n 0.00273399f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_c_306_n N_A_138_47#_c_344_n 0.00972546f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_c_305_n N_A_138_47#_c_358_n 0.011459f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_184 N_VGND_c_306_n N_A_138_47#_c_358_n 0.00644035f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_306_n A_458_47# 0.00706721f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__or4bb_1.spice
* Created: Thu Aug 27 14:44:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or4bb_1.pex.spice"
.subckt sky130_fd_sc_hd__or4bb_1  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_N_M1008_g N_A_27_410#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1092 PD=0.715 PS=1.36 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_205_93#_M1009_d N_D_N_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.06195 PD=1.36 PS=0.715 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_311_413#_M1003_d N_A_205_93#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.05985 AS=0.1092 PD=0.705 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_27_410#_M1006_g N_A_311_413#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.05985 PD=0.69 PS=0.705 NRD=0 NRS=2.856 M=1 R=2.8
+ SA=75000.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_A_311_413#_M1007_d N_B_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_311_413#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0567 PD=0.777196 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_311_413#_M1000_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.123773 PD=1.85 PS=1.2028 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_C_N_M1011_g N_A_27_410#_M1011_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.122612 AS=0.1092 PD=1.32 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_205_93#_M1013_d N_D_N_M1013_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.122612 PD=1.4 PS=1.32 NRD=0 NRS=111.128 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_393_413# N_A_205_93#_M1005_g N_A_311_413#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1215 AS=0.1092 PD=1.33 PS=1.36 NRD=109.887 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_489_297# N_A_27_410#_M1004_g A_393_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1215 PD=0.63 PS=1.33 NRD=23.443 NRS=109.887 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 A_561_297# N_B_M1001_g A_489_297# VPB PHIGHVT L=0.15 W=0.42 AD=0.05985
+ AS=0.0441 PD=0.705 PS=0.63 NRD=41.0351 NRS=23.443 M=1 R=2.8 SA=75000.5
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_561_297# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0876972 AS=0.05985 PD=0.792676 PS=0.705 NRD=72.1217 NRS=41.0351 M=1 R=2.8
+ SA=75001 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_311_413#_M1002_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1
+ AD=0.275 AS=0.208803 PD=2.55 PS=1.88732 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
c_92 VPB 0 1.14153e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__or4bb_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__and4_1.pxi.spice
* Created: Thu Aug 27 14:08:20 2020
* 
x_PM_SKY130_FD_SC_HD__AND4_1%A N_A_M1008_g N_A_M1005_g A N_A_c_62_n
+ PM_SKY130_FD_SC_HD__AND4_1%A
x_PM_SKY130_FD_SC_HD__AND4_1%B N_B_M1003_g N_B_M1004_g B B N_B_c_92_n
+ PM_SKY130_FD_SC_HD__AND4_1%B
x_PM_SKY130_FD_SC_HD__AND4_1%C N_C_M1001_g N_C_M1000_g C C C N_C_c_128_n
+ PM_SKY130_FD_SC_HD__AND4_1%C
x_PM_SKY130_FD_SC_HD__AND4_1%D N_D_M1006_g N_D_M1007_g D N_D_c_162_n
+ PM_SKY130_FD_SC_HD__AND4_1%D
x_PM_SKY130_FD_SC_HD__AND4_1%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1005_d
+ N_A_27_47#_M1000_d N_A_27_47#_c_195_n N_A_27_47#_M1002_g N_A_27_47#_M1009_g
+ N_A_27_47#_c_196_n N_A_27_47#_c_201_n N_A_27_47#_c_202_n N_A_27_47#_c_203_n
+ N_A_27_47#_c_204_n N_A_27_47#_c_205_n N_A_27_47#_c_215_n N_A_27_47#_c_206_n
+ N_A_27_47#_c_207_n N_A_27_47#_c_197_n N_A_27_47#_c_198_n
+ PM_SKY130_FD_SC_HD__AND4_1%A_27_47#
x_PM_SKY130_FD_SC_HD__AND4_1%VPWR N_VPWR_M1005_s N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n VPWR
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_280_n N_VPWR_c_289_n
+ N_VPWR_c_290_n PM_SKY130_FD_SC_HD__AND4_1%VPWR
x_PM_SKY130_FD_SC_HD__AND4_1%X N_X_M1002_d N_X_M1009_d X X X X X X X N_X_c_327_n
+ X PM_SKY130_FD_SC_HD__AND4_1%X
x_PM_SKY130_FD_SC_HD__AND4_1%VGND N_VGND_M1006_d N_VGND_c_348_n VGND
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n
+ PM_SKY130_FD_SC_HD__AND4_1%VGND
cc_1 VNB N_A_M1008_g 0.0335276f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A 0.0241094f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_c_62_n 0.0358837f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_B_M1003_g 0.0289451f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_5 VNB B 0.00436529f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_B_c_92_n 0.022258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_C_M1001_g 0.0295654f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_8 VNB C 0.00405215f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_9 VNB N_C_c_128_n 0.0211841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_D_M1006_g 0.0327756f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_11 VNB D 0.00552985f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB N_D_c_162_n 0.0240404f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_13 VNB N_A_27_47#_c_195_n 0.022188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_196_n 0.00423441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_197_n 0.00176185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_198_n 0.0332007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_280_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0248614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_327_n 0.0203838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_348_n 0.007123f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_21 VNB N_VGND_c_349_n 0.0651496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_350_n 0.0181367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_351_n 0.180805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_352_n 0.00519339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A_M1005_g 0.0542317f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_26 VPB A 0.0375855f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_27 VPB N_A_c_62_n 0.0116644f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_28 VPB N_B_M1004_g 0.0535426f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_29 VPB B 0.00197498f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_30 VPB N_B_c_92_n 0.00452167f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_C_M1000_g 0.0514578f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_32 VPB C 0.00151186f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_33 VPB N_C_c_128_n 0.00444518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_D_M1007_g 0.0582549f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_35 VPB D 2.17214e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_36 VPB N_D_c_162_n 0.00533442f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_37 VPB N_A_27_47#_M1009_g 0.0244277f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_38 VPB N_A_27_47#_c_196_n 0.00182681f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_201_n 0.00802631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_202_n 0.0141766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_203_n 0.00876314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_204_n 0.00479623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_205_n 0.00196007f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_206_n 0.00907375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_207_n 0.00580186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_198_n 0.00945264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_281_n 0.0101372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_282_n 0.0120325f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_49 VPB N_VPWR_c_283_n 0.012113f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_284_n 0.0055866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_285_n 0.0169225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_286_n 0.0262431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_287_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_280_n 0.0429404f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_289_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_290_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB X 0.0366158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB X 0.0105533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 N_A_M1008_g N_B_M1003_g 0.0246474f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_B_M1004_g 0.0269783f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_61 N_A_M1008_g B 9.50824e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_62 N_A_c_62_n N_B_c_92_n 0.0246474f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_M1008_g N_A_27_47#_c_196_n 0.013587f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_A_27_47#_c_196_n 0.00345914f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_65 A N_A_27_47#_c_196_n 0.0522899f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A_c_62_n N_A_27_47#_c_196_n 0.00830241f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_M1005_g N_A_27_47#_c_201_n 0.00412063f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_68 A N_A_27_47#_c_201_n 0.0232492f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_M1008_g N_A_27_47#_c_215_n 0.0130729f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_70 A N_A_27_47#_c_215_n 0.0123303f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_c_62_n N_A_27_47#_c_215_n 0.00201045f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_A_27_47#_c_206_n 0.00703313f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_73 A N_A_27_47#_c_206_n 0.0139295f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 A N_VPWR_M1005_s 0.00226676f $X=0.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_75 N_A_M1005_g N_VPWR_c_282_n 0.00909987f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_76 A N_VPWR_c_282_n 0.0188536f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_M1005_g N_VPWR_c_285_n 0.0046653f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_VPWR_c_280_n 0.00810316f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_79 A N_VPWR_c_280_n 0.00141964f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_M1008_g N_VGND_c_349_n 0.00357877f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_M1008_g N_VGND_c_351_n 0.00625807f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_82 A N_VGND_c_351_n 0.0038518f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_C_M1001_g 0.0256661f $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_84 B N_C_M1001_g 0.00712225f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_85 N_B_M1004_g N_C_M1000_g 0.0295302f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_86 N_B_M1003_g C 5.58864e-19 $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_87 B C 0.0725053f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_88 N_B_c_92_n C 3.10814e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_92_n N_C_c_128_n 0.015329f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_M1003_g N_A_27_47#_c_196_n 0.00476538f $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_A_27_47#_c_196_n 0.00336034f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_92 B N_A_27_47#_c_196_n 0.0459143f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_93 N_B_M1004_g N_A_27_47#_c_201_n 0.00822678f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_94 N_B_M1004_g N_A_27_47#_c_202_n 0.0158289f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_95 B N_A_27_47#_c_202_n 0.0278359f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_96 N_B_c_92_n N_A_27_47#_c_202_n 0.00216998f $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_A_27_47#_c_215_n 0.00423688f $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_98 B N_A_27_47#_c_215_n 0.014844f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_99 N_B_c_92_n N_A_27_47#_c_206_n 4.83855e-19 $X=0.97 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B_M1004_g N_VPWR_c_282_n 5.02781e-19 $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_101 N_B_M1004_g N_VPWR_c_283_n 0.00377488f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_102 N_B_M1004_g N_VPWR_c_285_n 0.00585385f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_VPWR_c_280_n 0.0109266f $X=0.97 $Y=2.275 $X2=0 $Y2=0
cc_104 B A_197_47# 0.00599816f $X=1.065 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_105 N_B_M1003_g N_VGND_c_349_n 0.00448953f $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_106 B N_VGND_c_349_n 0.013239f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_107 N_B_M1003_g N_VGND_c_351_n 0.00756059f $X=0.91 $Y=0.445 $X2=0 $Y2=0
cc_108 B N_VGND_c_351_n 0.0121789f $X=1.065 $Y=0.425 $X2=0 $Y2=0
cc_109 N_C_M1001_g N_D_M1006_g 0.0312763f $X=1.44 $Y=0.445 $X2=0 $Y2=0
cc_110 C N_D_M1006_g 0.00652967f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_111 N_C_M1000_g N_D_M1007_g 0.0381082f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_112 N_C_M1001_g D 5.6497e-19 $X=1.44 $Y=0.445 $X2=0 $Y2=0
cc_113 C D 0.0718202f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_114 N_C_c_128_n D 3.26806e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_115 N_C_c_128_n N_D_c_162_n 0.0204483f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_M1000_g N_A_27_47#_c_202_n 0.0154362f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_117 C N_A_27_47#_c_202_n 0.0125111f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_118 N_C_c_128_n N_A_27_47#_c_202_n 0.00217887f $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_119 N_C_M1000_g N_A_27_47#_c_203_n 0.00813665f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_120 C N_A_27_47#_c_207_n 0.0123056f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_121 N_C_c_128_n N_A_27_47#_c_207_n 4.35311e-19 $X=1.5 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C_M1000_g N_VPWR_c_283_n 0.0050897f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_123 N_C_M1000_g N_VPWR_c_286_n 0.00585385f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_124 N_C_M1000_g N_VPWR_c_280_n 0.0107669f $X=1.49 $Y=2.275 $X2=0 $Y2=0
cc_125 C A_303_47# 0.00458281f $X=1.525 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_126 N_C_M1001_g N_VGND_c_349_n 0.00448323f $X=1.44 $Y=0.445 $X2=0 $Y2=0
cc_127 C N_VGND_c_349_n 0.0113736f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_128 N_C_M1001_g N_VGND_c_351_n 0.00765234f $X=1.44 $Y=0.445 $X2=0 $Y2=0
cc_129 C N_VGND_c_351_n 0.0103942f $X=1.525 $Y=0.425 $X2=0 $Y2=0
cc_130 N_D_M1006_g N_A_27_47#_c_195_n 0.00937516f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_131 D N_A_27_47#_c_195_n 0.00269728f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_132 N_D_M1007_g N_A_27_47#_M1009_g 0.0153486f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_133 N_D_M1007_g N_A_27_47#_c_203_n 0.00761453f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_134 N_D_M1007_g N_A_27_47#_c_204_n 0.0179779f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_135 D N_A_27_47#_c_204_n 0.0218354f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_136 N_D_c_162_n N_A_27_47#_c_204_n 0.00381149f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_137 N_D_M1007_g N_A_27_47#_c_205_n 0.00352692f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_138 D N_A_27_47#_c_197_n 0.0186662f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_139 N_D_c_162_n N_A_27_47#_c_197_n 8.48156e-19 $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_140 D N_A_27_47#_c_198_n 0.00251865f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_141 N_D_c_162_n N_A_27_47#_c_198_n 0.0185899f $X=1.98 $Y=1.16 $X2=0 $Y2=0
cc_142 N_D_M1007_g N_VPWR_c_284_n 0.00906378f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_143 N_D_M1007_g N_VPWR_c_286_n 0.00585385f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_144 N_D_M1007_g N_VPWR_c_280_n 0.0115579f $X=1.92 $Y=2.275 $X2=0 $Y2=0
cc_145 D N_VGND_M1006_d 0.00441165f $X=1.985 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_146 N_D_M1006_g N_VGND_c_348_n 0.0057931f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_147 D N_VGND_c_348_n 0.0401038f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_148 N_D_M1006_g N_VGND_c_349_n 0.00447066f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_149 D N_VGND_c_349_n 0.0105628f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_150 N_D_M1006_g N_VGND_c_351_n 0.00810262f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_151 D N_VGND_c_351_n 0.00972626f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_204_n N_VPWR_M1007_d 0.0220757f $X=2.37 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_201_n N_VPWR_c_283_n 0.0101331f $X=0.72 $Y=2.3 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_202_n N_VPWR_c_283_n 0.0211463f $X=1.58 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_203_n N_VPWR_c_283_n 0.0114393f $X=1.705 $Y=2.3 $X2=0 $Y2=0
cc_156 N_A_27_47#_M1009_g N_VPWR_c_284_n 0.00908063f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_203_n N_VPWR_c_284_n 0.0165215f $X=1.705 $Y=2.3 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_204_n N_VPWR_c_284_n 0.0280671f $X=2.37 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_198_n N_VPWR_c_284_n 8.55454e-19 $X=2.75 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_201_n N_VPWR_c_285_n 0.0170214f $X=0.72 $Y=2.3 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_203_n N_VPWR_c_286_n 0.0145827f $X=1.705 $Y=2.3 $X2=0 $Y2=0
cc_162 N_A_27_47#_M1009_g N_VPWR_c_287_n 0.00541359f $X=2.75 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1005_d N_VPWR_c_280_n 0.00626597f $X=0.545 $Y=2.065 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1000_d N_VPWR_c_280_n 0.00327378f $X=1.565 $Y=2.065 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_M1009_g N_VPWR_c_280_n 0.0113018f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_201_n N_VPWR_c_280_n 0.00955092f $X=0.72 $Y=2.3 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_203_n N_VPWR_c_280_n 0.00955092f $X=1.705 $Y=2.3 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_195_n X 0.0186821f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_205_n X 0.0116249f $X=2.527 $Y=1.495 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_197_n X 0.018994f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_195_n N_X_c_327_n 0.00730409f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_27_47#_M1009_g X 0.00440054f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_196_n A_109_47# 8.25779e-19 $X=0.58 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_27_47#_c_215_n A_109_47# 0.00429836f $X=0.58 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_27_47#_c_195_n N_VGND_c_348_n 0.00902138f $X=2.75 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_204_n N_VGND_c_348_n 4.22529e-19 $X=2.37 $Y=1.58 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_197_n N_VGND_c_348_n 0.0199489f $X=2.535 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_198_n N_VGND_c_348_n 0.00566811f $X=2.75 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_215_n N_VGND_c_349_n 0.0289623f $X=0.58 $Y=0.42 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_195_n N_VGND_c_350_n 0.00542953f $X=2.75 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1008_s N_VGND_c_351_n 0.0022878f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_195_n N_VGND_c_351_n 0.0113045f $X=2.75 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_215_n N_VGND_c_351_n 0.0179555f $X=0.58 $Y=0.42 $X2=0 $Y2=0
cc_184 N_VPWR_c_280_n N_X_M1009_d 0.00209319f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_185 N_VPWR_c_287_n X 0.0216305f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_186 N_VPWR_c_280_n X 0.0127342f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_187 N_X_c_327_n N_VGND_c_350_n 0.0172989f $X=2.96 $Y=0.38 $X2=0 $Y2=0
cc_188 N_X_M1002_d N_VGND_c_351_n 0.00211564f $X=2.825 $Y=0.235 $X2=0 $Y2=0
cc_189 N_X_c_327_n N_VGND_c_351_n 0.0125287f $X=2.96 $Y=0.38 $X2=0 $Y2=0
cc_190 A_109_47# N_VGND_c_351_n 0.00822242f $X=0.545 $Y=0.235 $X2=0.72 $Y2=2.3
cc_191 A_197_47# N_VGND_c_351_n 0.00770534f $X=0.985 $Y=0.235 $X2=0 $Y2=0
cc_192 A_303_47# N_VGND_c_351_n 0.0072757f $X=1.515 $Y=0.235 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__nand2b_2.spice
* Created: Thu Aug 27 14:29:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand2b_2.spice.pex"
.subckt sky130_fd_sc_hd__nand2b_2  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_N_M1009_g N_A_27_93#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.194 AS=0.1092 PD=1.95 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_27_93#_M1002_g N_A_229_47#_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1002_d N_A_27_93#_M1005_g N_A_229_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1007 N_A_229_47#_M1005_s N_B_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_229_47#_M1008_d N_B_M1008_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_N_M1004_g N_A_27_93#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0868394 AS=0.1092 PD=0.792676 PS=1.36 NRD=71.1761 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1004_d N_A_27_93#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.206761 AS=0.165 PD=1.88732 PS=1.33 NRD=0 NRS=4.9053 M=1 R=6.66667
+ SA=75000.4 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_93#_M1006_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.335 AS=0.165 PD=1.67 PS=1.33 NRD=0 NRS=4.9053 M=1 R=6.66667 SA=75000.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1006_d N_B_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.335
+ AS=0.135 PD=1.67 PS=1.27 NRD=10.8153 NRS=0 M=1 R=6.66667 SA=75001.7 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1 AD=0.275
+ AS=0.135 PD=2.55 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.1 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_37 VNB 0 5.82644e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hd__nand2b_2.spice.SKY130_FD_SC_HD__NAND2B_2.pxi"
*
.ends
*
*

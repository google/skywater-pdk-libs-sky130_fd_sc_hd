* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hd__macro_sparecell VGND VNB VPB VPWR LO
*.PININFO VGND:I VNB:I VPB:I VPWR:I LO:O
XI1 net59 LO VGND VNB VPB VPWR / scs8hd_conb_1
XI6 nor2right invright VGND VNB VPB VPWR / scs8hd_inv_2
XI7 nor2left invleft VGND VNB VPB VPWR / scs8hd_inv_2
XI4 nd2right nd2right nor2right VGND VNB VPB VPWR / scs8hd_nor2_2
XI5 nd2left nd2left nor2left VGND VNB VPB VPWR / scs8hd_nor2_2
XI2 LO LO nd2right VGND VNB VPB VPWR / scs8hd_nand2_2
XI3 LO LO nd2left VGND VNB VPB VPWR / scs8hd_nand2_2
.ENDS sky130_fd_sc_hd__macro_sparecell

* File: sky130_fd_sc_hd__o21ai_2.spice
* Created: Thu Aug 27 14:35:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ai_2.spice.pex"
.subckt sky130_fd_sc_hd__o21ai_2  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_A_29_47#_M1009_d N_A1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.091 PD=1.83 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 N_A_29_47#_M1000_d N_A2_M1000_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002 A=0.0975 P=1.6 MULT=1
MM1004 N_A_29_47#_M1000_d N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.12675 PD=0.93 PS=1.04 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_29_47#_M1011_d N_A1_M1011_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.12675 PD=0.93 PS=1.04 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75001.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_29_47#_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1002_d N_B1_M1007_g N_A_29_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_112_297#_M1003_d N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1005 N_A_112_297#_M1003_d N_A2_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75002
+ A=0.15 P=2.3 MULT=1
MM1010 N_A_112_297#_M1010_d N_A2_M1010_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.14 PD=1.35 PS=1.28 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_112_297#_M1010_d N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.175 AS=0.16 PD=1.35 PS=1.32 NRD=3.9203 NRS=2.9353 M=1 R=6.66667
+ SA=75001.5 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1008_s N_B1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=4.9053 NRS=0 M=1 R=6.66667 SA=75002 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.265
+ AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hd__o21ai_2.spice.SKY130_FD_SC_HD__O21AI_2.pxi"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_hd__and3_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
M1000 a_27_47# B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=3.9785e+11p ps=4.05e+06u
M1001 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.633e+11p ps=2.28e+06u
M1002 a_181_47# B a_109_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1003 VGND C a_181_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1006 a_109_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1007 VPWR C a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


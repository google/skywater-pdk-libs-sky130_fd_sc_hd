* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X3 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X4 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X15 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends

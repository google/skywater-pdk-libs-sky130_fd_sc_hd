* File: sky130_fd_sc_hd__nor3b_4.spice
* Created: Thu Aug 27 14:32:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nor3b_4.pex.spice"
.subckt sky130_fd_sc_hd__nor3b_4  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_C_N_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1017_d N_A_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1010_d N_A_M1016_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_A_M1021_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1011 N_Y_M1002_d N_B_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1012_d N_B_M1012_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1025 N_Y_M1012_d N_B_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1025_s N_A_27_47#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.5
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_27_47#_M1005_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1005_d N_A_27_47#_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_27_47#_M1009_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_C_N_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1004_d N_A_M1014_g N_A_197_297#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_A_197_297#_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1018_d N_A_M1019_g N_A_197_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_A_197_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_197_297#_M1000_d N_B_M1000_g N_A_555_297#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.1 A=0.15 P=2.3 MULT=1
MM1003 N_A_197_297#_M1000_d N_B_M1003_g N_A_555_297#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1006 N_A_197_297#_M1006_d N_B_M1006_g N_A_555_297#_M1003_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.3 A=0.15 P=2.3 MULT=1
MM1013 N_A_197_297#_M1006_d N_B_M1013_g N_A_555_297#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1015 N_Y_M1015_d N_A_27_47#_M1015_g N_A_555_297#_M1013_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.4 A=0.15 P=2.3 MULT=1
MM1020 N_Y_M1015_d N_A_27_47#_M1020_g N_A_555_297#_M1020_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1023 N_Y_M1023_d N_A_27_47#_M1023_g N_A_555_297#_M1020_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1024 N_Y_M1023_d N_A_27_47#_M1024_g N_A_555_297#_M1024_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.1
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX26_noxref VNB VPB NWDIODE A=11.6844 P=17.77
*
.include "sky130_fd_sc_hd__nor3b_4.pxi.spice"
*
.ends
*
*

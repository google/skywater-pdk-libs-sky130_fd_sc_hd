# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.12000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095000 1.020000 7.745000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.960000 1.020000 9.990000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.020000 5.650000 1.275000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.020000 3.745000 1.275000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 1.020000 1.845000 1.275000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.009500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 7.620000 0.785000 ;
        RECT 0.145000 0.785000 0.320000 1.475000 ;
        RECT 0.145000 1.475000 1.720000 1.655000 ;
        RECT 0.530000 1.655000 1.720000 1.685000 ;
        RECT 0.530000 1.685000 0.860000 2.085000 ;
        RECT 0.615000 0.455000 0.790000 0.615000 ;
        RECT 1.390000 1.685000 1.720000 2.085000 ;
        RECT 1.460000 0.455000 1.650000 0.615000 ;
        RECT 2.400000 0.455000 2.590000 0.615000 ;
        RECT 3.260000 0.455000 3.510000 0.615000 ;
        RECT 4.180000 0.455000 4.420000 0.615000 ;
        RECT 5.090000 0.455000 5.275000 0.615000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.120000 0.085000 ;
        RECT 0.115000  0.085000  0.445000 0.445000 ;
        RECT 0.960000  0.085000  1.290000 0.445000 ;
        RECT 1.820000  0.085000  2.230000 0.445000 ;
        RECT 2.760000  0.085000  3.090000 0.445000 ;
        RECT 3.680000  0.085000  4.010000 0.445000 ;
        RECT 4.590000  0.085000  4.920000 0.445000 ;
        RECT 5.445000  0.085000  5.780000 0.445000 ;
        RECT 8.245000  0.085000  8.575000 0.445000 ;
        RECT 9.105000  0.085000  9.435000 0.445000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.120000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.120000 2.805000 ;
        RECT 6.220000 1.785000  6.550000 2.635000 ;
        RECT 7.080000 1.805000  7.410000 2.635000 ;
        RECT 8.080000 1.895000  8.410000 2.635000 ;
        RECT 9.030000 1.915000  9.360000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.120000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.100000 1.835000 0.360000 2.255000 ;
      RECT 0.100000 2.255000 3.870000 2.445000 ;
      RECT 1.030000 1.855000 1.220000 2.255000 ;
      RECT 1.890000 1.855000 2.080000 2.255000 ;
      RECT 2.250000 1.475000 5.680000 1.655000 ;
      RECT 2.250000 1.655000 3.440000 1.685000 ;
      RECT 2.250000 1.685000 2.580000 2.085000 ;
      RECT 2.750000 1.855000 2.940000 2.255000 ;
      RECT 3.110000 1.685000 3.440000 2.085000 ;
      RECT 3.610000 1.835000 3.870000 2.255000 ;
      RECT 4.060000 1.835000 4.320000 2.255000 ;
      RECT 4.060000 2.255000 5.180000 2.275000 ;
      RECT 4.060000 2.275000 6.050000 2.445000 ;
      RECT 4.490000 1.655000 5.680000 1.685000 ;
      RECT 4.490000 1.685000 4.820000 2.085000 ;
      RECT 4.990000 1.855000 5.180000 2.255000 ;
      RECT 5.350000 1.685000 5.680000 2.085000 ;
      RECT 5.860000 1.445000 9.770000 1.615000 ;
      RECT 5.860000 1.615000 6.050000 2.275000 ;
      RECT 5.980000 0.275000 8.075000 0.445000 ;
      RECT 6.720000 1.615000 6.910000 2.315000 ;
      RECT 7.580000 1.615000 9.770000 1.665000 ;
      RECT 7.580000 1.665000 7.910000 2.315000 ;
      RECT 7.885000 0.445000 8.075000 0.615000 ;
      RECT 7.885000 0.615000 9.865000 0.785000 ;
      RECT 8.580000 1.665000 9.770000 1.670000 ;
      RECT 8.580000 1.670000 8.840000 2.290000 ;
      RECT 8.745000 0.300000 8.935000 0.615000 ;
      RECT 9.530000 1.670000 9.770000 2.260000 ;
      RECT 9.605000 0.290000 9.865000 0.615000 ;
  END
END sky130_fd_sc_hd__a2111oi_4
END LIBRARY

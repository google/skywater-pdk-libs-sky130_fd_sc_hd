* File: sky130_fd_sc_hd__and4b_1.pex.spice
* Created: Tue Sep  1 18:58:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4B_1%A_N 3 7 9 10 17
c33 17 0 1.66235e-19 $X=0.47 $Y=1.16
r34 14 17 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.47 $Y2=1.16
r35 9 10 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.267 $Y=1.16
+ $X2=0.267 $Y2=1.53
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r37 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r38 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=2.275
r39 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r40 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%A_27_47# 1 2 7 9 11 13 15 18 22 24 25 26 27
+ 29 31 35
c77 26 0 1.66235e-19 $X=0.63 $Y=1.93
r78 36 38 78.4908 $w=2.18e-07 $l=3.55e-07 $layer=POLY_cond $X=0.895 $Y=1.16
+ $X2=0.895 $Y2=0.805
r79 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.895
+ $Y=1.16 $X2=0.895 $Y2=1.16
r80 32 35 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.895 $Y2=1.16
r81 30 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=1.325
+ $X2=0.715 $Y2=1.16
r82 30 31 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.715 $Y=1.325
+ $X2=0.715 $Y2=1.845
r83 29 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=0.995
+ $X2=0.715 $Y2=1.16
r84 28 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.715 $Y=0.825
+ $X2=0.715 $Y2=0.995
r85 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=1.93
+ $X2=0.715 $Y2=1.845
r86 26 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.63 $Y=1.93
+ $X2=0.345 $Y2=1.93
r87 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=0.74
+ $X2=0.715 $Y2=0.825
r88 24 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.63 $Y=0.74
+ $X2=0.345 $Y2=0.74
r89 20 27 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=2.015
+ $X2=0.345 $Y2=1.93
r90 20 22 18.0623 $w=1.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.257 $Y=2.015
+ $X2=0.257 $Y2=2.3
r91 16 25 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.655
+ $X2=0.345 $Y2=0.74
r92 16 18 14.8935 $w=1.73e-07 $l=2.35e-07 $layer=LI1_cond $X=0.257 $Y=0.655
+ $X2=0.257 $Y2=0.42
r93 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.41 $Y=0.73 $X2=1.41
+ $Y2=0.445
r94 12 38 11.5617 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.03 $Y=0.805
+ $X2=0.895 $Y2=0.805
r95 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=0.805
+ $X2=1.41 $Y2=0.73
r96 11 12 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.335 $Y=0.805
+ $X2=1.03 $Y2=0.805
r97 7 36 41.2111 $w=2.18e-07 $l=1.67481e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.895 $Y2=1.16
r98 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=2.275
r99 2 22 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r100 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%B 3 7 9 10 11 12 22
r38 20 22 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=1.655 $Y=1.27
+ $X2=1.77 $Y2=1.27
r39 17 20 32.2152 $w=2.7e-07 $l=1.45e-07 $layer=POLY_cond $X=1.51 $Y=1.27
+ $X2=1.655 $Y2=1.27
r40 11 12 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.66 $Y=1.19 $X2=1.66
+ $Y2=1.53
r41 11 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.27 $X2=1.655 $Y2=1.27
r42 10 11 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.66 $Y=0.85 $X2=1.66
+ $Y2=1.19
r43 9 10 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.66 $Y=0.51 $X2=1.66
+ $Y2=0.85
r44 5 22 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.77 $Y=1.135
+ $X2=1.77 $Y2=1.27
r45 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.77 $Y=1.135 $X2=1.77
+ $Y2=0.445
r46 1 17 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.51 $Y=1.405
+ $X2=1.51 $Y2=1.27
r47 1 3 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.51 $Y=1.405 $X2=1.51
+ $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%C 3 7 9 10 11 12 18
r38 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.16
+ $X2=2.21 $Y2=1.325
r39 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.16
+ $X2=2.21 $Y2=0.995
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.16 $X2=2.21 $Y2=1.16
r41 11 12 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=1.19
+ $X2=2.16 $Y2=1.53
r42 11 19 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.16 $Y=1.19 $X2=2.16
+ $Y2=1.16
r43 10 19 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.16 $Y=0.85
+ $X2=2.16 $Y2=1.16
r44 9 10 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=0.51 $X2=2.16
+ $Y2=0.85
r45 7 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.27 $Y=2.275
+ $X2=2.27 $Y2=1.325
r46 3 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.27 $Y=0.445
+ $X2=2.27 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%D 3 7 9 10 11 16
c42 16 0 1.99282e-19 $X=2.69 $Y=1.16
r43 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=1.325
r44 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=0.995
r45 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r46 10 11 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.655 $Y=1.19
+ $X2=2.655 $Y2=1.53
r47 10 17 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=2.655 $Y=1.19
+ $X2=2.655 $Y2=1.16
r48 9 17 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=2.655 $Y=0.85
+ $X2=2.655 $Y2=1.16
r49 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.325
r50 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.71 $Y=0.445
+ $X2=2.71 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%A_193_413# 1 2 3 12 15 18 21 23 27 29 32 34
+ 37 38 42 43 46
c93 38 0 1.99282e-19 $X=2.525 $Y=1.96
r94 43 47 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.17 $Y2=1.325
r95 43 46 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.17 $Y2=0.995
r96 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.16 $X2=3.17 $Y2=1.16
r97 39 42 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.08 $Y=1.16 $X2=3.17
+ $Y2=1.16
r98 34 36 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0.42
+ $X2=1.205 $Y2=0.585
r99 31 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.16
r100 31 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.08 $Y=1.325
+ $X2=3.08 $Y2=1.875
r101 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.96
+ $X2=2.525 $Y2=1.96
r102 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=1.96
+ $X2=3.08 $Y2=1.875
r103 29 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.995 $Y=1.96
+ $X2=2.61 $Y2=1.96
r104 25 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=2.045
+ $X2=2.525 $Y2=1.96
r105 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.525 $Y=2.045
+ $X2=2.525 $Y2=2.3
r106 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=1.96
+ $X2=1.235 $Y2=1.96
r107 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=1.96
+ $X2=2.525 $Y2=1.96
r108 23 24 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=2.44 $Y=1.96
+ $X2=1.32 $Y2=1.96
r109 19 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.045
+ $X2=1.235 $Y2=1.96
r110 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.235 $Y=2.045
+ $X2=1.235 $Y2=2.3
r111 18 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=1.875
+ $X2=1.235 $Y2=1.96
r112 18 36 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=1.235 $Y=1.875
+ $X2=1.235 $Y2=0.585
r113 15 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.21 $Y=1.985
+ $X2=3.21 $Y2=1.325
r114 12 46 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.56
+ $X2=3.21 $Y2=0.995
r115 3 27 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=2.065 $X2=2.525 $Y2=2.3
r116 2 21 600 $w=1.7e-07 $l=3.69256e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=2.065 $X2=1.235 $Y2=2.3
r117 1 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%VPWR 1 2 3 12 18 20 22 27 34 35 38 43 49 51
r60 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 47 49 9.81967 $w=5.78e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=2.515
+ $X2=2.225 $Y2=2.515
r62 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 45 47 0.20622 $w=5.78e-07 $l=1e-08 $layer=LI1_cond $X=2.06 $Y=2.515 $X2=2.07
+ $Y2=2.515
r64 42 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 41 45 9.27992 $w=5.78e-07 $l=4.5e-07 $layer=LI1_cond $X=1.61 $Y=2.515
+ $X2=2.06 $Y2=2.515
r66 41 43 7.75746 $w=5.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.61 $Y=2.515
+ $X2=1.555 $Y2=2.515
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r69 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 35 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r72 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=2.975 $Y2=2.72
r73 32 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.14 $Y=2.72
+ $X2=3.45 $Y2=2.72
r74 31 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 31 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 30 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.225 $Y2=2.72
r77 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 27 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.975 $Y2=2.72
r79 27 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.81 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 22 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r81 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r82 20 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 20 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r84 16 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.72
r85 16 18 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.975 $Y=2.635
+ $X2=2.975 $Y2=2.31
r86 15 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r87 15 43 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.555 $Y2=2.72
r88 10 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r89 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r90 3 18 600 $w=1.7e-07 $l=3.16938e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.065 $X2=2.975 $Y2=2.31
r91 2 45 300 $w=1.7e-07 $l=5.84808e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=2.065 $X2=2.06 $Y2=2.31
r92 1 12 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%X 1 2 7 9 10 11 12 13 18
r20 12 13 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.465 $Y=1.87
+ $X2=3.465 $Y2=2.21
r21 12 18 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=3.465 $Y=1.87
+ $X2=3.465 $Y2=1.66
r22 11 25 4.67847 $w=3.39e-07 $l=1.3e-07 $layer=LI1_cond $X=3.425 $Y=0.51
+ $X2=3.425 $Y2=0.38
r23 9 18 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.465 $Y=1.625
+ $X2=3.465 $Y2=1.66
r24 9 10 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.465 $Y=1.625
+ $X2=3.465 $Y2=1.495
r25 7 11 13.6456 $w=3.39e-07 $l=3.34813e-07 $layer=LI1_cond $X=3.51 $Y=0.805
+ $X2=3.425 $Y2=0.51
r26 7 10 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.51 $Y=0.805 $X2=3.51
+ $Y2=1.495
r27 2 18 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.485 $X2=3.42 $Y2=1.66
r28 1 25 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND4B_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r57 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r59 33 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r60 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r61 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=2.92
+ $Y2=0
r62 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.45
+ $Y2=0
r63 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r64 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r65 26 29 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r66 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r67 25 28 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r68 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r70 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r71 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.92
+ $Y2=0
r72 22 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.53
+ $Y2=0
r73 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r74 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r75 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r78 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.38
r79 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085 $X2=0.68
+ $Y2=0
r80 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r81 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.235 $X2=2.92 $Y2=0.38
r82 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__and2b_4.spice
* Created: Thu Aug 27 14:07:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and2b_4.spice.pex"
.subckt sky130_fd_sc_hd__and2b_4  VNB VPB B A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* B	B
* VPB	VPB
* VNB	VNB
MM1012 A_109_47# N_A_33_199#_M1012_g N_A_27_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.0715 AS=0.169 PD=0.87 PS=1.82 NRD=10.152 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g A_109_47# VNB NSHORT L=0.15 W=0.65 AD=0.1365
+ AS=0.0715 PD=1.07 PS=0.87 NRD=11.988 NRS=10.152 M=1 R=4.33333 SA=75000.6
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.1365 PD=0.93 PS=1.07 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75001.1
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1003_d N_A_27_47#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0.912 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1008_d N_A_27_47#_M1008_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75002
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1008_d N_A_27_47#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.129696 PD=0.93 PS=1.22103 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1004 N_A_33_199#_M1004_d N_A_N_M1004_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0838037 PD=1.37 PS=0.788972 NRD=0 NRS=41.292 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_27_47#_M1010_d N_A_33_199#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_27_47#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.185 AS=0.135 PD=1.37 PS=1.27 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.2 A=0.15 P=2.3 MULT=1
MM1000 N_X_M1000_d N_A_27_47#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.185 PD=1.3 PS=1.37 NRD=4.9053 NRS=7.8603 M=1 R=6.66667 SA=75001.1
+ SB=75001.7 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1000_d N_A_27_47#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.15 AS=0.135 PD=1.3 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.6
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1007 N_X_M1007_d N_A_27_47#_M1007_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002
+ SB=75000.8 A=0.15 P=2.3 MULT=1
MM1013 N_X_M1007_d N_A_27_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.219366 PD=1.27 PS=1.90845 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75000.4 A=0.15 P=2.3 MULT=1
MM1002 N_A_33_199#_M1002_d N_A_N_M1002_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0921338 PD=1.37 PS=0.801549 NRD=0 NRS=77.0861 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
DX14_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_68 VPB 0 1.19177e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__and2b_4.spice.SKY130_FD_SC_HD__AND2B_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__diode_2.pxi.spice
* Created: Thu Aug 27 14:16:11 2020
* 
x_PM_SKY130_FD_SC_HD__DIODE_2%DIODE N_DIODE_D0_noxref_neg DIODE DIODE DIODE
+ DIODE DIODE DIODE N_DIODE_c_6_n PM_SKY130_FD_SC_HD__DIODE_2%DIODE
cc_1 VNB N_DIODE_c_6_n 0.100756f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=0.37
cc_2 VNB VGND 0.111926f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=0.195
cc_3 VNB VPWR 0.0420108f $X=-0.19 $Y=-0.24 $X2=0.155 $Y2=0.195
cc_4 VPB N_DIODE_c_6_n 0.132027f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=0.37
cc_5 VPB VPWR 0.0750482f $X=-0.19 $Y=1.305 $X2=0.155 $Y2=0.195
cc_6 N_DIODE_D0_noxref_neg VGND 0.00601196f $X=0.155 $Y=0.195 $X2=-0.19
+ $Y2=-0.24
cc_7 N_DIODE_c_6_n VGND 0.0815688f $X=0.66 $Y=0.37 $X2=-0.19 $Y2=-0.24
cc_8 N_DIODE_c_6_n VPWR 0.0824348f $X=0.66 $Y=0.37 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__o41ai_2.spice.SKY130_FD_SC_HD__O41AI_2.pxi
* Created: Thu Aug 27 14:42:13 2020
* 
x_PM_SKY130_FD_SC_HD__O41AI_2%B1 N_B1_c_100_n N_B1_M1009_g N_B1_M1002_g
+ N_B1_c_101_n N_B1_M1019_g N_B1_M1015_g B1 N_B1_c_103_n
+ PM_SKY130_FD_SC_HD__O41AI_2%B1
x_PM_SKY130_FD_SC_HD__O41AI_2%A4 N_A4_M1001_g N_A4_M1016_g N_A4_c_144_n
+ N_A4_M1004_g N_A4_M1017_g A4 A4 PM_SKY130_FD_SC_HD__O41AI_2%A4
x_PM_SKY130_FD_SC_HD__O41AI_2%A3 N_A3_c_194_n N_A3_M1010_g N_A3_M1006_g
+ N_A3_c_195_n N_A3_M1011_g N_A3_M1013_g A3 A3 N_A3_c_197_n
+ PM_SKY130_FD_SC_HD__O41AI_2%A3
x_PM_SKY130_FD_SC_HD__O41AI_2%A2 N_A2_c_245_n N_A2_M1005_g N_A2_M1014_g
+ N_A2_c_247_n N_A2_M1007_g N_A2_M1018_g A2 A2 PM_SKY130_FD_SC_HD__O41AI_2%A2
x_PM_SKY130_FD_SC_HD__O41AI_2%A1 N_A1_M1003_g N_A1_M1000_g N_A1_M1012_g
+ N_A1_M1008_g N_A1_c_301_n A1 A1 A1 N_A1_c_303_n PM_SKY130_FD_SC_HD__O41AI_2%A1
x_PM_SKY130_FD_SC_HD__O41AI_2%VPWR N_VPWR_M1002_d N_VPWR_M1015_d N_VPWR_M1000_s
+ N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n
+ N_VPWR_c_348_n VPWR N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_342_n
+ N_VPWR_c_352_n PM_SKY130_FD_SC_HD__O41AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O41AI_2%Y N_Y_M1009_s N_Y_M1002_s N_Y_M1016_s N_Y_c_419_n
+ N_Y_c_415_n N_Y_c_416_n Y Y Y N_Y_c_430_n Y PM_SKY130_FD_SC_HD__O41AI_2%Y
x_PM_SKY130_FD_SC_HD__O41AI_2%A_299_297# N_A_299_297#_M1016_d
+ N_A_299_297#_M1017_d N_A_299_297#_M1013_d N_A_299_297#_c_460_n
+ N_A_299_297#_c_465_n N_A_299_297#_c_461_n N_A_299_297#_c_482_n
+ N_A_299_297#_c_462_n N_A_299_297#_c_463_n N_A_299_297#_c_464_n
+ PM_SKY130_FD_SC_HD__O41AI_2%A_299_297#
x_PM_SKY130_FD_SC_HD__O41AI_2%A_549_297# N_A_549_297#_M1006_s
+ N_A_549_297#_M1014_s N_A_549_297#_c_499_n N_A_549_297#_c_498_n
+ N_A_549_297#_c_502_n N_A_549_297#_c_506_n
+ PM_SKY130_FD_SC_HD__O41AI_2%A_549_297#
x_PM_SKY130_FD_SC_HD__O41AI_2%A_743_297# N_A_743_297#_M1014_d
+ N_A_743_297#_M1018_d N_A_743_297#_M1008_d N_A_743_297#_c_522_n
+ N_A_743_297#_c_546_n N_A_743_297#_c_523_n N_A_743_297#_c_524_n
+ N_A_743_297#_c_525_n N_A_743_297#_c_526_n N_A_743_297#_c_527_n
+ PM_SKY130_FD_SC_HD__O41AI_2%A_743_297#
x_PM_SKY130_FD_SC_HD__O41AI_2%A_27_47# N_A_27_47#_M1009_d N_A_27_47#_M1019_d
+ N_A_27_47#_M1001_d N_A_27_47#_M1010_s N_A_27_47#_M1005_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1012_d N_A_27_47#_c_561_n N_A_27_47#_c_562_n N_A_27_47#_c_580_n
+ N_A_27_47#_c_563_n N_A_27_47#_c_564_n N_A_27_47#_c_565_n N_A_27_47#_c_566_n
+ N_A_27_47#_c_589_n N_A_27_47#_c_567_n N_A_27_47#_c_593_n N_A_27_47#_c_568_n
+ N_A_27_47#_c_569_n N_A_27_47#_c_570_n N_A_27_47#_c_616_n N_A_27_47#_c_571_n
+ N_A_27_47#_c_572_n N_A_27_47#_c_573_n N_A_27_47#_c_574_n N_A_27_47#_c_575_n
+ N_A_27_47#_c_576_n PM_SKY130_FD_SC_HD__O41AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O41AI_2%VGND N_VGND_M1001_s N_VGND_M1004_s N_VGND_M1011_d
+ N_VGND_M1005_s N_VGND_M1003_s N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n
+ N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n
+ VGND N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n
+ PM_SKY130_FD_SC_HD__O41AI_2%VGND
cc_1 VNB N_B1_c_100_n 0.0218118f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_2 VNB N_B1_c_101_n 0.0213711f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1
cc_3 VNB B1 0.00739817f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_B1_c_103_n 0.0577137f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.155
cc_5 VNB N_A4_M1001_g 0.0230908f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_6 VNB N_A4_c_144_n 0.0440469f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_7 VNB N_A4_M1004_g 0.0175655f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.31
cc_8 VNB A4 0.00398645f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_9 VNB N_A3_c_194_n 0.0167892f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_10 VNB N_A3_c_195_n 0.0223573f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1
cc_11 VNB A3 0.0104884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A3_c_197_n 0.0404228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_245_n 0.0210751f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1
cc_14 VNB N_A2_M1014_g 5.70301e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_15 VNB N_A2_c_247_n 0.0678892f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1
cc_16 VNB N_A2_M1018_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_17 VNB A2 0.00147452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A1_M1003_g 0.0175639f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB N_A1_M1000_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A1_M1012_g 0.0238771f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.31
cc_21 VNB N_A1_M1008_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_A1_c_301_n 0.0244845f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.155
cc_23 VNB A1 0.0226217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A1_c_303_n 0.035956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_342_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.00102834f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.155
cc_27 VNB N_A_27_47#_c_561_n 0.00929764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_562_n 0.0186192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_563_n 0.00218672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_564_n 0.00292811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_565_n 0.00950017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_566_n 0.00438747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_567_n 0.00502844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_568_n 0.012193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_569_n 0.00495287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_570_n 0.00217793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_571_n 0.0110652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_572_n 0.0183265f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_573_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_574_n 0.00222758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_c_575_n 0.00273991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_576_n 0.00348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_697_n 0.00784154f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_44 VNB N_VGND_c_698_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_699_n 0.00725923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_700_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_701_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_702_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_703_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_704_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_705_n 0.00448912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_706_n 0.0189035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_707_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_708_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_709_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_710_n 0.0363931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_711_n 0.0229659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_712_n 0.308393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_713_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VPB N_B1_M1002_g 0.0271346f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_61 VPB N_B1_M1015_g 0.0256664f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_62 VPB N_B1_c_103_n 0.0117486f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.155
cc_63 VPB N_A4_M1016_g 0.0266409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A4_c_144_n 0.00808891f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_65 VPB N_A4_M1017_g 0.0196003f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_66 VPB N_A3_M1006_g 0.0191806f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_A3_M1013_g 0.0262448f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_A3_c_197_n 0.00699813f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A2_M1014_g 0.0266417f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_70 VPB N_A2_M1018_g 0.0194911f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_71 VPB N_A1_M1000_g 0.0192639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A1_M1008_g 0.026498f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_73 VPB N_VPWR_c_343_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_74 VPB N_VPWR_c_344_n 0.0426886f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_75 VPB N_VPWR_c_345_n 0.0108458f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_76 VPB N_VPWR_c_346_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_347_n 0.0874296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_348_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_349_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_350_n 0.0208797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_342_n 0.0616801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_352_n 0.00477947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_Y_c_415_n 0.0204941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_Y_c_416_n 0.00223596f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_85 VPB Y 0.0012699f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.155
cc_86 VPB Y 4.31737e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_299_297#_c_460_n 0.00443954f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_88 VPB N_A_299_297#_c_461_n 0.00181821f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_89 VPB N_A_299_297#_c_462_n 0.00672436f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.155
cc_90 VPB N_A_299_297#_c_463_n 0.00290214f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.155
cc_91 VPB N_A_299_297#_c_464_n 0.00463043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_549_297#_c_498_n 0.0119191f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.31
cc_93 VPB N_A_743_297#_c_522_n 0.00321875f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_94 VPB N_A_743_297#_c_523_n 0.00293165f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_95 VPB N_A_743_297#_c_524_n 0.00867926f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.155
cc_96 VPB N_A_743_297#_c_525_n 0.0313172f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_743_297#_c_526_n 0.00854254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_743_297#_c_527_n 0.00223793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 N_B1_c_103_n N_A4_c_144_n 0.00661769f $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_100 N_B1_c_103_n A4 0.00100487f $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_101 N_B1_M1002_g N_VPWR_c_344_n 0.00321781f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_102 B1 N_VPWR_c_344_n 0.0154705f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B1_c_103_n N_VPWR_c_344_n 0.00546397f $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_104 N_B1_M1015_g N_VPWR_c_345_n 0.00321269f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B1_M1002_g N_VPWR_c_349_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_M1015_g N_VPWR_c_349_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B1_M1002_g N_VPWR_c_342_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_108 N_B1_M1015_g N_VPWR_c_342_n 0.0108276f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_109 N_B1_M1002_g N_Y_c_419_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_110 N_B1_M1015_g N_Y_c_419_n 0.0145598f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_111 N_B1_M1015_g N_Y_c_415_n 0.0185401f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_112 N_B1_c_100_n Y 0.00252419f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_113 N_B1_M1002_g Y 0.00334195f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_114 N_B1_c_101_n Y 0.00513102f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_115 N_B1_M1015_g Y 0.00673635f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_116 B1 Y 0.0145749f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_117 N_B1_c_103_n Y 0.0246239f $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_118 N_B1_M1002_g Y 0.00409939f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_119 N_B1_M1015_g Y 9.33329e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_120 N_B1_c_100_n N_Y_c_430_n 0.00389361f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_121 N_B1_c_101_n N_Y_c_430_n 0.00314611f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_122 N_B1_c_100_n N_A_27_47#_c_562_n 4.72894e-19 $X=0.47 $Y=1 $X2=0 $Y2=0
cc_123 B1 N_A_27_47#_c_562_n 0.0194124f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B1_c_103_n N_A_27_47#_c_562_n 0.00581864f $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_125 N_B1_c_100_n N_A_27_47#_c_580_n 0.011676f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_126 N_B1_c_101_n N_A_27_47#_c_580_n 0.0124471f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_127 B1 N_A_27_47#_c_580_n 0.00168026f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_c_103_n N_A_27_47#_c_580_n 2.99017e-19 $X=0.89 $Y=1.155 $X2=0 $Y2=0
cc_129 N_B1_c_101_n N_A_27_47#_c_566_n 4.59762e-19 $X=0.89 $Y=1 $X2=0 $Y2=0
cc_130 N_B1_c_101_n N_VGND_c_697_n 0.00229957f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_131 N_B1_c_100_n N_VGND_c_710_n 0.00357877f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_132 N_B1_c_101_n N_VGND_c_710_n 0.00357877f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_133 N_B1_c_100_n N_VGND_c_712_n 0.00617937f $X=0.47 $Y=1 $X2=0 $Y2=0
cc_134 N_B1_c_101_n N_VGND_c_712_n 0.00655123f $X=0.89 $Y=1 $X2=0 $Y2=0
cc_135 N_A4_M1004_g N_A3_c_194_n 0.0195612f $X=2.25 $Y=0.56 $X2=-0.19 $Y2=-0.24
cc_136 N_A4_M1017_g N_A3_M1006_g 0.0195612f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_137 N_A4_c_144_n A3 2.49913e-19 $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_138 A4 A3 0.0115402f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A4_c_144_n N_A3_c_197_n 0.0195612f $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_140 A4 N_A3_c_197_n 2.49913e-19 $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A4_M1016_g N_VPWR_c_345_n 0.00229957f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A4_M1016_g N_VPWR_c_347_n 0.00357877f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A4_M1017_g N_VPWR_c_347_n 0.00357877f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A4_M1016_g N_VPWR_c_342_n 0.00655123f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A4_M1017_g N_VPWR_c_342_n 0.00525237f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A4_M1016_g N_Y_c_415_n 0.0127129f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_147 N_A4_c_144_n N_Y_c_415_n 0.00580397f $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_148 A4 N_Y_c_415_n 0.0272059f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A4_M1016_g N_Y_c_416_n 0.0124577f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A4_c_144_n N_Y_c_416_n 0.00210083f $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_151 N_A4_M1017_g N_Y_c_416_n 0.00834752f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_152 A4 N_Y_c_416_n 0.0266429f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A4_c_144_n Y 6.83861e-19 $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_154 A4 Y 0.00499079f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A4_M1016_g N_A_299_297#_c_465_n 0.00926693f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A4_M1017_g N_A_299_297#_c_465_n 0.0112878f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A4_M1017_g N_A_299_297#_c_463_n 3.16391e-19 $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_158 N_A4_M1001_g N_A_27_47#_c_564_n 0.00283431f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_159 N_A4_M1001_g N_A_27_47#_c_565_n 0.0106049f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A4_c_144_n N_A_27_47#_c_565_n 0.00597682f $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_161 A4 N_A_27_47#_c_565_n 0.0266587f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A4_M1001_g N_A_27_47#_c_589_n 0.00749409f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A4_M1004_g N_A_27_47#_c_589_n 0.00655349f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A4_M1004_g N_A_27_47#_c_567_n 0.00845772f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_165 A4 N_A_27_47#_c_567_n 0.00820272f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A4_M1004_g N_A_27_47#_c_593_n 5.77985e-19 $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A4_M1001_g N_A_27_47#_c_573_n 0.00110555f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_168 N_A4_c_144_n N_A_27_47#_c_573_n 0.0021496f $X=2.25 $Y=1.025 $X2=0 $Y2=0
cc_169 N_A4_M1004_g N_A_27_47#_c_573_n 0.00110555f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_170 A4 N_A_27_47#_c_573_n 0.0265408f $X=2.01 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A4_M1001_g N_VGND_c_697_n 0.00321269f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A4_M1004_g N_VGND_c_698_n 0.00146448f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_173 N_A4_M1001_g N_VGND_c_702_n 0.00424416f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A4_M1004_g N_VGND_c_702_n 0.00424416f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A4_M1001_g N_VGND_c_712_n 0.00706214f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A4_M1004_g N_VGND_c_712_n 0.00576327f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A3_c_197_n N_A2_M1014_g 3.85179e-19 $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A3_c_195_n N_A2_c_247_n 5.45993e-19 $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_179 A3 N_A2_c_247_n 9.01325e-19 $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A3_c_197_n N_A2_c_247_n 0.0086443f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_181 A3 A2 0.0156078f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A3_M1006_g N_VPWR_c_347_n 0.00539841f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A3_M1013_g N_VPWR_c_347_n 0.00357835f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A3_M1006_g N_VPWR_c_342_n 0.00961452f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_185 N_A3_M1013_g N_VPWR_c_342_n 0.0066022f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A3_M1006_g N_A_299_297#_c_462_n 0.0124513f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A3_M1013_g N_A_299_297#_c_462_n 0.01284f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_188 A3 N_A_299_297#_c_462_n 0.0645678f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_189 N_A3_c_197_n N_A_299_297#_c_462_n 0.00629998f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A3_M1006_g N_A_549_297#_c_499_n 0.00525097f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A3_M1013_g N_A_549_297#_c_499_n 0.0110455f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_192 N_A3_M1013_g N_A_549_297#_c_498_n 0.0122179f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A3_M1006_g N_A_549_297#_c_502_n 0.00200125f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A3_M1013_g N_A_549_297#_c_502_n 7.04098e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A3_M1013_g N_A_743_297#_c_526_n 4.35828e-19 $X=3.09 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A3_c_194_n N_A_27_47#_c_589_n 5.77985e-19 $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_197 N_A3_c_194_n N_A_27_47#_c_567_n 0.00845772f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_198 A3 N_A_27_47#_c_567_n 0.00820272f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A3_c_194_n N_A_27_47#_c_593_n 0.00655349f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_200 N_A3_c_195_n N_A_27_47#_c_593_n 0.00764499f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_201 N_A3_c_195_n N_A_27_47#_c_568_n 0.0106049f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_202 A3 N_A_27_47#_c_568_n 0.0391474f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A3_c_197_n N_A_27_47#_c_568_n 0.00427365f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_204 N_A3_c_195_n N_A_27_47#_c_569_n 0.0032209f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_205 N_A3_c_194_n N_A_27_47#_c_574_n 0.00110555f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_206 N_A3_c_195_n N_A_27_47#_c_574_n 0.00110555f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_207 A3 N_A_27_47#_c_574_n 0.0265407f $X=3.39 $Y=1.105 $X2=0 $Y2=0
cc_208 N_A3_c_197_n N_A_27_47#_c_574_n 0.00221933f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A3_c_194_n N_VGND_c_698_n 0.00146448f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_210 N_A3_c_195_n N_VGND_c_699_n 0.00320466f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_211 N_A3_c_194_n N_VGND_c_704_n 0.00424416f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_212 N_A3_c_195_n N_VGND_c_704_n 0.00424416f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_213 N_A3_c_194_n N_VGND_c_712_n 0.00576327f $X=2.67 $Y=1.01 $X2=0 $Y2=0
cc_214 N_A3_c_195_n N_VGND_c_712_n 0.00706214f $X=3.09 $Y=1.01 $X2=0 $Y2=0
cc_215 N_A2_c_247_n N_A1_M1003_g 0.0150149f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_216 N_A2_M1018_g N_A1_M1000_g 0.0150149f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A2_c_247_n N_A1_c_301_n 0.0150149f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_218 N_A2_c_247_n A1 0.00159684f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_219 A2 A1 0.0169012f $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_220 N_A2_M1018_g N_VPWR_c_346_n 0.00130019f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A2_M1014_g N_VPWR_c_347_n 0.00357835f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A2_M1018_g N_VPWR_c_347_n 0.00539841f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A2_M1014_g N_VPWR_c_342_n 0.0066022f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A2_M1018_g N_VPWR_c_342_n 0.00961452f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A2_M1014_g N_A_299_297#_c_462_n 4.35828e-19 $X=4.07 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A2_M1014_g N_A_549_297#_c_498_n 0.012922f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A2_M1018_g N_A_549_297#_c_498_n 0.00202057f $X=4.49 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A2_M1014_g N_A_549_297#_c_506_n 0.0110455f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_229 N_A2_M1018_g N_A_549_297#_c_506_n 0.00525096f $X=4.49 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A2_M1014_g N_A_743_297#_c_522_n 0.0128841f $X=4.07 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A2_c_247_n N_A_743_297#_c_522_n 0.00315957f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_232 N_A2_M1018_g N_A_743_297#_c_522_n 0.0128516f $X=4.49 $Y=1.985 $X2=0 $Y2=0
cc_233 A2 N_A_743_297#_c_522_n 0.042003f $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_234 N_A2_c_247_n N_A_743_297#_c_526_n 0.00386993f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_235 A2 N_A_743_297#_c_526_n 0.0134547f $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_236 N_A2_c_245_n N_A_27_47#_c_569_n 0.00655349f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_237 N_A2_c_247_n N_A_27_47#_c_569_n 5.77985e-19 $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_238 N_A2_c_245_n N_A_27_47#_c_570_n 0.00850187f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_239 N_A2_c_247_n N_A_27_47#_c_570_n 0.0106979f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_240 A2 N_A_27_47#_c_570_n 0.0359509f $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_241 N_A2_c_245_n N_A_27_47#_c_616_n 5.77985e-19 $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_242 N_A2_c_247_n N_A_27_47#_c_616_n 0.00655349f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_243 N_A2_c_245_n N_A_27_47#_c_575_n 0.00134339f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_244 N_A2_c_247_n N_A_27_47#_c_575_n 0.00545145f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_245 A2 N_A_27_47#_c_575_n 0.0197652f $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_246 N_A2_c_247_n N_A_27_47#_c_576_n 0.00136675f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_247 A2 N_A_27_47#_c_576_n 3.84034e-19 $X=4.33 $Y=1.105 $X2=0 $Y2=0
cc_248 N_A2_c_245_n N_VGND_c_699_n 0.00208329f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_249 N_A2_c_245_n N_VGND_c_700_n 0.00268723f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_250 N_A2_c_247_n N_VGND_c_700_n 0.00146448f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_251 N_A2_c_245_n N_VGND_c_706_n 0.00424416f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_252 N_A2_c_247_n N_VGND_c_708_n 0.00424416f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_253 N_A2_c_245_n N_VGND_c_712_n 0.00706214f $X=4.07 $Y=0.99 $X2=0 $Y2=0
cc_254 N_A2_c_247_n N_VGND_c_712_n 0.00576327f $X=4.49 $Y=0.99 $X2=0 $Y2=0
cc_255 N_A1_M1000_g N_VPWR_c_346_n 0.0130033f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A1_M1008_g N_VPWR_c_346_n 0.0137667f $X=5.33 $Y=1.985 $X2=0 $Y2=0
cc_257 N_A1_M1000_g N_VPWR_c_347_n 0.0046653f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_258 N_A1_M1008_g N_VPWR_c_350_n 0.0046653f $X=5.33 $Y=1.985 $X2=0 $Y2=0
cc_259 N_A1_M1000_g N_VPWR_c_342_n 0.007919f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A1_M1008_g N_VPWR_c_342_n 0.00897951f $X=5.33 $Y=1.985 $X2=0 $Y2=0
cc_261 N_A1_M1000_g N_A_743_297#_c_523_n 0.0124912f $X=4.91 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A1_M1008_g N_A_743_297#_c_523_n 0.0128263f $X=5.33 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A1_c_301_n N_A_743_297#_c_523_n 0.00198252f $X=5.405 $Y=1.16 $X2=0
+ $Y2=0
cc_264 A1 N_A_743_297#_c_523_n 0.0474586f $X=5.71 $Y=1.105 $X2=0 $Y2=0
cc_265 N_A1_c_303_n N_A_743_297#_c_523_n 0.00107937f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_266 A1 N_A_743_297#_c_524_n 0.0203859f $X=5.71 $Y=1.105 $X2=0 $Y2=0
cc_267 N_A1_c_303_n N_A_743_297#_c_524_n 0.00573441f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_268 A1 N_A_743_297#_c_527_n 0.00555139f $X=5.71 $Y=1.105 $X2=0 $Y2=0
cc_269 N_A1_M1003_g N_A_27_47#_c_616_n 0.00655349f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A1_M1012_g N_A_27_47#_c_616_n 5.77985e-19 $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A1_M1003_g N_A_27_47#_c_571_n 0.00850187f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_272 N_A1_M1012_g N_A_27_47#_c_571_n 0.00976996f $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A1_c_301_n N_A_27_47#_c_571_n 0.00205431f $X=5.405 $Y=1.16 $X2=0 $Y2=0
cc_274 A1 N_A_27_47#_c_571_n 0.0625867f $X=5.71 $Y=1.105 $X2=0 $Y2=0
cc_275 N_A1_c_303_n N_A_27_47#_c_571_n 0.00709394f $X=5.57 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A1_M1003_g N_A_27_47#_c_572_n 5.77985e-19 $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A1_M1012_g N_A_27_47#_c_572_n 0.00655349f $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A1_M1003_g N_A_27_47#_c_576_n 0.00110056f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_279 A1 N_A_27_47#_c_576_n 0.0120882f $X=5.71 $Y=1.105 $X2=0 $Y2=0
cc_280 N_A1_M1003_g N_VGND_c_701_n 0.00146448f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A1_M1012_g N_VGND_c_701_n 0.00268723f $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A1_M1003_g N_VGND_c_708_n 0.00424416f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A1_M1012_g N_VGND_c_711_n 0.00424416f $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A1_M1003_g N_VGND_c_712_n 0.00576327f $X=4.91 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A1_M1012_g N_VGND_c_712_n 0.00682379f $X=5.33 $Y=0.56 $X2=0 $Y2=0
cc_286 N_VPWR_c_342_n N_Y_M1002_s 0.00215201f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_c_342_n N_Y_M1016_s 0.00216833f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_c_349_n N_Y_c_419_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_342_n N_Y_c_419_n 0.0122217f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_M1015_d N_Y_c_415_n 0.00296777f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_291 N_VPWR_c_345_n N_Y_c_415_n 0.0201604f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_292 N_VPWR_c_342_n N_A_299_297#_M1016_d 0.00209324f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_293 N_VPWR_c_342_n N_A_299_297#_M1017_d 0.00385313f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_342_n N_A_299_297#_M1013_d 0.00226545f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_345_n N_A_299_297#_c_460_n 0.033926f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_296 N_VPWR_c_347_n N_A_299_297#_c_465_n 0.0358391f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_342_n N_A_299_297#_c_465_n 0.0234424f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_345_n N_A_299_297#_c_461_n 0.0136295f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_299 N_VPWR_c_347_n N_A_299_297#_c_461_n 0.0172955f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_342_n N_A_299_297#_c_461_n 0.0096036f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_347_n N_A_299_297#_c_482_n 0.0114668f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_342_n N_A_299_297#_c_482_n 0.00653655f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_342_n N_A_549_297#_M1006_s 0.00215201f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_304 N_VPWR_c_342_n N_A_549_297#_M1014_s 0.00215201f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_347_n N_A_549_297#_c_498_n 0.0833579f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_342_n N_A_549_297#_c_498_n 0.0510191f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_347_n N_A_549_297#_c_502_n 0.0189579f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_342_n N_A_549_297#_c_502_n 0.0122647f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_342_n N_A_743_297#_M1014_d 0.00226545f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_310 N_VPWR_c_342_n N_A_743_297#_M1018_d 0.00562358f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_342_n N_A_743_297#_M1008_d 0.00399293f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_347_n N_A_743_297#_c_546_n 0.0113958f $X=4.955 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_342_n N_A_743_297#_c_546_n 0.00646998f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_M1000_s N_A_743_297#_c_523_n 0.00165831f $X=4.985 $Y=1.485 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_346_n N_A_743_297#_c_523_n 0.0171101f $X=5.12 $Y=2 $X2=0 $Y2=0
cc_316 N_VPWR_c_350_n N_A_743_297#_c_525_n 0.0172566f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_342_n N_A_743_297#_c_525_n 0.00955092f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_344_n N_A_27_47#_c_562_n 7.42972e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_319 N_Y_c_415_n N_A_299_297#_M1016_d 0.00296777f $X=1.875 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_320 N_Y_c_415_n N_A_299_297#_c_460_n 0.020037f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_321 N_Y_M1016_s N_A_299_297#_c_465_n 0.00312348f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_322 N_Y_c_415_n N_A_299_297#_c_465_n 0.00277146f $X=1.875 $Y=1.555 $X2=0
+ $Y2=0
cc_323 N_Y_c_416_n N_A_299_297#_c_465_n 0.015949f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_324 N_Y_c_416_n N_A_299_297#_c_463_n 0.00902116f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_325 Y N_A_27_47#_c_562_n 0.00110995f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_326 N_Y_M1009_s N_A_27_47#_c_580_n 0.00304606f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_c_430_n N_A_27_47#_c_580_n 0.0161347f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_328 N_Y_c_415_n N_A_27_47#_c_565_n 0.0080857f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_329 N_Y_c_415_n N_A_27_47#_c_566_n 0.00958572f $X=1.875 $Y=1.555 $X2=0 $Y2=0
cc_330 N_Y_c_430_n N_A_27_47#_c_566_n 0.00722085f $X=0.68 $Y=0.72 $X2=0 $Y2=0
cc_331 N_Y_M1009_s N_VGND_c_712_n 0.00216833f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_332 N_A_299_297#_c_462_n N_A_549_297#_M1006_s 0.00185611f $X=3.215 $Y=1.53
+ $X2=-0.19 $Y2=1.305
cc_333 N_A_299_297#_c_462_n N_A_549_297#_c_499_n 0.0139142f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_334 N_A_299_297#_M1013_d N_A_549_297#_c_498_n 0.00539485f $X=3.165 $Y=1.485
+ $X2=0 $Y2=0
cc_335 N_A_299_297#_c_464_n N_A_549_297#_c_498_n 0.0184944f $X=3.3 $Y=1.62 $X2=0
+ $Y2=0
cc_336 N_A_299_297#_c_462_n N_A_743_297#_c_526_n 0.0128664f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_337 N_A_299_297#_c_464_n N_A_743_297#_c_526_n 0.0329033f $X=3.3 $Y=1.62 $X2=0
+ $Y2=0
cc_338 N_A_299_297#_c_462_n N_A_27_47#_c_567_n 0.00167329f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_339 N_A_299_297#_c_463_n N_A_27_47#_c_567_n 0.00642736f $X=2.545 $Y=1.53
+ $X2=0 $Y2=0
cc_340 N_A_549_297#_c_498_n N_A_743_297#_M1014_d 0.00539485f $X=4.115 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_341 N_A_549_297#_M1014_s N_A_743_297#_c_522_n 0.00185611f $X=4.145 $Y=1.485
+ $X2=0 $Y2=0
cc_342 N_A_549_297#_c_506_n N_A_743_297#_c_522_n 0.0139142f $X=4.28 $Y=2 $X2=0
+ $Y2=0
cc_343 N_A_549_297#_c_498_n N_A_743_297#_c_526_n 0.0184944f $X=4.115 $Y=2.38
+ $X2=0 $Y2=0
cc_344 N_A_743_297#_c_526_n N_A_27_47#_c_575_n 0.00354305f $X=3.86 $Y=1.61 $X2=0
+ $Y2=0
cc_345 N_A_743_297#_c_522_n N_A_27_47#_c_576_n 0.00259965f $X=4.615 $Y=1.53
+ $X2=0 $Y2=0
cc_346 N_A_743_297#_c_527_n N_A_27_47#_c_576_n 0.00437653f $X=4.7 $Y=1.61 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_565_n N_VGND_M1001_s 0.00286661f $X=1.875 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_348 N_A_27_47#_c_567_n N_VGND_M1004_s 0.00169589f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_349 N_A_27_47#_c_568_n N_VGND_M1011_d 0.00324897f $X=3.695 $Y=0.82 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_570_n N_VGND_M1005_s 0.00169589f $X=4.535 $Y=0.82 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_571_n N_VGND_M1003_s 0.00169589f $X=5.375 $Y=0.82 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_563_n N_VGND_c_697_n 0.0168365f $X=1.14 $Y=0.465 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_564_n N_VGND_c_697_n 0.00586968f $X=1.1 $Y=0.72 $X2=0 $Y2=0
cc_354 N_A_27_47#_c_565_n N_VGND_c_697_n 0.0173651f $X=1.875 $Y=0.82 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_567_n N_VGND_c_698_n 0.0111177f $X=2.715 $Y=0.82 $X2=0 $Y2=0
cc_356 N_A_27_47#_c_568_n N_VGND_c_699_n 0.0161898f $X=3.695 $Y=0.82 $X2=0 $Y2=0
cc_357 N_A_27_47#_c_569_n N_VGND_c_699_n 0.0182479f $X=3.86 $Y=0.38 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_570_n N_VGND_c_700_n 0.0111177f $X=4.535 $Y=0.82 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_571_n N_VGND_c_701_n 0.0111177f $X=5.375 $Y=0.82 $X2=0 $Y2=0
cc_360 N_A_27_47#_c_565_n N_VGND_c_702_n 0.00193763f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_589_n N_VGND_c_702_n 0.0188551f $X=2.04 $Y=0.38 $X2=0 $Y2=0
cc_362 N_A_27_47#_c_567_n N_VGND_c_702_n 0.00193763f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_567_n N_VGND_c_704_n 0.00193763f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_593_n N_VGND_c_704_n 0.0188551f $X=2.88 $Y=0.38 $X2=0 $Y2=0
cc_365 N_A_27_47#_c_568_n N_VGND_c_704_n 0.00193763f $X=3.695 $Y=0.82 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_c_568_n N_VGND_c_706_n 0.00364836f $X=3.695 $Y=0.82 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_c_569_n N_VGND_c_706_n 0.0209479f $X=3.86 $Y=0.38 $X2=0 $Y2=0
cc_368 N_A_27_47#_c_570_n N_VGND_c_706_n 0.00193763f $X=4.535 $Y=0.82 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_570_n N_VGND_c_708_n 0.00193763f $X=4.535 $Y=0.82 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_c_616_n N_VGND_c_708_n 0.0188551f $X=4.7 $Y=0.38 $X2=0 $Y2=0
cc_371 N_A_27_47#_c_571_n N_VGND_c_708_n 0.00193763f $X=5.375 $Y=0.82 $X2=0
+ $Y2=0
cc_372 N_A_27_47#_c_561_n N_VGND_c_710_n 0.0180491f $X=0.215 $Y=0.465 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_580_n N_VGND_c_710_n 0.0362386f $X=1.015 $Y=0.36 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_563_n N_VGND_c_710_n 0.0173343f $X=1.14 $Y=0.465 $X2=0 $Y2=0
cc_375 N_A_27_47#_c_565_n N_VGND_c_710_n 0.00282598f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_571_n N_VGND_c_711_n 0.00193763f $X=5.375 $Y=0.82 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_572_n N_VGND_c_711_n 0.0209479f $X=5.54 $Y=0.38 $X2=0 $Y2=0
cc_378 N_A_27_47#_M1009_d N_VGND_c_712_n 0.00209324f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_M1019_d N_VGND_c_712_n 0.00209324f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_M1001_d N_VGND_c_712_n 0.00215201f $X=1.905 $Y=0.235 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_M1010_s N_VGND_c_712_n 0.00215201f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_M1005_d N_VGND_c_712_n 0.00225715f $X=3.715 $Y=0.235 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_M1007_d N_VGND_c_712_n 0.00215201f $X=4.565 $Y=0.235 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_M1012_d N_VGND_c_712_n 0.00225715f $X=5.405 $Y=0.235 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_561_n N_VGND_c_712_n 0.0100013f $X=0.215 $Y=0.465 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_580_n N_VGND_c_712_n 0.023553f $X=1.015 $Y=0.36 $X2=0 $Y2=0
cc_387 N_A_27_47#_c_563_n N_VGND_c_712_n 0.00961652f $X=1.14 $Y=0.465 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_565_n N_VGND_c_712_n 0.00980173f $X=1.875 $Y=0.82 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_589_n N_VGND_c_712_n 0.0122069f $X=2.04 $Y=0.38 $X2=0 $Y2=0
cc_390 N_A_27_47#_c_567_n N_VGND_c_712_n 0.00828806f $X=2.715 $Y=0.82 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_593_n N_VGND_c_712_n 0.0122069f $X=2.88 $Y=0.38 $X2=0 $Y2=0
cc_392 N_A_27_47#_c_568_n N_VGND_c_712_n 0.011185f $X=3.695 $Y=0.82 $X2=0 $Y2=0
cc_393 N_A_27_47#_c_569_n N_VGND_c_712_n 0.0124119f $X=3.86 $Y=0.38 $X2=0 $Y2=0
cc_394 N_A_27_47#_c_570_n N_VGND_c_712_n 0.00828806f $X=4.535 $Y=0.82 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_616_n N_VGND_c_712_n 0.0122069f $X=4.7 $Y=0.38 $X2=0 $Y2=0
cc_396 N_A_27_47#_c_571_n N_VGND_c_712_n 0.00828806f $X=5.375 $Y=0.82 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_572_n N_VGND_c_712_n 0.0124119f $X=5.54 $Y=0.38 $X2=0 $Y2=0

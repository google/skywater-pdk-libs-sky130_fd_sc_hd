* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
M1000 a_285_47# A VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=5.525e+11p ps=5.6e+06u
M1001 VGND a_35_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=5.005e+11p ps=2.84e+06u
M1002 VPWR B a_285_297# VPB phighvt w=1e+06u l=150000u
+  ad=5.3e+11p pd=5.06e+06u as=5.3e+11p ps=5.06e+06u
M1003 X B a_285_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_285_297# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_35_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1006 VPWR A a_117_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1007 X a_35_297# a_285_297# VPB phighvt w=1e+06u l=150000u
+  ad=3e+11p pd=2.6e+06u as=0p ps=0u
M1008 VGND A a_35_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_297# B a_35_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.6e+11p ps=2.52e+06u
.ends

* File: sky130_fd_sc_hd__clkinv_4.pex.spice
* Created: Tue Sep  1 19:01:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKINV_4%A 3 7 11 13 17 21 23 27 31 33 37 41 45 47
+ 48 49 50 51 53 54 55 56 57 58 59
r98 69 70 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r99 59 70 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=2.53 $Y=1.177
+ $X2=2.36 $Y2=1.177
r100 58 70 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=2.07 $Y=1.177
+ $X2=2.36 $Y2=1.177
r101 57 58 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=1.177
+ $X2=2.07 $Y2=1.177
r102 56 57 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=1.177
+ $X2=1.61 $Y2=1.177
r103 55 56 25.0976 $w=2.23e-07 $l=4.9e-07 $layer=LI1_cond $X=0.66 $Y=1.177
+ $X2=1.15 $Y2=1.177
r104 55 66 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r105 54 69 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=2.59 $Y=1.16 $X2=2.36
+ $Y2=1.16
r106 52 69 11.1087 $w=2.7e-07 $l=5e-08 $layer=POLY_cond $X=2.31 $Y=1.16 $X2=2.36
+ $Y2=1.16
r107 52 53 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=1.16
+ $X2=2.235 $Y2=1.16
r108 48 66 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=0.87 $Y=1.16
+ $X2=0.66 $Y2=1.16
r109 48 49 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=0.87 $Y=1.16
+ $X2=0.945 $Y2=1.16
r110 47 66 15.5522 $w=2.7e-07 $l=7e-08 $layer=POLY_cond $X=0.59 $Y=1.16 $X2=0.66
+ $Y2=1.16
r111 43 54 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.59 $Y2=1.16
r112 43 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.665 $Y=1.295
+ $X2=2.665 $Y2=1.985
r113 39 53 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.295
+ $X2=2.235 $Y2=1.16
r114 39 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.235 $Y=1.295
+ $X2=2.235 $Y2=1.985
r115 35 53 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.235 $Y=1.025
+ $X2=2.235 $Y2=1.16
r116 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.235 $Y=1.025
+ $X2=2.235 $Y2=0.445
r117 34 51 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.805 $Y2=1.16
r118 33 53 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=1.16
+ $X2=2.235 $Y2=1.16
r119 33 34 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.16 $Y=1.16
+ $X2=1.88 $Y2=1.16
r120 29 51 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.805 $Y=1.295
+ $X2=1.805 $Y2=1.16
r121 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.805 $Y=1.295
+ $X2=1.805 $Y2=1.985
r122 25 51 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.805 $Y=1.025
+ $X2=1.805 $Y2=1.16
r123 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.805 $Y=1.025
+ $X2=1.805 $Y2=0.445
r124 24 50 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.16
+ $X2=1.375 $Y2=1.16
r125 23 51 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.805 $Y2=1.16
r126 23 24 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.45 $Y2=1.16
r127 19 50 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.375 $Y2=1.16
r128 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.375 $Y=1.295
+ $X2=1.375 $Y2=1.985
r129 15 50 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.375 $Y=1.025
+ $X2=1.375 $Y2=1.16
r130 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.375 $Y=1.025
+ $X2=1.375 $Y2=0.445
r131 14 49 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=0.945 $Y2=1.16
r132 13 50 13.3889 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.3 $Y=1.16
+ $X2=1.375 $Y2=1.16
r133 13 14 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.3 $Y=1.16
+ $X2=1.02 $Y2=1.16
r134 9 49 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.945 $Y=1.295
+ $X2=0.945 $Y2=1.16
r135 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.945 $Y=1.295
+ $X2=0.945 $Y2=1.985
r136 5 49 43.38 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=1.16
r137 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=0.445
r138 1 47 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.515 $Y=1.295
+ $X2=0.59 $Y2=1.16
r139 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.515 $Y=1.295
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 34
+ 43 51 55
r52 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 46 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 43 54 5.33458 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.75 $Y=2.72
+ $X2=2.985 $Y2=2.72
r57 43 45 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.75 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 42 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r59 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 39 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.29 $Y=2.72 $X2=1.16
+ $Y2=2.72
r62 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.29 $Y=2.72 $X2=1.61
+ $Y2=2.72
r63 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 35 48 4.96256 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=2.72
+ $X2=0.215 $Y2=2.72
r66 35 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.43 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 34 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.03 $Y=2.72 $X2=1.16
+ $Y2=2.72
r68 34 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.03 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 32 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 30 41 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.89 $Y=2.72
+ $X2=1.61 $Y2=2.72
r72 30 31 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.89 $Y=2.72 $X2=2.02
+ $Y2=2.72
r73 29 45 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r74 29 31 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.15 $Y=2.72 $X2=2.02
+ $Y2=2.72
r75 25 54 2.90564 $w=3.85e-07 $l=1.04307e-07 $layer=LI1_cond $X=2.942 $Y=2.635
+ $X2=2.985 $Y2=2.72
r76 25 27 20.0555 $w=3.83e-07 $l=6.7e-07 $layer=LI1_cond $X=2.942 $Y=2.635
+ $X2=2.942 $Y2=1.965
r77 21 31 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=2.635
+ $X2=2.02 $Y2=2.72
r78 21 23 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=2.02 $Y=2.635
+ $X2=2.02 $Y2=1.965
r79 17 51 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=2.635
+ $X2=1.16 $Y2=2.72
r80 17 19 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.16 $Y=2.635
+ $X2=1.16 $Y2=1.965
r81 13 48 2.93137 $w=3.45e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.215 $Y2=2.72
r82 13 15 22.3808 $w=3.43e-07 $l=6.7e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=1.965
r83 4 27 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.485 $X2=2.88 $Y2=1.965
r84 3 23 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.485 $X2=2.02 $Y2=1.965
r85 2 19 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=1.485 $X2=1.16 $Y2=1.965
r86 1 15 300 $w=1.7e-07 $l=5.56417e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.3 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_4%Y 1 2 3 4 5 17 18 19 20 21 24 26 30 32 36
+ 38 42 44 48 50 52 53 54 55 56 57 58 59 65 66
r107 59 66 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=1.545
+ $X2=2.985 $Y2=1.46
r108 59 66 0.307318 $w=2.98e-07 $l=8e-09 $layer=LI1_cond $X=2.985 $Y=1.452
+ $X2=2.985 $Y2=1.46
r109 58 59 10.0647 $w=2.98e-07 $l=2.62e-07 $layer=LI1_cond $X=2.985 $Y=1.19
+ $X2=2.985 $Y2=1.452
r110 57 65 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.81
+ $X2=2.985 $Y2=0.895
r111 57 58 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=2.985 $Y=0.915
+ $X2=2.985 $Y2=1.19
r112 57 65 0.768295 $w=2.98e-07 $l=2e-08 $layer=LI1_cond $X=2.985 $Y=0.915
+ $X2=2.985 $Y2=0.895
r113 51 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.58 $Y=1.545
+ $X2=2.45 $Y2=1.545
r114 50 59 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.835 $Y=1.545
+ $X2=2.985 $Y2=1.545
r115 50 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.835 $Y=1.545
+ $X2=2.58 $Y2=1.545
r116 46 56 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=1.63
+ $X2=2.45 $Y2=1.545
r117 46 48 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=2.45 $Y=1.63 $X2=2.45
+ $Y2=1.83
r118 45 55 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.145 $Y=0.81
+ $X2=2.017 $Y2=0.81
r119 44 57 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.835 $Y=0.81
+ $X2=2.985 $Y2=0.81
r120 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.835 $Y=0.81
+ $X2=2.145 $Y2=0.81
r121 40 55 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.017 $Y=0.725
+ $X2=2.017 $Y2=0.81
r122 40 42 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.017 $Y=0.725
+ $X2=2.017 $Y2=0.445
r123 39 54 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.72 $Y=1.545
+ $X2=1.592 $Y2=1.545
r124 38 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.32 $Y=1.545
+ $X2=2.45 $Y2=1.545
r125 38 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.32 $Y=1.545
+ $X2=1.72 $Y2=1.545
r126 34 54 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.592 $Y=1.63
+ $X2=1.592 $Y2=1.545
r127 34 36 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=1.592 $Y=1.63
+ $X2=1.592 $Y2=1.83
r128 33 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.29 $Y=0.81
+ $X2=1.16 $Y2=0.81
r129 32 55 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.89 $Y=0.81
+ $X2=2.017 $Y2=0.81
r130 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.89 $Y=0.81 $X2=1.29
+ $Y2=0.81
r131 28 53 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.725
+ $X2=1.16 $Y2=0.81
r132 28 30 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.16 $Y=0.725
+ $X2=1.16 $Y2=0.445
r133 27 52 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.86 $Y=1.545
+ $X2=0.732 $Y2=1.545
r134 26 54 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.465 $Y=1.545
+ $X2=1.592 $Y2=1.545
r135 26 27 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.465 $Y=1.545
+ $X2=0.86 $Y2=1.545
r136 22 52 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.732 $Y=1.63
+ $X2=0.732 $Y2=1.545
r137 22 24 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=0.732 $Y=1.63
+ $X2=0.732 $Y2=1.83
r138 20 52 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.605 $Y=1.545
+ $X2=0.732 $Y2=1.545
r139 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.605 $Y=1.545
+ $X2=0.275 $Y2=1.545
r140 18 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.03 $Y=0.81
+ $X2=1.16 $Y2=0.81
r141 18 19 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.03 $Y=0.81
+ $X2=0.275 $Y2=0.81
r142 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=1.46
+ $X2=0.275 $Y2=1.545
r143 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.275 $Y2=0.81
r144 16 17 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.19 $Y2=1.46
r145 5 48 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=2.31
+ $Y=1.485 $X2=2.45 $Y2=1.83
r146 4 36 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.485 $X2=1.59 $Y2=1.83
r147 3 24 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.73 $Y2=1.83
r148 2 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.02 $Y2=0.445
r149 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.16 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKINV_4%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r45 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r47 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r49 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r50 39 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.465
+ $Y2=0
r51 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.99
+ $Y2=0
r52 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r53 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r54 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r55 35 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=1.59
+ $Y2=0
r56 35 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.72 $Y=0 $X2=2.07
+ $Y2=0
r57 34 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.465
+ $Y2=0
r58 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.07
+ $Y2=0
r59 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r60 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r61 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 30 45 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=0.712
+ $Y2=0
r63 30 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0 $X2=1.15
+ $Y2=0
r64 29 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.59
+ $Y2=0
r65 29 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.15
+ $Y2=0
r66 24 45 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.712
+ $Y2=0
r67 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.23
+ $Y2=0
r68 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 18 51 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0
r71 18 20 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0.085
+ $X2=2.465 $Y2=0.39
r72 14 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r73 14 16 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.39
r74 10 45 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r75 10 12 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.39
r76 3 20 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.235 $X2=2.45 $Y2=0.39
r77 2 16 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.59 $Y2=0.39
r78 1 12 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=0.54
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__nand4b_4.pxi.spice
* Created: Tue Sep  1 19:17:10 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4B_4%A_N N_A_N_c_145_n N_A_N_M1030_g N_A_N_M1024_g A_N
+ N_A_N_c_147_n PM_SKY130_FD_SC_HD__NAND4B_4%A_N
x_PM_SKY130_FD_SC_HD__NAND4B_4%A_27_47# N_A_27_47#_M1030_s N_A_27_47#_M1024_s
+ N_A_27_47#_M1005_g N_A_27_47#_M1001_g N_A_27_47#_M1008_g N_A_27_47#_M1020_g
+ N_A_27_47#_M1012_g N_A_27_47#_M1025_g N_A_27_47#_M1019_g N_A_27_47#_M1027_g
+ N_A_27_47#_c_183_n N_A_27_47#_c_196_n N_A_27_47#_c_197_n N_A_27_47#_c_184_n
+ N_A_27_47#_c_185_n N_A_27_47#_c_198_n N_A_27_47#_c_186_n N_A_27_47#_c_187_n
+ N_A_27_47#_c_188_n N_A_27_47#_c_189_n N_A_27_47#_c_190_n N_A_27_47#_c_191_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND4B_4%B N_B_M1010_g N_B_M1014_g N_B_M1013_g N_B_M1016_g
+ N_B_M1017_g N_B_M1021_g N_B_M1018_g N_B_M1028_g B B B B N_B_c_312_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%B
x_PM_SKY130_FD_SC_HD__NAND4B_4%C N_C_M1000_g N_C_M1002_g N_C_M1003_g N_C_M1022_g
+ N_C_M1006_g N_C_M1029_g N_C_M1033_g N_C_M1031_g C C C C N_C_c_398_n
+ N_C_c_399_n N_C_c_400_n PM_SKY130_FD_SC_HD__NAND4B_4%C
x_PM_SKY130_FD_SC_HD__NAND4B_4%D N_D_M1004_g N_D_M1015_g N_D_M1007_g N_D_M1023_g
+ N_D_M1009_g N_D_M1026_g N_D_M1011_g N_D_M1032_g D D D D N_D_c_480_n
+ N_D_c_481_n PM_SKY130_FD_SC_HD__NAND4B_4%D
x_PM_SKY130_FD_SC_HD__NAND4B_4%VPWR N_VPWR_M1024_d N_VPWR_M1001_s N_VPWR_M1020_s
+ N_VPWR_M1027_s N_VPWR_M1016_s N_VPWR_M1028_s N_VPWR_M1022_d N_VPWR_M1031_d
+ N_VPWR_M1023_d N_VPWR_M1032_d N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n
+ N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n
+ N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n
+ N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n
+ N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n
+ VPWR N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n
+ N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_562_n PM_SKY130_FD_SC_HD__NAND4B_4%VPWR
x_PM_SKY130_FD_SC_HD__NAND4B_4%Y N_Y_M1005_s N_Y_M1012_s N_Y_M1001_d N_Y_M1025_d
+ N_Y_M1014_d N_Y_M1021_d N_Y_M1002_s N_Y_M1029_s N_Y_M1015_s N_Y_M1026_s
+ N_Y_c_697_n N_Y_c_699_n N_Y_c_725_n N_Y_c_700_n N_Y_c_732_n N_Y_c_735_n
+ N_Y_c_701_n N_Y_c_754_n N_Y_c_702_n N_Y_c_779_n N_Y_c_703_n N_Y_c_786_n
+ N_Y_c_704_n N_Y_c_791_n N_Y_c_705_n N_Y_c_706_n N_Y_c_813_n N_Y_c_707_n
+ N_Y_c_708_n N_Y_c_709_n N_Y_c_710_n N_Y_c_711_n N_Y_c_712_n Y Y Y N_Y_c_745_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%Y
x_PM_SKY130_FD_SC_HD__NAND4B_4%VGND N_VGND_M1030_d N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n
+ VGND N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n N_VGND_c_879_n
+ N_VGND_c_880_n N_VGND_c_881_n PM_SKY130_FD_SC_HD__NAND4B_4%VGND
x_PM_SKY130_FD_SC_HD__NAND4B_4%A_215_47# N_A_215_47#_M1005_d N_A_215_47#_M1008_d
+ N_A_215_47#_M1019_d N_A_215_47#_M1013_s N_A_215_47#_M1018_s
+ N_A_215_47#_c_972_n N_A_215_47#_c_973_n N_A_215_47#_c_974_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%A_215_47#
x_PM_SKY130_FD_SC_HD__NAND4B_4%A_633_47# N_A_633_47#_M1010_d N_A_633_47#_M1017_d
+ N_A_633_47#_M1000_s N_A_633_47#_M1006_s N_A_633_47#_c_1016_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%A_633_47#
x_PM_SKY130_FD_SC_HD__NAND4B_4%A_991_47# N_A_991_47#_M1000_d N_A_991_47#_M1003_d
+ N_A_991_47#_M1033_d N_A_991_47#_M1007_d N_A_991_47#_M1011_d
+ N_A_991_47#_c_1050_n N_A_991_47#_c_1060_n N_A_991_47#_c_1061_n
+ N_A_991_47#_c_1051_n N_A_991_47#_c_1052_n N_A_991_47#_c_1068_n
+ N_A_991_47#_c_1053_n N_A_991_47#_c_1054_n N_A_991_47#_c_1055_n
+ PM_SKY130_FD_SC_HD__NAND4B_4%A_991_47#
cc_1 VNB N_A_N_c_145_n 0.0248249f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB A_N 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_147_n 0.0394785f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_A_27_47#_M1005_g 0.0215979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_M1001_g 5.56194e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_6 VNB N_A_27_47#_M1008_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1020_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1012_g 0.0172529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1025_g 4.47552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1019_g 0.0171875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1027_g 4.28089e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_183_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_184_n 0.00234584f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_185_n 0.00924007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_186_n 0.0041304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_187_n 7.89459e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_188_n 0.00934767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_189_n 0.00250524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_190_n 0.0330574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_191_n 0.0585093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B_M1010_g 0.0176939f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_B_M1014_g 4.64995e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B_M1013_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_24 VNB N_B_M1016_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_B_M1017_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_M1021_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_B_M1018_g 0.023095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB B 0.00341317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_B_c_312_n 0.0748536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_C_M1000_g 0.0237399f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_31 VNB N_C_M1002_g 5.64907e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_C_M1003_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_33 VNB N_C_M1022_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_C_M1006_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_C_M1029_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_C_M1033_g 0.0176998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_C_M1031_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_C_c_398_n 0.0331062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_C_c_399_n 0.00184776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_C_c_400_n 0.0582445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_D_M1004_g 0.017551f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_42 VNB N_D_M1015_g 4.65797e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_D_M1007_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_44 VNB N_D_M1023_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_D_M1009_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_D_M1026_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_D_M1011_g 0.0230765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB D 0.00946594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_D_c_480_n 0.0589025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_D_c_481_n 0.029112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VPWR_c_562_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_697_n 0.00505016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB Y 0.00123574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_871_n 0.00858498f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_55 VNB N_VGND_c_872_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_873_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_874_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_875_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_876_n 0.0171909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_877_n 0.142193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_878_n 0.0184638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_879_n 0.42228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_880_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_881_n 0.00323567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_215_47#_c_972_n 0.00217944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_215_47#_c_973_n 0.00643123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_215_47#_c_974_n 0.00252967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_633_47#_c_1016_n 0.0256487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_991_47#_c_1050_n 0.00245677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_991_47#_c_1051_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_991_47#_c_1052_n 0.00353671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_991_47#_c_1053_n 0.0112299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_991_47#_c_1054_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_991_47#_c_1055_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VPB N_A_N_M1024_g 0.0293659f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_76 VPB N_A_N_c_147_n 0.00860623f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_77 VPB N_A_27_47#_M1001_g 0.0241952f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_78 VPB N_A_27_47#_M1020_g 0.0191612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_M1025_g 0.019143f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_M1027_g 0.0188875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_196_n 0.00769697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_197_n 0.0314532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_198_n 0.00130953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_187_n 0.00459877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_B_M1014_g 0.0194556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_B_M1016_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_B_M1021_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_B_M1028_g 0.0266409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_B_c_312_n 0.00387272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_C_M1002_g 0.026721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_C_M1022_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_C_M1029_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_C_M1031_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_D_M1015_g 0.0194869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_D_M1023_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_D_M1026_g 0.0191843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_D_M1032_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_D_c_481_n 0.00976317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_563_n 0.0100313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_564_n 0.00466099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_565_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_566_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_567_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_568_n 0.00645473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_569_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_570_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_571_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_572_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_573_n 0.0112234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_574_n 0.0457449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_575_n 0.00644865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_576_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_577_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_578_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_579_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_580_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_581_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_582_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_583_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_584_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_585_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_586_n 0.0178188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_587_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_588_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_589_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_590_n 0.0132394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_591_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_562_n 0.0456476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Y_c_699_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Y_c_700_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_Y_c_701_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_Y_c_702_n 0.00714557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_Y_c_703_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_Y_c_704_n 0.0051021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_Y_c_705_n 0.00219943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_Y_c_706_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_Y_c_707_n 0.00714987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_Y_c_708_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_Y_c_709_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_Y_c_710_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Y_c_711_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_Y_c_712_n 0.00223815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB Y 0.00133154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB Y 6.61229e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 N_A_N_c_145_n N_A_27_47#_c_183_n 0.00749409f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_N_M1024_g N_A_27_47#_c_196_n 9.46316e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_147 A_N N_A_27_47#_c_196_n 0.0184258f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A_N_c_147_n N_A_27_47#_c_196_n 0.00604186f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_N_M1024_g N_A_27_47#_c_197_n 0.0106625f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_N_c_145_n N_A_27_47#_c_184_n 0.0111694f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_151 A_N N_A_27_47#_c_184_n 9.95686e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A_N_c_145_n N_A_27_47#_c_185_n 0.00126954f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_153 A_N N_A_27_47#_c_185_n 0.0254514f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_N_c_147_n N_A_27_47#_c_185_n 0.00695726f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_N_M1024_g N_A_27_47#_c_198_n 0.0134143f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_156 A_N N_A_27_47#_c_198_n 8.10212e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A_N_c_145_n N_A_27_47#_c_186_n 0.00608685f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_N_c_147_n N_A_27_47#_c_187_n 0.00836542f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_159 A_N N_A_27_47#_c_189_n 0.0167772f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_160 N_A_N_c_147_n N_A_27_47#_c_189_n 0.00240443f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_N_c_147_n N_A_27_47#_c_190_n 0.0056585f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_N_M1024_g N_VPWR_c_563_n 0.0048073f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_N_M1024_g N_VPWR_c_564_n 0.00320962f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_N_M1024_g N_VPWR_c_586_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_N_M1024_g N_VPWR_c_562_n 0.0117818f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_N_c_145_n N_VGND_c_871_n 0.0044954f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_N_c_145_n N_VGND_c_876_n 0.00424416f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_N_c_145_n N_VGND_c_879_n 0.00801635f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_N_c_145_n N_A_215_47#_c_973_n 0.00354381f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1019_g N_B_M1010_g 0.0269031f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_27_47#_M1027_g N_B_M1014_g 0.0301081f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_191_n B 0.0016612f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_191_n N_B_c_312_n 0.0187797f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_198_n N_VPWR_M1024_d 0.00486366f $X=0.61 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_27_47#_c_187_n N_VPWR_M1024_d 2.96637e-19 $X=0.707 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_27_47#_M1001_g N_VPWR_c_563_n 0.0033532f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_197_n N_VPWR_c_564_n 0.00532029f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_198_n N_VPWR_c_564_n 0.0135165f $X=0.61 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_188_n N_VPWR_c_564_n 0.0188025f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_190_n N_VPWR_c_564_n 0.00621923f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1020_g N_VPWR_c_565_n 0.00146448f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1025_g N_VPWR_c_565_n 0.00146448f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_M1027_g N_VPWR_c_566_n 0.00146448f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_198_n N_VPWR_c_575_n 0.0180607f $X=0.61 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_188_n N_VPWR_c_575_n 0.00706024f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_M1001_g N_VPWR_c_576_n 0.00541359f $X=1.41 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_M1020_g N_VPWR_c_576_n 0.00541359f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1025_g N_VPWR_c_578_n 0.00541359f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_M1027_g N_VPWR_c_578_n 0.00541359f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_197_n N_VPWR_c_586_n 0.0213966f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_191 N_A_27_47#_M1024_s N_VPWR_c_562_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1001_g N_VPWR_c_562_n 0.0108276f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1020_g N_VPWR_c_562_n 0.00950154f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1025_g N_VPWR_c_562_n 0.00950154f $X=2.25 $Y=1.985 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_M1027_g N_VPWR_c_562_n 0.00952874f $X=2.67 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_197_n N_VPWR_c_562_n 0.0126193f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_197 N_A_27_47#_M1005_g N_Y_c_697_n 0.00398755f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1008_g N_Y_c_697_n 0.0112239f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1012_g N_Y_c_697_n 0.0125587f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_188_n N_Y_c_697_n 0.0555084f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_191_n N_Y_c_697_n 0.00415773f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1001_g N_Y_c_699_n 0.00388437f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_27_47#_M1020_g N_Y_c_699_n 0.00149073f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_187_n N_Y_c_699_n 0.00141121f $X=0.707 $Y=1.495 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_188_n N_Y_c_699_n 0.026643f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_191_n N_Y_c_699_n 0.00206439f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1001_g N_Y_c_725_n 0.00902485f $X=1.41 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1020_g N_Y_c_725_n 0.00975139f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_209 N_A_27_47#_M1025_g N_Y_c_725_n 6.1949e-19 $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1020_g N_Y_c_700_n 0.0120357f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_27_47#_M1025_g N_Y_c_700_n 0.0130373f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_188_n N_Y_c_700_n 0.0304181f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_191_n N_Y_c_700_n 0.0019951f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_27_47#_M1020_g N_Y_c_732_n 6.1949e-19 $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1025_g N_Y_c_732_n 0.00975139f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_27_47#_M1027_g N_Y_c_732_n 0.00975139f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1027_g N_Y_c_735_n 6.1949e-19 $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_218 N_A_27_47#_M1027_g N_Y_c_707_n 0.0140789f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A_27_47#_M1012_g Y 0.00309532f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A_27_47#_M1025_g Y 0.00387565f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1019_g Y 0.00330868f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_27_47#_M1027_g Y 0.00414987f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_188_n Y 0.0155586f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_191_n Y 0.0199186f $X=2.67 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1025_g Y 0.00180793f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A_27_47#_M1027_g Y 0.00209341f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1019_g N_Y_c_745_n 0.00573509f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_184_n N_VGND_M1030_d 0.00464211f $X=0.61 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_229 N_A_27_47#_M1005_g N_VGND_c_871_n 0.00229957f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_184_n N_VGND_c_871_n 0.015871f $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_188_n N_VGND_c_871_n 0.00148402f $X=2.04 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_183_n N_VGND_c_876_n 0.0213324f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_184_n N_VGND_c_876_n 0.00193763f $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_234 N_A_27_47#_M1005_g N_VGND_c_877_n 0.00357877f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1008_g N_VGND_c_877_n 0.00357877f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_236 N_A_27_47#_M1012_g N_VGND_c_877_n 0.00357877f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A_27_47#_M1019_g N_VGND_c_877_n 0.00357877f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A_27_47#_M1030_s N_VGND_c_879_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1005_g N_VGND_c_879_n 0.00655123f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_240 N_A_27_47#_M1008_g N_VGND_c_879_n 0.00522516f $X=1.83 $Y=0.56 $X2=0 $Y2=0
cc_241 N_A_27_47#_M1012_g N_VGND_c_879_n 0.00522516f $X=2.25 $Y=0.56 $X2=0 $Y2=0
cc_242 N_A_27_47#_M1019_g N_VGND_c_879_n 0.00525237f $X=2.67 $Y=0.56 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_183_n N_VGND_c_879_n 0.0126042f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_184_n N_VGND_c_879_n 0.00474294f $X=0.61 $Y=0.82 $X2=0 $Y2=0
cc_245 N_A_27_47#_M1005_g N_A_215_47#_c_973_n 4.61765e-19 $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_183_n N_A_215_47#_c_973_n 0.0055786f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_184_n N_A_215_47#_c_973_n 0.0116908f $X=0.61 $Y=0.82 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_188_n N_A_215_47#_c_973_n 0.0201437f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_190_n N_A_215_47#_c_973_n 0.00588114f $X=1.335 $Y=1.16 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1005_g N_A_215_47#_c_974_n 0.0103313f $X=1.41 $Y=0.56 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1008_g N_A_215_47#_c_974_n 0.00866705f $X=1.83 $Y=0.56 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_M1012_g N_A_215_47#_c_974_n 0.00866705f $X=2.25 $Y=0.56 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_M1019_g N_A_215_47#_c_974_n 0.0119423f $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_188_n N_A_215_47#_c_974_n 0.00348394f $X=2.04 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_191_n N_A_215_47#_c_974_n 2.87379e-19 $X=2.67 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1019_g N_A_633_47#_c_1016_n 7.78229e-19 $X=2.67 $Y=0.56 $X2=0
+ $Y2=0
cc_257 N_B_c_312_n N_C_M1000_g 2.44664e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B_c_312_n N_C_M1002_g 2.44664e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_259 B N_C_c_398_n 2.32928e-19 $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_260 N_B_c_312_n N_C_c_398_n 0.0171123f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_261 B N_C_c_399_n 0.0156078f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_262 N_B_c_312_n N_C_c_399_n 7.96599e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B_M1014_g N_VPWR_c_566_n 0.00146448f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_264 N_B_M1016_g N_VPWR_c_567_n 0.00146448f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_265 N_B_M1021_g N_VPWR_c_567_n 0.00146448f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_266 N_B_M1028_g N_VPWR_c_568_n 0.0158595f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_267 N_B_M1014_g N_VPWR_c_580_n 0.00541359f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_268 N_B_M1016_g N_VPWR_c_580_n 0.00541359f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_269 N_B_M1021_g N_VPWR_c_587_n 0.00541359f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_270 N_B_M1028_g N_VPWR_c_587_n 0.00541359f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_271 N_B_M1014_g N_VPWR_c_562_n 0.00952874f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_272 N_B_M1016_g N_VPWR_c_562_n 0.00950154f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_273 N_B_M1021_g N_VPWR_c_562_n 0.00950154f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_274 N_B_M1028_g N_VPWR_c_562_n 0.0109543f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_275 N_B_M1014_g N_Y_c_732_n 6.1949e-19 $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_276 N_B_M1014_g N_Y_c_735_n 0.00975139f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_277 N_B_M1016_g N_Y_c_735_n 0.00975139f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_278 N_B_M1021_g N_Y_c_735_n 6.1949e-19 $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_279 N_B_M1016_g N_Y_c_701_n 0.0120357f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_280 N_B_M1021_g N_Y_c_701_n 0.0120357f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_281 B N_Y_c_701_n 0.0366837f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_282 N_B_c_312_n N_Y_c_701_n 0.0019951f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_283 N_B_M1016_g N_Y_c_754_n 6.1949e-19 $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_284 N_B_M1021_g N_Y_c_754_n 0.00975139f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_285 N_B_M1028_g N_Y_c_754_n 0.0145598f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_286 N_B_M1028_g N_Y_c_702_n 0.0147646f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_287 B N_Y_c_702_n 0.0205565f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_288 N_B_c_312_n N_Y_c_702_n 0.00375551f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B_M1014_g N_Y_c_707_n 0.0119784f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_290 B N_Y_c_707_n 0.0147425f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_291 N_B_c_312_n N_Y_c_707_n 0.00133007f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_292 N_B_M1014_g N_Y_c_708_n 0.00149073f $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_293 N_B_M1016_g N_Y_c_708_n 0.00149073f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_294 B N_Y_c_708_n 0.026643f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_295 N_B_c_312_n N_Y_c_708_n 0.00206439f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_296 N_B_M1021_g N_Y_c_709_n 0.00149073f $X=3.93 $Y=1.985 $X2=0 $Y2=0
cc_297 N_B_M1028_g N_Y_c_709_n 0.00149073f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_298 B N_Y_c_709_n 0.026643f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_299 N_B_c_312_n N_Y_c_709_n 0.00206439f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_300 N_B_M1010_g Y 6.04393e-19 $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_301 N_B_M1014_g Y 7.57491e-19 $X=3.09 $Y=1.985 $X2=0 $Y2=0
cc_302 B Y 0.0110559f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_303 N_B_c_312_n Y 6.42444e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_304 N_B_M1010_g N_Y_c_745_n 8.12273e-19 $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_305 N_B_M1010_g N_VGND_c_877_n 0.00357877f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_306 N_B_M1013_g N_VGND_c_877_n 0.00357877f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_307 N_B_M1017_g N_VGND_c_877_n 0.00357877f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_308 N_B_M1018_g N_VGND_c_877_n 0.00357877f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_309 N_B_M1010_g N_VGND_c_879_n 0.00525237f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_310 N_B_M1013_g N_VGND_c_879_n 0.00522516f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_311 N_B_M1017_g N_VGND_c_879_n 0.00522516f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_312 N_B_M1018_g N_VGND_c_879_n 0.00655123f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_313 N_B_M1010_g N_A_215_47#_c_974_n 0.0103313f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_314 N_B_M1013_g N_A_215_47#_c_974_n 0.00866705f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_315 N_B_M1017_g N_A_215_47#_c_974_n 0.00866705f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_316 N_B_M1018_g N_A_215_47#_c_974_n 0.00866705f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_317 B N_A_215_47#_c_974_n 0.00441672f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_318 N_B_c_312_n N_A_215_47#_c_974_n 7.82777e-19 $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_319 N_B_M1010_g N_A_633_47#_c_1016_n 0.00563386f $X=3.09 $Y=0.56 $X2=0 $Y2=0
cc_320 N_B_M1013_g N_A_633_47#_c_1016_n 0.0112239f $X=3.51 $Y=0.56 $X2=0 $Y2=0
cc_321 N_B_M1017_g N_A_633_47#_c_1016_n 0.0112239f $X=3.93 $Y=0.56 $X2=0 $Y2=0
cc_322 N_B_M1018_g N_A_633_47#_c_1016_n 0.0145787f $X=4.35 $Y=0.56 $X2=0 $Y2=0
cc_323 B N_A_633_47#_c_1016_n 0.107394f $X=4.31 $Y=1.105 $X2=0 $Y2=0
cc_324 N_B_c_312_n N_A_633_47#_c_1016_n 0.0101499f $X=4.35 $Y=1.16 $X2=0 $Y2=0
cc_325 N_C_M1033_g N_D_M1004_g 0.0200474f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_326 N_C_M1031_g N_D_M1015_g 0.0200474f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_327 N_C_c_399_n D 0.0068506f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_328 N_C_c_400_n D 7.60646e-19 $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_329 N_C_c_399_n N_D_c_480_n 7.68131e-19 $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_330 N_C_c_400_n N_D_c_480_n 0.0200474f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_331 N_C_M1002_g N_VPWR_c_568_n 0.0158595f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_332 N_C_M1022_g N_VPWR_c_569_n 0.00146448f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_333 N_C_M1029_g N_VPWR_c_569_n 0.00146448f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_334 N_C_M1031_g N_VPWR_c_570_n 0.00146448f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_335 N_C_M1002_g N_VPWR_c_582_n 0.00541359f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_336 N_C_M1022_g N_VPWR_c_582_n 0.00541359f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_337 N_C_M1029_g N_VPWR_c_584_n 0.00541359f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_338 N_C_M1031_g N_VPWR_c_584_n 0.00541359f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_339 N_C_M1002_g N_VPWR_c_562_n 0.0109543f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_340 N_C_M1022_g N_VPWR_c_562_n 0.00950154f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_341 N_C_M1029_g N_VPWR_c_562_n 0.00950154f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_342 N_C_M1031_g N_VPWR_c_562_n 0.00952874f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_343 N_C_M1002_g N_Y_c_702_n 0.0147646f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_344 N_C_c_398_n N_Y_c_702_n 0.00873655f $X=5.215 $Y=1.16 $X2=0 $Y2=0
cc_345 N_C_c_399_n N_Y_c_702_n 0.0398476f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_346 N_C_M1002_g N_Y_c_779_n 0.0145598f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_347 N_C_M1022_g N_Y_c_779_n 0.00975139f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_348 N_C_M1029_g N_Y_c_779_n 6.1949e-19 $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_349 N_C_M1022_g N_Y_c_703_n 0.0120357f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_350 N_C_M1029_g N_Y_c_703_n 0.0120357f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_351 N_C_c_399_n N_Y_c_703_n 0.0366837f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_352 N_C_c_400_n N_Y_c_703_n 0.0019951f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_353 N_C_M1022_g N_Y_c_786_n 6.1949e-19 $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_354 N_C_M1029_g N_Y_c_786_n 0.00975139f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_355 N_C_M1031_g N_Y_c_786_n 0.00975139f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_356 N_C_M1031_g N_Y_c_704_n 0.0155716f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_357 N_C_c_399_n N_Y_c_704_n 3.14784e-19 $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_358 N_C_M1031_g N_Y_c_791_n 6.1949e-19 $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_359 N_C_M1002_g N_Y_c_710_n 0.00149073f $X=5.29 $Y=1.985 $X2=0 $Y2=0
cc_360 N_C_M1022_g N_Y_c_710_n 0.00149073f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_361 N_C_c_399_n N_Y_c_710_n 0.026643f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_362 N_C_c_400_n N_Y_c_710_n 0.00206439f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_363 N_C_M1029_g N_Y_c_711_n 0.00149073f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_364 N_C_M1031_g N_Y_c_711_n 0.00149073f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_365 N_C_c_399_n N_Y_c_711_n 0.026643f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_366 N_C_c_400_n N_Y_c_711_n 0.00206439f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_367 N_C_M1000_g N_VGND_c_877_n 0.00357877f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_368 N_C_M1003_g N_VGND_c_877_n 0.00357877f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_369 N_C_M1006_g N_VGND_c_877_n 0.00357877f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_370 N_C_M1033_g N_VGND_c_877_n 0.00357877f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_371 N_C_M1000_g N_VGND_c_879_n 0.00655123f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_372 N_C_M1003_g N_VGND_c_879_n 0.00522516f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_373 N_C_M1006_g N_VGND_c_879_n 0.00522516f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_374 N_C_M1033_g N_VGND_c_879_n 0.00525237f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_375 N_C_M1000_g N_A_633_47#_c_1016_n 0.0145787f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_376 N_C_M1003_g N_A_633_47#_c_1016_n 0.0112239f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_377 N_C_M1006_g N_A_633_47#_c_1016_n 0.0112239f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_378 N_C_M1033_g N_A_633_47#_c_1016_n 0.00383287f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_379 N_C_c_398_n N_A_633_47#_c_1016_n 0.00910351f $X=5.215 $Y=1.16 $X2=0 $Y2=0
cc_380 N_C_c_399_n N_A_633_47#_c_1016_n 0.127005f $X=6.345 $Y=1.16 $X2=0 $Y2=0
cc_381 N_C_c_400_n N_A_633_47#_c_1016_n 0.0062366f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_382 N_C_M1000_g N_A_991_47#_c_1050_n 0.00866705f $X=5.29 $Y=0.56 $X2=0 $Y2=0
cc_383 N_C_M1003_g N_A_991_47#_c_1050_n 0.00866705f $X=5.71 $Y=0.56 $X2=0 $Y2=0
cc_384 N_C_M1006_g N_A_991_47#_c_1050_n 0.00866705f $X=6.13 $Y=0.56 $X2=0 $Y2=0
cc_385 N_C_M1033_g N_A_991_47#_c_1050_n 0.0123292f $X=6.55 $Y=0.56 $X2=0 $Y2=0
cc_386 N_D_M1015_g N_VPWR_c_570_n 0.00146448f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_387 N_D_M1015_g N_VPWR_c_571_n 0.00541359f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_388 N_D_M1023_g N_VPWR_c_571_n 0.00541359f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_389 N_D_M1023_g N_VPWR_c_572_n 0.00146448f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_390 N_D_M1026_g N_VPWR_c_572_n 0.00146448f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_391 N_D_M1032_g N_VPWR_c_574_n 0.0041053f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_392 D N_VPWR_c_574_n 0.0206302f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_393 N_D_c_481_n N_VPWR_c_574_n 0.00595724f $X=8.47 $Y=1.16 $X2=0 $Y2=0
cc_394 N_D_M1026_g N_VPWR_c_588_n 0.00541359f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_395 N_D_M1032_g N_VPWR_c_588_n 0.00541359f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_396 N_D_M1015_g N_VPWR_c_562_n 0.00952874f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_397 N_D_M1023_g N_VPWR_c_562_n 0.00950154f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_398 N_D_M1026_g N_VPWR_c_562_n 0.00950154f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_399 N_D_M1032_g N_VPWR_c_562_n 0.010492f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_400 N_D_M1015_g N_Y_c_786_n 6.1949e-19 $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_401 N_D_M1015_g N_Y_c_704_n 0.013439f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_402 N_D_M1015_g N_Y_c_791_n 0.00975139f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_403 N_D_M1023_g N_Y_c_791_n 0.00975139f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_404 N_D_M1026_g N_Y_c_791_n 6.1949e-19 $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_405 N_D_M1023_g N_Y_c_705_n 0.0120357f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_406 N_D_M1026_g N_Y_c_705_n 0.0120357f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_407 D N_Y_c_705_n 0.0366837f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_408 N_D_c_480_n N_Y_c_705_n 0.0019951f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_409 N_D_M1026_g N_Y_c_706_n 0.00149073f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_410 N_D_M1032_g N_Y_c_706_n 0.00331821f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_411 D N_Y_c_706_n 0.026643f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_412 N_D_c_480_n N_Y_c_706_n 0.00206439f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_413 N_D_M1023_g N_Y_c_813_n 6.1949e-19 $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_414 N_D_M1026_g N_Y_c_813_n 0.00975139f $X=7.81 $Y=1.985 $X2=0 $Y2=0
cc_415 N_D_M1032_g N_Y_c_813_n 0.00902485f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_416 N_D_M1015_g N_Y_c_712_n 0.00149073f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_417 N_D_M1023_g N_Y_c_712_n 0.00149073f $X=7.39 $Y=1.985 $X2=0 $Y2=0
cc_418 D N_Y_c_712_n 0.026643f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_419 N_D_c_480_n N_Y_c_712_n 0.00206439f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_420 N_D_M1004_g N_VGND_c_872_n 0.00268723f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_421 N_D_M1007_g N_VGND_c_872_n 0.00146448f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_422 N_D_M1009_g N_VGND_c_873_n 0.00146448f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_423 N_D_M1011_g N_VGND_c_873_n 0.00268723f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_424 N_D_M1007_g N_VGND_c_874_n 0.00424416f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_425 N_D_M1009_g N_VGND_c_874_n 0.00424416f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_426 N_D_M1004_g N_VGND_c_877_n 0.00422898f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_427 N_D_M1011_g N_VGND_c_878_n 0.00424416f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_428 N_D_M1004_g N_VGND_c_879_n 0.00577235f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_429 N_D_M1007_g N_VGND_c_879_n 0.00573607f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_430 N_D_M1009_g N_VGND_c_879_n 0.00573607f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_431 N_D_M1011_g N_VGND_c_879_n 0.00672653f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_432 N_D_M1004_g N_A_991_47#_c_1060_n 0.00244813f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_433 N_D_M1004_g N_A_991_47#_c_1061_n 0.00411304f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_434 N_D_M1007_g N_A_991_47#_c_1061_n 5.17008e-19 $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_435 N_D_M1004_g N_A_991_47#_c_1051_n 0.00958113f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_436 N_D_M1007_g N_A_991_47#_c_1051_n 0.00845772f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_437 D N_A_991_47#_c_1051_n 0.0298076f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_438 N_D_c_480_n N_A_991_47#_c_1051_n 0.00205431f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_439 N_D_M1004_g N_A_991_47#_c_1052_n 0.00144629f $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_440 N_D_M1004_g N_A_991_47#_c_1068_n 5.77985e-19 $X=6.97 $Y=0.56 $X2=0 $Y2=0
cc_441 N_D_M1007_g N_A_991_47#_c_1068_n 0.00655349f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_442 N_D_M1009_g N_A_991_47#_c_1068_n 0.00655349f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_443 N_D_M1011_g N_A_991_47#_c_1068_n 5.77985e-19 $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_444 N_D_M1009_g N_A_991_47#_c_1053_n 0.00850187f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_445 N_D_M1011_g N_A_991_47#_c_1053_n 0.00977142f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_446 D N_A_991_47#_c_1053_n 0.0629925f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_447 N_D_c_480_n N_A_991_47#_c_1053_n 0.00205431f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_448 N_D_c_481_n N_A_991_47#_c_1053_n 0.00740456f $X=8.47 $Y=1.16 $X2=0 $Y2=0
cc_449 N_D_M1009_g N_A_991_47#_c_1054_n 5.77896e-19 $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_450 N_D_M1011_g N_A_991_47#_c_1054_n 0.00655349f $X=8.23 $Y=0.56 $X2=0 $Y2=0
cc_451 N_D_M1007_g N_A_991_47#_c_1055_n 0.00110555f $X=7.39 $Y=0.56 $X2=0 $Y2=0
cc_452 N_D_M1009_g N_A_991_47#_c_1055_n 0.00110555f $X=7.81 $Y=0.56 $X2=0 $Y2=0
cc_453 D N_A_991_47#_c_1055_n 0.0265408f $X=8.425 $Y=1.105 $X2=0 $Y2=0
cc_454 N_D_c_480_n N_A_991_47#_c_1055_n 0.00213429f $X=8.305 $Y=1.16 $X2=0 $Y2=0
cc_455 N_VPWR_c_562_n N_Y_M1001_d 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_c_562_n N_Y_M1025_d 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_457 N_VPWR_c_562_n N_Y_M1014_d 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_562_n N_Y_M1021_d 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_562_n N_Y_M1002_s 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_562_n N_Y_M1029_s 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_461 N_VPWR_c_562_n N_Y_M1015_s 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_562_n N_Y_M1026_s 0.00215201f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_463 N_VPWR_c_576_n N_Y_c_725_n 0.0189039f $X=1.955 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_562_n N_Y_c_725_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_M1020_s N_Y_c_700_n 0.00167154f $X=1.905 $Y=1.485 $X2=0 $Y2=0
cc_466 N_VPWR_c_565_n N_Y_c_700_n 0.0129161f $X=2.04 $Y=2 $X2=0 $Y2=0
cc_467 N_VPWR_c_578_n N_Y_c_732_n 0.0189039f $X=2.795 $Y=2.72 $X2=0 $Y2=0
cc_468 N_VPWR_c_562_n N_Y_c_732_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_469 N_VPWR_c_580_n N_Y_c_735_n 0.0189039f $X=3.635 $Y=2.72 $X2=0 $Y2=0
cc_470 N_VPWR_c_562_n N_Y_c_735_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_M1016_s N_Y_c_701_n 0.00167154f $X=3.585 $Y=1.485 $X2=0 $Y2=0
cc_472 N_VPWR_c_567_n N_Y_c_701_n 0.0129161f $X=3.72 $Y=2 $X2=0 $Y2=0
cc_473 N_VPWR_c_587_n N_Y_c_754_n 0.0189039f $X=4.475 $Y=2.72 $X2=0 $Y2=0
cc_474 N_VPWR_c_562_n N_Y_c_754_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_475 N_VPWR_M1028_s N_Y_c_702_n 0.0115037f $X=4.425 $Y=1.485 $X2=0 $Y2=0
cc_476 N_VPWR_c_568_n N_Y_c_702_n 0.0559698f $X=5 $Y=2 $X2=0 $Y2=0
cc_477 N_VPWR_c_582_n N_Y_c_779_n 0.0189039f $X=5.835 $Y=2.72 $X2=0 $Y2=0
cc_478 N_VPWR_c_562_n N_Y_c_779_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_479 N_VPWR_M1022_d N_Y_c_703_n 0.00167154f $X=5.785 $Y=1.485 $X2=0 $Y2=0
cc_480 N_VPWR_c_569_n N_Y_c_703_n 0.0129161f $X=5.92 $Y=2 $X2=0 $Y2=0
cc_481 N_VPWR_c_584_n N_Y_c_786_n 0.0189039f $X=6.675 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_562_n N_Y_c_786_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_M1031_d N_Y_c_704_n 0.00167154f $X=6.625 $Y=1.485 $X2=0 $Y2=0
cc_484 N_VPWR_c_570_n N_Y_c_704_n 0.0129161f $X=6.76 $Y=2 $X2=0 $Y2=0
cc_485 N_VPWR_c_571_n N_Y_c_791_n 0.0189039f $X=7.515 $Y=2.72 $X2=0 $Y2=0
cc_486 N_VPWR_c_562_n N_Y_c_791_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_487 N_VPWR_M1023_d N_Y_c_705_n 0.00167154f $X=7.465 $Y=1.485 $X2=0 $Y2=0
cc_488 N_VPWR_c_572_n N_Y_c_705_n 0.0129161f $X=7.6 $Y=2 $X2=0 $Y2=0
cc_489 N_VPWR_c_574_n N_Y_c_706_n 0.0108343f $X=8.44 $Y=1.66 $X2=0 $Y2=0
cc_490 N_VPWR_c_588_n N_Y_c_813_n 0.0189039f $X=8.355 $Y=2.72 $X2=0 $Y2=0
cc_491 N_VPWR_c_562_n N_Y_c_813_n 0.0122217f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_492 N_VPWR_M1027_s N_Y_c_707_n 0.00167154f $X=2.745 $Y=1.485 $X2=0 $Y2=0
cc_493 N_VPWR_c_566_n N_Y_c_707_n 0.0129161f $X=2.88 $Y=2 $X2=0 $Y2=0
cc_494 N_Y_M1005_s N_VGND_c_879_n 0.00216833f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_495 N_Y_M1012_s N_VGND_c_879_n 0.00216833f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_496 N_Y_c_697_n N_A_215_47#_M1008_d 0.00162207f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_497 N_Y_c_697_n N_A_215_47#_c_973_n 0.0120104f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_498 N_Y_M1005_s N_A_215_47#_c_974_n 0.00305599f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_499 N_Y_M1012_s N_A_215_47#_c_974_n 0.00305226f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_500 N_Y_c_697_n N_A_215_47#_c_974_n 0.0447682f $X=2.375 $Y=0.77 $X2=0 $Y2=0
cc_501 N_Y_c_745_n N_A_215_47#_c_974_n 0.0154172f $X=2.507 $Y=0.905 $X2=0 $Y2=0
cc_502 N_Y_c_702_n N_A_633_47#_c_1016_n 0.00714173f $X=5.335 $Y=1.555 $X2=0
+ $Y2=0
cc_503 N_Y_c_745_n N_A_633_47#_c_1016_n 0.00943676f $X=2.507 $Y=0.905 $X2=0
+ $Y2=0
cc_504 N_Y_c_704_n N_A_991_47#_c_1051_n 0.00238597f $X=7.015 $Y=1.555 $X2=0
+ $Y2=0
cc_505 N_Y_c_704_n N_A_991_47#_c_1052_n 0.00933129f $X=7.015 $Y=1.555 $X2=0
+ $Y2=0
cc_506 N_VGND_c_879_n N_A_215_47#_M1005_d 0.00209324f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_507 N_VGND_c_879_n N_A_215_47#_M1008_d 0.00215227f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_879_n N_A_215_47#_M1019_d 0.00215227f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_879_n N_A_215_47#_M1013_s 0.00215227f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_879_n N_A_215_47#_M1018_s 0.00209344f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_871_n N_A_215_47#_c_972_n 0.0168365f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_512 N_VGND_c_877_n N_A_215_47#_c_972_n 0.0173346f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_879_n N_A_215_47#_c_972_n 0.00961661f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_871_n N_A_215_47#_c_973_n 0.00586968f $X=0.68 $Y=0.38 $X2=0
+ $Y2=0
cc_515 N_VGND_c_877_n N_A_215_47#_c_974_n 0.192442f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_879_n N_A_215_47#_c_974_n 0.122676f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_879_n N_A_633_47#_M1010_d 0.00216833f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_518 N_VGND_c_879_n N_A_633_47#_M1017_d 0.00216833f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_879_n N_A_633_47#_M1000_s 0.00216833f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_879_n N_A_633_47#_M1006_s 0.00216833f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_877_n N_A_633_47#_c_1016_n 0.00358979f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_879_n N_A_633_47#_c_1016_n 0.0118623f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_879_n N_A_991_47#_M1000_d 0.00209344f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_524 N_VGND_c_879_n N_A_991_47#_M1003_d 0.00215227f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_879_n N_A_991_47#_M1033_d 0.00215206f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_879_n N_A_991_47#_M1007_d 0.00215201f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_879_n N_A_991_47#_M1011_d 0.00209319f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_877_n N_A_991_47#_c_1050_n 0.098916f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_879_n N_A_991_47#_c_1050_n 0.0628327f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_877_n N_A_991_47#_c_1060_n 0.0152108f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_879_n N_A_991_47#_c_1060_n 0.00940698f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_M1004_s N_A_991_47#_c_1051_n 0.00169589f $X=7.045 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_VGND_c_872_n N_A_991_47#_c_1051_n 0.0111177f $X=7.18 $Y=0.38 $X2=0
+ $Y2=0
cc_534 N_VGND_c_874_n N_A_991_47#_c_1051_n 0.00193763f $X=7.935 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_c_877_n N_A_991_47#_c_1051_n 0.00193763f $X=7.095 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_879_n N_A_991_47#_c_1051_n 0.00828806f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_874_n N_A_991_47#_c_1068_n 0.0188551f $X=7.935 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_879_n N_A_991_47#_c_1068_n 0.0122069f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_M1009_s N_A_991_47#_c_1053_n 0.00169589f $X=7.885 $Y=0.235 $X2=0
+ $Y2=0
cc_540 N_VGND_c_873_n N_A_991_47#_c_1053_n 0.0111177f $X=8.02 $Y=0.38 $X2=0
+ $Y2=0
cc_541 N_VGND_c_874_n N_A_991_47#_c_1053_n 0.00193763f $X=7.935 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_c_878_n N_A_991_47#_c_1053_n 0.00193763f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_879_n N_A_991_47#_c_1053_n 0.00828806f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_878_n N_A_991_47#_c_1054_n 0.0213324f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_879_n N_A_991_47#_c_1054_n 0.0126042f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_546 N_A_215_47#_c_974_n N_A_633_47#_M1010_d 0.00305599f $X=4.56 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_547 N_A_215_47#_c_974_n N_A_633_47#_M1017_d 0.00305599f $X=4.56 $Y=0.38 $X2=0
+ $Y2=0
cc_548 N_A_215_47#_M1013_s N_A_633_47#_c_1016_n 0.00162207f $X=3.585 $Y=0.235
+ $X2=0 $Y2=0
cc_549 N_A_215_47#_M1018_s N_A_633_47#_c_1016_n 0.00321334f $X=4.425 $Y=0.235
+ $X2=0 $Y2=0
cc_550 N_A_215_47#_c_974_n N_A_633_47#_c_1016_n 0.083864f $X=4.56 $Y=0.38 $X2=0
+ $Y2=0
cc_551 N_A_215_47#_c_974_n N_A_991_47#_c_1050_n 0.0180051f $X=4.56 $Y=0.38 $X2=0
+ $Y2=0
cc_552 N_A_633_47#_c_1016_n N_A_991_47#_M1000_d 0.00321334f $X=6.34 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_553 N_A_633_47#_c_1016_n N_A_991_47#_M1003_d 0.00162207f $X=6.34 $Y=0.72
+ $X2=0 $Y2=0
cc_554 N_A_633_47#_M1000_s N_A_991_47#_c_1050_n 0.00305599f $X=5.365 $Y=0.235
+ $X2=0 $Y2=0
cc_555 N_A_633_47#_M1006_s N_A_991_47#_c_1050_n 0.00305599f $X=6.205 $Y=0.235
+ $X2=0 $Y2=0
cc_556 N_A_633_47#_c_1016_n N_A_991_47#_c_1050_n 0.083864f $X=6.34 $Y=0.72 $X2=0
+ $Y2=0
cc_557 N_A_633_47#_c_1016_n N_A_991_47#_c_1052_n 0.00799569f $X=6.34 $Y=0.72
+ $X2=0 $Y2=0

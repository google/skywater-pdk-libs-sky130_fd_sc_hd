* NGSPICE file created from sky130_fd_sc_hd__nand4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
M1000 Y a_27_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=1.08e+12p pd=1.016e+07u as=2.1392e+12p ps=1.542e+07u
M1001 VGND D a_655_47# VNB nshort w=650000u l=150000u
+  ad=2.847e+11p pd=3.2e+06u as=5.72e+11p ps=5.66e+06u
M1002 a_215_47# a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=5.135e+11p pd=5.48e+06u as=1.755e+11p ps=1.84e+06u
M1003 Y a_27_47# a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_465_47# C a_655_47# VNB nshort w=650000u l=150000u
+  ad=3.51e+11p pd=3.68e+06u as=0p ps=0u
M1005 a_655_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_465_47# B a_215_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1008 VPWR D Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_215_47# B a_465_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y D VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_655_47# C a_465_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_27_47# Y VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends


* File: sky130_fd_sc_hd__clkbuf_16.spice.SKY130_FD_SC_HD__CLKBUF_16.pxi
* Created: Thu Aug 27 14:10:41 2020
* 
x_PM_SKY130_FD_SC_HD__CLKBUF_16%A N_A_M1012_g N_A_c_151_n N_A_M1009_g
+ N_A_M1022_g N_A_c_152_n N_A_M1019_g N_A_M1026_g N_A_c_153_n N_A_M1021_g
+ N_A_M1039_g N_A_c_154_n N_A_M1038_g A A N_A_c_150_n
+ PM_SKY130_FD_SC_HD__CLKBUF_16%A
x_PM_SKY130_FD_SC_HD__CLKBUF_16%A_110_47# N_A_110_47#_M1012_d
+ N_A_110_47#_M1026_d N_A_110_47#_M1009_s N_A_110_47#_M1021_s
+ N_A_110_47#_M1002_g N_A_110_47#_M1000_g N_A_110_47#_M1003_g
+ N_A_110_47#_M1001_g N_A_110_47#_M1004_g N_A_110_47#_M1005_g
+ N_A_110_47#_M1007_g N_A_110_47#_M1006_g N_A_110_47#_M1008_g
+ N_A_110_47#_M1010_g N_A_110_47#_M1015_g N_A_110_47#_M1011_g
+ N_A_110_47#_M1017_g N_A_110_47#_M1013_g N_A_110_47#_M1018_g
+ N_A_110_47#_M1014_g N_A_110_47#_M1020_g N_A_110_47#_M1016_g
+ N_A_110_47#_M1023_g N_A_110_47#_M1024_g N_A_110_47#_M1029_g
+ N_A_110_47#_M1025_g N_A_110_47#_M1031_g N_A_110_47#_M1027_g
+ N_A_110_47#_M1032_g N_A_110_47#_M1028_g N_A_110_47#_M1033_g
+ N_A_110_47#_M1030_g N_A_110_47#_M1036_g N_A_110_47#_M1034_g
+ N_A_110_47#_c_224_n N_A_110_47#_M1037_g N_A_110_47#_M1035_g
+ N_A_110_47#_c_226_n N_A_110_47#_c_246_n N_A_110_47#_c_259_n
+ N_A_110_47#_c_227_n N_A_110_47#_c_247_n N_A_110_47#_c_228_n
+ N_A_110_47#_c_267_n N_A_110_47#_c_269_n
+ PM_SKY130_FD_SC_HD__CLKBUF_16%A_110_47#
x_PM_SKY130_FD_SC_HD__CLKBUF_16%VPWR N_VPWR_M1009_d N_VPWR_M1019_d
+ N_VPWR_M1038_d N_VPWR_M1001_s N_VPWR_M1006_s N_VPWR_M1011_s N_VPWR_M1014_s
+ N_VPWR_M1024_s N_VPWR_M1027_s N_VPWR_M1030_s N_VPWR_M1035_s N_VPWR_c_498_n
+ N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n
+ N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n VPWR
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_497_n
+ PM_SKY130_FD_SC_HD__CLKBUF_16%VPWR
x_PM_SKY130_FD_SC_HD__CLKBUF_16%X N_X_M1002_s N_X_M1004_s N_X_M1008_s
+ N_X_M1017_s N_X_M1020_s N_X_M1029_s N_X_M1032_s N_X_M1036_s N_X_M1000_d
+ N_X_M1005_d N_X_M1010_d N_X_M1013_d N_X_M1016_d N_X_M1025_d N_X_M1028_d
+ N_X_M1034_d N_X_c_642_n N_X_c_643_n N_X_c_644_n N_X_c_678_n N_X_c_645_n
+ N_X_c_646_n N_X_c_688_n N_X_c_647_n N_X_c_648_n N_X_c_698_n N_X_c_649_n
+ N_X_c_650_n N_X_c_709_n N_X_c_651_n N_X_c_652_n N_X_c_719_n N_X_c_653_n
+ N_X_c_654_n N_X_c_729_n N_X_c_655_n N_X_c_656_n N_X_c_657_n N_X_c_739_n
+ N_X_c_658_n N_X_c_743_n N_X_c_659_n N_X_c_747_n N_X_c_660_n N_X_c_752_n
+ N_X_c_661_n N_X_c_757_n N_X_c_662_n N_X_c_762_n N_X_c_663_n X X X X
+ N_X_c_666_n PM_SKY130_FD_SC_HD__CLKBUF_16%X
x_PM_SKY130_FD_SC_HD__CLKBUF_16%VGND N_VGND_M1012_s N_VGND_M1022_s
+ N_VGND_M1039_s N_VGND_M1003_d N_VGND_M1007_d N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1023_d N_VGND_M1031_d N_VGND_M1033_d N_VGND_M1037_d N_VGND_c_873_n
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n
+ N_VGND_c_879_n N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n N_VGND_c_883_n
+ N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n N_VGND_c_888_n
+ N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n
+ N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n VGND
+ N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n N_VGND_c_901_n N_VGND_c_902_n
+ N_VGND_c_903_n N_VGND_c_904_n N_VGND_c_905_n
+ PM_SKY130_FD_SC_HD__CLKBUF_16%VGND
cc_1 VNB N_A_M1012_g 0.0293898f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_M1022_g 0.0229781f $X=-0.19 $Y=-0.24 $X2=0.905 $Y2=0.445
cc_3 VNB N_A_M1026_g 0.0229774f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.445
cc_4 VNB N_A_M1039_g 0.0234436f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.445
cc_5 VNB A 0.0236322f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_150_n 0.109553f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.155
cc_7 VNB N_A_110_47#_M1002_g 0.0260664f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=0.9
cc_8 VNB N_A_110_47#_M1003_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=0.445
cc_9 VNB N_A_110_47#_M1004_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_110_47#_M1007_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.155
cc_11 VNB N_A_110_47#_M1008_g 0.0241433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_110_47#_M1015_g 0.0241428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1017_g 0.0238169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_M1018_g 0.0240545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_M1020_g 0.0240466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_110_47#_M1023_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_110_47#_M1029_g 0.0241355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_110_47#_M1031_g 0.0241431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_110_47#_M1032_g 0.0241328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_110_47#_M1033_g 0.0241116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_110_47#_M1036_g 0.0237673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_110_47#_c_224_n 0.300055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_110_47#_M1037_g 0.0320587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_110_47#_c_226_n 0.00439944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_110_47#_c_227_n 0.00481736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_110_47#_c_228_n 0.00429043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_497_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_642_n 0.00160391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_643_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_644_n 0.00419804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_645_n 0.00126237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_646_n 0.00514258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_647_n 0.00125415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_648_n 0.00501892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_649_n 6.22964e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_650_n 0.00491776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_651_n 0.00125437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_652_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_653_n 0.00126258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_654_n 0.00522562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_655_n 0.00126798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_656_n 4.84646e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_657_n 0.00137779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_658_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_659_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_X_c_660_n 0.00217463f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_661_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_662_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_663_n 0.00207149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB X 0.0318745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_873_n 0.0107531f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_52 VNB N_VGND_c_874_n 0.0190761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_875_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.155
cc_54 VNB N_VGND_c_876_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_877_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_878_n 0.00400996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_879_n 0.00390627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_880_n 0.0157899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_881_n 0.00395785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_882_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_883_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_884_n 0.00397944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_885_n 0.00402207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_886_n 0.0135264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_887_n 0.0178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_888_n 0.0167416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_889_n 0.00500104f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_890_n 0.0160902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_891_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_892_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_893_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_894_n 0.0154623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_895_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_896_n 0.0157075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_897_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_898_n 0.0167416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_899_n 0.0157442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_900_n 0.0154599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_901_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_902_n 0.0046855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_903_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_904_n 0.00478165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_905_n 0.430355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VPB N_A_c_151_n 0.0192408f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.41
cc_85 VPB N_A_c_152_n 0.0143973f $X=-0.19 $Y=1.305 $X2=0.905 $Y2=1.41
cc_86 VPB N_A_c_153_n 0.0143972f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.41
cc_87 VPB N_A_c_154_n 0.0145802f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.41
cc_88 VPB A 0.00127249f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_89 VPB N_A_c_150_n 0.0444013f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.155
cc_90 VPB N_A_110_47#_M1000_g 0.0190615f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.41
cc_91 VPB N_A_110_47#_M1001_g 0.0187483f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.985
cc_92 VPB N_A_110_47#_M1005_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_93 VPB N_A_110_47#_M1006_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_110_47#_M1010_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_110_47#_M1011_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_110_47#_M1013_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_110_47#_M1014_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_A_110_47#_M1016_g 0.0186881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_110_47#_M1024_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_110_47#_M1025_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_110_47#_M1027_g 0.0187483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_110_47#_M1028_g 0.0187387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_110_47#_M1030_g 0.0186963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_110_47#_M1034_g 0.0173762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_110_47#_c_224_n 0.0522358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_110_47#_M1035_g 0.0224494f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_110_47#_c_246_n 0.00130522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_110_47#_c_247_n 0.00130663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_110_47#_c_228_n 0.00459688f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_498_n 0.0108797f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_111 VPB N_VPWR_c_499_n 0.0303682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_500_n 0.00397494f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.155
cc_113 VPB N_VPWR_c_501_n 0.0038747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_502_n 0.0038747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_503_n 0.0038747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_504_n 0.0038747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_505_n 0.0167159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_506_n 0.00381264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_507_n 0.0171833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_508_n 0.00383029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_509_n 0.00383029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_510_n 0.00390012f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_511_n 0.012949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_512_n 0.0275421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_513_n 0.0167191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_514_n 0.00506696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_515_n 0.0167159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_516_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_517_n 0.0167159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_518_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_519_n 0.0167159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_520_n 0.00502323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_521_n 0.0171833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_522_n 0.00497107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_523_n 0.0167435f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_524_n 0.0171833f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_525_n 0.0172466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_526_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_527_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_528_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_529_n 0.00473193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_497_n 0.0471568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB X 0.0102708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_X_c_666_n 0.00995053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 N_A_M1039_g N_A_110_47#_M1002_g 0.0222446f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_c_154_n N_A_110_47#_M1000_g 0.0222446f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_150_n N_A_110_47#_c_224_n 0.0222446f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_148 N_A_M1012_g N_A_110_47#_c_226_n 0.00404849f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_M1022_g N_A_110_47#_c_226_n 0.00359298f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_150 A N_A_110_47#_c_226_n 0.0237393f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_151 N_A_c_150_n N_A_110_47#_c_226_n 0.0135245f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_152 N_A_c_151_n N_A_110_47#_c_246_n 0.00324761f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_152_n N_A_110_47#_c_246_n 0.00234025f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_150_n N_A_110_47#_c_246_n 0.0103199f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_155 N_A_c_150_n N_A_110_47#_c_259_n 0.0576342f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_156 N_A_M1026_g N_A_110_47#_c_227_n 0.00352135f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_M1039_g N_A_110_47#_c_227_n 0.00356184f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_c_150_n N_A_110_47#_c_227_n 0.0139367f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_159 N_A_c_153_n N_A_110_47#_c_247_n 0.00216105f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_154_n N_A_110_47#_c_247_n 0.00314608f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_150_n N_A_110_47#_c_247_n 0.00809327f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_162 N_A_c_150_n N_A_110_47#_c_228_n 0.0213857f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_163 A N_A_110_47#_c_267_n 0.0198893f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_164 N_A_c_150_n N_A_110_47#_c_267_n 0.00950927f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_165 N_A_c_150_n N_A_110_47#_c_269_n 0.00588528f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_166 N_A_c_151_n N_VPWR_c_499_n 0.00341694f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_167 A N_VPWR_c_499_n 0.0100578f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A_c_150_n N_VPWR_c_499_n 0.00611048f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_169 N_A_c_152_n N_VPWR_c_500_n 0.00161372f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_153_n N_VPWR_c_500_n 0.00161372f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_150_n N_VPWR_c_500_n 0.00223472f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_172 N_A_c_154_n N_VPWR_c_501_n 0.00161372f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_153_n N_VPWR_c_513_n 0.00585385f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_154_n N_VPWR_c_513_n 0.00585385f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_151_n N_VPWR_c_523_n 0.00585385f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_152_n N_VPWR_c_523_n 0.00585385f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_151_n N_VPWR_c_497_n 0.0114221f $X=0.475 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_152_n N_VPWR_c_497_n 0.0104895f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_153_n N_VPWR_c_497_n 0.0105664f $X=1.335 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_154_n N_VPWR_c_497_n 0.0105915f $X=1.765 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_M1012_g N_VGND_c_874_n 0.0038241f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_182 A N_VGND_c_874_n 0.0245931f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_183 N_A_c_150_n N_VGND_c_874_n 0.00149294f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_184 N_A_M1022_g N_VGND_c_875_n 0.00168046f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_M1026_g N_VGND_c_875_n 0.00168046f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A_c_150_n N_VGND_c_875_n 0.00255763f $X=1.765 $Y=1.155 $X2=0 $Y2=0
cc_187 N_A_M1039_g N_VGND_c_876_n 0.00170359f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_M1026_g N_VGND_c_888_n 0.00585385f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_M1039_g N_VGND_c_888_n 0.00585385f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_M1012_g N_VGND_c_898_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A_M1022_g N_VGND_c_898_n 0.00585385f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_M1012_g N_VGND_c_905_n 0.011499f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_M1022_g N_VGND_c_905_n 0.010643f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_M1026_g N_VGND_c_905_n 0.010643f $X=1.335 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_M1039_g N_VGND_c_905_n 0.0106694f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_196 A N_VGND_c_905_n 0.00157507f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_197 N_A_110_47#_c_259_n N_VPWR_c_500_n 0.0071967f $X=1.43 $Y=1.2 $X2=0 $Y2=0
cc_198 N_A_110_47#_M1000_g N_VPWR_c_501_n 0.00161372f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_110_47#_c_228_n N_VPWR_c_501_n 0.0081125f $X=7.505 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_110_47#_M1001_g N_VPWR_c_502_n 0.00248982f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_110_47#_M1005_g N_VPWR_c_502_n 0.00248982f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_202 N_A_110_47#_M1006_g N_VPWR_c_503_n 0.00248982f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_203 N_A_110_47#_M1010_g N_VPWR_c_503_n 0.00248982f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_204 N_A_110_47#_M1011_g N_VPWR_c_504_n 0.00248982f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_110_47#_M1013_g N_VPWR_c_504_n 0.00248982f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_110_47#_M1013_g N_VPWR_c_505_n 0.00591536f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_110_47#_M1014_g N_VPWR_c_505_n 0.00591536f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_208 N_A_110_47#_M1014_g N_VPWR_c_506_n 0.00245982f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_110_47#_M1016_g N_VPWR_c_506_n 0.00241885f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_110_47#_M1016_g N_VPWR_c_507_n 0.00591536f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_211 N_A_110_47#_M1024_g N_VPWR_c_507_n 0.00591536f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_212 N_A_110_47#_M1024_g N_VPWR_c_508_n 0.00247084f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_213 N_A_110_47#_M1025_g N_VPWR_c_508_n 0.00244044f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_214 N_A_110_47#_M1027_g N_VPWR_c_509_n 0.00247084f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_215 N_A_110_47#_M1028_g N_VPWR_c_509_n 0.00244044f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_216 N_A_110_47#_M1030_g N_VPWR_c_510_n 0.0024762f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_217 N_A_110_47#_M1034_g N_VPWR_c_510_n 0.00252673f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_218 N_A_110_47#_c_224_n N_VPWR_c_510_n 3.54728e-19 $X=8.64 $Y=0.95 $X2=0
+ $Y2=0
cc_219 N_A_110_47#_M1035_g N_VPWR_c_512_n 0.00722026f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_220 N_A_110_47#_c_247_n N_VPWR_c_513_n 0.0141362f $X=1.55 $Y=1.92 $X2=0 $Y2=0
cc_221 N_A_110_47#_M1000_g N_VPWR_c_515_n 0.00591536f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_222 N_A_110_47#_M1001_g N_VPWR_c_515_n 0.00591536f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A_110_47#_M1005_g N_VPWR_c_517_n 0.00591536f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_110_47#_M1006_g N_VPWR_c_517_n 0.00591536f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_110_47#_M1010_g N_VPWR_c_519_n 0.00591536f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_110_47#_M1011_g N_VPWR_c_519_n 0.00591536f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_110_47#_M1028_g N_VPWR_c_521_n 0.00591536f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_110_47#_M1030_g N_VPWR_c_521_n 0.00591536f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_229 N_A_110_47#_c_246_n N_VPWR_c_523_n 0.0144053f $X=0.69 $Y=1.96 $X2=0 $Y2=0
cc_230 N_A_110_47#_M1025_g N_VPWR_c_524_n 0.00591536f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_110_47#_M1027_g N_VPWR_c_524_n 0.00591536f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_232 N_A_110_47#_M1034_g N_VPWR_c_525_n 0.00585385f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_233 N_A_110_47#_M1035_g N_VPWR_c_525_n 0.00556673f $X=8.64 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_110_47#_M1009_s N_VPWR_c_497_n 0.00344736f $X=0.55 $Y=1.485 $X2=0
+ $Y2=0
cc_235 N_A_110_47#_M1021_s N_VPWR_c_497_n 0.00336062f $X=1.41 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_A_110_47#_M1000_g N_VPWR_c_497_n 0.0105781f $X=2.195 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_110_47#_M1001_g N_VPWR_c_497_n 0.0106294f $X=2.625 $Y=1.985 $X2=0
+ $Y2=0
cc_238 N_A_110_47#_M1005_g N_VPWR_c_497_n 0.0106294f $X=3.055 $Y=1.985 $X2=0
+ $Y2=0
cc_239 N_A_110_47#_M1006_g N_VPWR_c_497_n 0.0106294f $X=3.485 $Y=1.985 $X2=0
+ $Y2=0
cc_240 N_A_110_47#_M1010_g N_VPWR_c_497_n 0.0106294f $X=3.915 $Y=1.985 $X2=0
+ $Y2=0
cc_241 N_A_110_47#_M1011_g N_VPWR_c_497_n 0.0106294f $X=4.345 $Y=1.985 $X2=0
+ $Y2=0
cc_242 N_A_110_47#_M1013_g N_VPWR_c_497_n 0.0106294f $X=4.775 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_110_47#_M1014_g N_VPWR_c_497_n 0.0106158f $X=5.205 $Y=1.985 $X2=0
+ $Y2=0
cc_244 N_A_110_47#_M1016_g N_VPWR_c_497_n 0.0106386f $X=5.63 $Y=1.985 $X2=0
+ $Y2=0
cc_245 N_A_110_47#_M1024_g N_VPWR_c_497_n 0.0106408f $X=6.06 $Y=1.985 $X2=0
+ $Y2=0
cc_246 N_A_110_47#_M1025_g N_VPWR_c_497_n 0.0106522f $X=6.49 $Y=1.985 $X2=0
+ $Y2=0
cc_247 N_A_110_47#_M1027_g N_VPWR_c_497_n 0.0106408f $X=6.92 $Y=1.985 $X2=0
+ $Y2=0
cc_248 N_A_110_47#_M1028_g N_VPWR_c_497_n 0.0106522f $X=7.35 $Y=1.985 $X2=0
+ $Y2=0
cc_249 N_A_110_47#_M1030_g N_VPWR_c_497_n 0.0106408f $X=7.78 $Y=1.985 $X2=0
+ $Y2=0
cc_250 N_A_110_47#_M1034_g N_VPWR_c_497_n 0.0106428f $X=8.21 $Y=1.985 $X2=0
+ $Y2=0
cc_251 N_A_110_47#_M1035_g N_VPWR_c_497_n 0.011058f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_252 N_A_110_47#_c_246_n N_VPWR_c_497_n 0.00935836f $X=0.69 $Y=1.96 $X2=0
+ $Y2=0
cc_253 N_A_110_47#_c_247_n N_VPWR_c_497_n 0.00952853f $X=1.55 $Y=1.92 $X2=0
+ $Y2=0
cc_254 N_A_110_47#_M1002_g N_X_c_642_n 0.00120255f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_255 N_A_110_47#_M1003_g N_X_c_642_n 0.00120255f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_256 N_A_110_47#_c_227_n N_X_c_642_n 0.00257148f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_257 N_A_110_47#_M1003_g N_X_c_643_n 0.0119364f $X=2.625 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A_110_47#_M1004_g N_X_c_643_n 0.0122327f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_110_47#_c_224_n N_X_c_643_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_260 N_A_110_47#_c_228_n N_X_c_643_n 0.0429599f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_110_47#_M1002_g N_X_c_644_n 0.00289158f $X=2.195 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_110_47#_c_224_n N_X_c_644_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_263 N_A_110_47#_c_227_n N_X_c_644_n 0.00599637f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_110_47#_c_228_n N_X_c_644_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_110_47#_M1001_g N_X_c_678_n 0.0151109f $X=2.625 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A_110_47#_M1005_g N_X_c_678_n 0.015045f $X=3.055 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A_110_47#_c_224_n N_X_c_678_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_268 N_A_110_47#_c_228_n N_X_c_678_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_110_47#_M1004_g N_X_c_645_n 0.00120255f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_110_47#_M1007_g N_X_c_645_n 0.00120255f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_271 N_A_110_47#_M1007_g N_X_c_646_n 0.0122792f $X=3.485 $Y=0.445 $X2=0 $Y2=0
cc_272 N_A_110_47#_M1008_g N_X_c_646_n 0.0122792f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_273 N_A_110_47#_c_224_n N_X_c_646_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_274 N_A_110_47#_c_228_n N_X_c_646_n 0.0429599f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_110_47#_M1006_g N_X_c_688_n 0.0151109f $X=3.485 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_110_47#_M1010_g N_X_c_688_n 0.0151109f $X=3.915 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_110_47#_c_224_n N_X_c_688_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_278 N_A_110_47#_c_228_n N_X_c_688_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_110_47#_M1008_g N_X_c_647_n 0.00120255f $X=3.915 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_110_47#_M1015_g N_X_c_647_n 0.00118828f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_281 N_A_110_47#_M1015_g N_X_c_648_n 0.0122792f $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_110_47#_M1017_g N_X_c_648_n 0.00994201f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_283 N_A_110_47#_c_224_n N_X_c_648_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_284 N_A_110_47#_c_228_n N_X_c_648_n 0.0418783f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_110_47#_M1011_g N_X_c_698_n 0.0151109f $X=4.345 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A_110_47#_M1013_g N_X_c_698_n 0.0150553f $X=4.775 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_110_47#_c_224_n N_X_c_698_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_288 N_A_110_47#_c_228_n N_X_c_698_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_110_47#_M1015_g N_X_c_649_n 5.05907e-19 $X=4.345 $Y=0.445 $X2=0 $Y2=0
cc_290 N_A_110_47#_M1017_g N_X_c_649_n 0.0062908f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_291 N_A_110_47#_M1018_g N_X_c_649_n 0.00119799f $X=5.205 $Y=0.445 $X2=0 $Y2=0
cc_292 N_A_110_47#_M1018_g N_X_c_650_n 0.0122482f $X=5.205 $Y=0.445 $X2=0 $Y2=0
cc_293 N_A_110_47#_M1020_g N_X_c_650_n 0.0101865f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_294 N_A_110_47#_c_224_n N_X_c_650_n 0.00253724f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_295 N_A_110_47#_c_228_n N_X_c_650_n 0.0418596f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_110_47#_M1014_g N_X_c_709_n 0.015067f $X=5.205 $Y=1.985 $X2=0 $Y2=0
cc_297 N_A_110_47#_M1016_g N_X_c_709_n 0.015067f $X=5.63 $Y=1.985 $X2=0 $Y2=0
cc_298 N_A_110_47#_c_224_n N_X_c_709_n 0.00220405f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_299 N_A_110_47#_c_228_n N_X_c_709_n 0.0378421f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_110_47#_M1020_g N_X_c_651_n 0.00121272f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_301 N_A_110_47#_M1023_g N_X_c_651_n 0.00117849f $X=6.06 $Y=0.445 $X2=0 $Y2=0
cc_302 N_A_110_47#_M1023_g N_X_c_652_n 0.0122792f $X=6.06 $Y=0.445 $X2=0 $Y2=0
cc_303 N_A_110_47#_M1029_g N_X_c_652_n 0.0102175f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_304 N_A_110_47#_c_224_n N_X_c_652_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_305 N_A_110_47#_c_228_n N_X_c_652_n 0.0429636f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_110_47#_M1024_g N_X_c_719_n 0.0151109f $X=6.06 $Y=1.985 $X2=0 $Y2=0
cc_307 N_A_110_47#_M1025_g N_X_c_719_n 0.0151109f $X=6.49 $Y=1.985 $X2=0 $Y2=0
cc_308 N_A_110_47#_c_224_n N_X_c_719_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_309 N_A_110_47#_c_228_n N_X_c_719_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_110_47#_M1029_g N_X_c_653_n 0.00122723f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_311 N_A_110_47#_M1031_g N_X_c_653_n 0.00117849f $X=6.92 $Y=0.445 $X2=0 $Y2=0
cc_312 N_A_110_47#_M1031_g N_X_c_654_n 0.0122792f $X=6.92 $Y=0.445 $X2=0 $Y2=0
cc_313 N_A_110_47#_M1032_g N_X_c_654_n 0.0102175f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_314 N_A_110_47#_c_224_n N_X_c_654_n 0.00267078f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_315 N_A_110_47#_c_228_n N_X_c_654_n 0.0429636f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_110_47#_M1027_g N_X_c_729_n 0.015107f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_317 N_A_110_47#_M1028_g N_X_c_729_n 0.0151109f $X=7.35 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A_110_47#_c_224_n N_X_c_729_n 0.00232005f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_319 N_A_110_47#_c_228_n N_X_c_729_n 0.0385727f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_110_47#_M1032_g N_X_c_655_n 0.00122723f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_321 N_A_110_47#_M1033_g N_X_c_655_n 0.00118774f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_322 N_A_110_47#_M1033_g N_X_c_656_n 0.0141891f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_323 N_A_110_47#_c_228_n N_X_c_656_n 3.30399e-19 $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_110_47#_M1036_g N_X_c_657_n 0.00121196f $X=8.21 $Y=0.445 $X2=0 $Y2=0
cc_325 N_A_110_47#_M1037_g N_X_c_657_n 0.00221636f $X=8.64 $Y=0.445 $X2=0 $Y2=0
cc_326 N_A_110_47#_c_224_n N_X_c_739_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_327 N_A_110_47#_c_228_n N_X_c_739_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_110_47#_c_224_n N_X_c_658_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_329 N_A_110_47#_c_228_n N_X_c_658_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_330 N_A_110_47#_c_224_n N_X_c_743_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_331 N_A_110_47#_c_228_n N_X_c_743_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_110_47#_c_224_n N_X_c_659_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_333 N_A_110_47#_c_228_n N_X_c_659_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_334 N_A_110_47#_c_224_n N_X_c_747_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_335 N_A_110_47#_c_228_n N_X_c_747_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_110_47#_M1017_g N_X_c_660_n 0.00211052f $X=4.775 $Y=0.445 $X2=0 $Y2=0
cc_337 N_A_110_47#_c_224_n N_X_c_660_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_338 N_A_110_47#_c_228_n N_X_c_660_n 0.0225791f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_339 N_A_110_47#_c_224_n N_X_c_752_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_340 N_A_110_47#_c_228_n N_X_c_752_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_110_47#_M1020_g N_X_c_661_n 0.00203048f $X=5.63 $Y=0.445 $X2=0 $Y2=0
cc_342 N_A_110_47#_c_224_n N_X_c_661_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_343 N_A_110_47#_c_228_n N_X_c_661_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_344 N_A_110_47#_c_224_n N_X_c_757_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_345 N_A_110_47#_c_228_n N_X_c_757_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_346 N_A_110_47#_M1029_g N_X_c_662_n 0.00203048f $X=6.49 $Y=0.445 $X2=0 $Y2=0
cc_347 N_A_110_47#_c_224_n N_X_c_662_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_348 N_A_110_47#_c_228_n N_X_c_662_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A_110_47#_c_224_n N_X_c_762_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_350 N_A_110_47#_c_228_n N_X_c_762_n 0.0168441f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A_110_47#_M1032_g N_X_c_663_n 0.00203048f $X=7.35 $Y=0.445 $X2=0 $Y2=0
cc_352 N_A_110_47#_c_224_n N_X_c_663_n 0.00277135f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_353 N_A_110_47#_c_228_n N_X_c_663_n 0.0213686f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A_110_47#_M1033_g X 0.00147955f $X=7.78 $Y=0.445 $X2=0 $Y2=0
cc_355 N_A_110_47#_M1030_g X 0.00539328f $X=7.78 $Y=1.985 $X2=0 $Y2=0
cc_356 N_A_110_47#_M1036_g X 0.011848f $X=8.21 $Y=0.445 $X2=0 $Y2=0
cc_357 N_A_110_47#_M1034_g X 0.00605481f $X=8.21 $Y=1.985 $X2=0 $Y2=0
cc_358 N_A_110_47#_c_224_n X 0.0567372f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_359 N_A_110_47#_M1037_g X 0.0136957f $X=8.64 $Y=0.445 $X2=0 $Y2=0
cc_360 N_A_110_47#_M1035_g X 0.00773738f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_361 N_A_110_47#_c_228_n X 0.0208936f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A_110_47#_M1030_g N_X_c_666_n 0.0165955f $X=7.78 $Y=1.985 $X2=0 $Y2=0
cc_363 N_A_110_47#_M1034_g N_X_c_666_n 0.0135796f $X=8.21 $Y=1.985 $X2=0 $Y2=0
cc_364 N_A_110_47#_c_224_n N_X_c_666_n 0.00238948f $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_365 N_A_110_47#_M1035_g N_X_c_666_n 0.0295096f $X=8.64 $Y=1.985 $X2=0 $Y2=0
cc_366 N_A_110_47#_c_228_n N_X_c_666_n 0.0170247f $X=7.505 $Y=1.16 $X2=0 $Y2=0
cc_367 N_A_110_47#_c_259_n N_VGND_c_875_n 0.00764914f $X=1.43 $Y=1.2 $X2=0 $Y2=0
cc_368 N_A_110_47#_M1002_g N_VGND_c_876_n 0.00170359f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_369 N_A_110_47#_c_228_n N_VGND_c_876_n 0.0091835f $X=7.505 $Y=1.16 $X2=0
+ $Y2=0
cc_370 N_A_110_47#_M1003_g N_VGND_c_877_n 0.00161372f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_110_47#_M1004_g N_VGND_c_877_n 0.00161372f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_110_47#_M1007_g N_VGND_c_878_n 0.00161372f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_373 N_A_110_47#_M1008_g N_VGND_c_878_n 0.00161372f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_110_47#_M1015_g N_VGND_c_879_n 0.00160579f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_375 N_A_110_47#_M1017_g N_VGND_c_879_n 0.0015619f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_110_47#_M1017_g N_VGND_c_880_n 0.00438144f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_110_47#_M1018_g N_VGND_c_880_n 0.00439206f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_110_47#_M1018_g N_VGND_c_881_n 0.00161724f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_110_47#_M1020_g N_VGND_c_881_n 0.00156827f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_380 N_A_110_47#_M1020_g N_VGND_c_882_n 0.00439206f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_381 N_A_110_47#_M1023_g N_VGND_c_882_n 0.00439206f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_A_110_47#_M1023_g N_VGND_c_883_n 0.00162174f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_110_47#_M1029_g N_VGND_c_883_n 0.00157905f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_384 N_A_110_47#_M1031_g N_VGND_c_884_n 0.00162174f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_110_47#_M1032_g N_VGND_c_884_n 0.00157905f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_110_47#_M1033_g N_VGND_c_885_n 0.00162705f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_110_47#_M1036_g N_VGND_c_885_n 0.00161372f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_110_47#_c_224_n N_VGND_c_885_n 4.7914e-19 $X=8.64 $Y=0.95 $X2=0 $Y2=0
cc_389 N_A_110_47#_M1037_g N_VGND_c_887_n 0.00341923f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_110_47#_c_227_n N_VGND_c_888_n 0.0137163f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_A_110_47#_M1002_g N_VGND_c_890_n 0.00585385f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_392 N_A_110_47#_M1003_g N_VGND_c_890_n 0.00439206f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_393 N_A_110_47#_M1004_g N_VGND_c_892_n 0.00439206f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_394 N_A_110_47#_M1007_g N_VGND_c_892_n 0.00439206f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_110_47#_M1008_g N_VGND_c_894_n 0.00439206f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_A_110_47#_M1015_g N_VGND_c_894_n 0.00439206f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_A_110_47#_M1032_g N_VGND_c_896_n 0.00439206f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_110_47#_M1033_g N_VGND_c_896_n 0.00439206f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_399 N_A_110_47#_c_226_n N_VGND_c_898_n 0.0137163f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_400 N_A_110_47#_M1029_g N_VGND_c_899_n 0.00439206f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_110_47#_M1031_g N_VGND_c_899_n 0.00439206f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_402 N_A_110_47#_M1036_g N_VGND_c_900_n 0.00439071f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_403 N_A_110_47#_M1037_g N_VGND_c_900_n 0.00439071f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_A_110_47#_M1012_d N_VGND_c_905_n 0.00336236f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_405 N_A_110_47#_M1026_d N_VGND_c_905_n 0.00336236f $X=1.41 $Y=0.235 $X2=0
+ $Y2=0
cc_406 N_A_110_47#_M1002_g N_VGND_c_905_n 0.0106694f $X=2.195 $Y=0.445 $X2=0
+ $Y2=0
cc_407 N_A_110_47#_M1003_g N_VGND_c_905_n 0.00590932f $X=2.625 $Y=0.445 $X2=0
+ $Y2=0
cc_408 N_A_110_47#_M1004_g N_VGND_c_905_n 0.00590932f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_409 N_A_110_47#_M1007_g N_VGND_c_905_n 0.00590932f $X=3.485 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_110_47#_M1008_g N_VGND_c_905_n 0.00590932f $X=3.915 $Y=0.445 $X2=0
+ $Y2=0
cc_411 N_A_110_47#_M1015_g N_VGND_c_905_n 0.00590932f $X=4.345 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_A_110_47#_M1017_g N_VGND_c_905_n 0.00587292f $X=4.775 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_110_47#_M1018_g N_VGND_c_905_n 0.00589619f $X=5.205 $Y=0.445 $X2=0
+ $Y2=0
cc_414 N_A_110_47#_M1020_g N_VGND_c_905_n 0.00592128f $X=5.63 $Y=0.445 $X2=0
+ $Y2=0
cc_415 N_A_110_47#_M1023_g N_VGND_c_905_n 0.00590932f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_416 N_A_110_47#_M1029_g N_VGND_c_905_n 0.00593441f $X=6.49 $Y=0.445 $X2=0
+ $Y2=0
cc_417 N_A_110_47#_M1031_g N_VGND_c_905_n 0.00590932f $X=6.92 $Y=0.445 $X2=0
+ $Y2=0
cc_418 N_A_110_47#_M1032_g N_VGND_c_905_n 0.00593441f $X=7.35 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_110_47#_M1033_g N_VGND_c_905_n 0.00590932f $X=7.78 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_A_110_47#_M1036_g N_VGND_c_905_n 0.00590684f $X=8.21 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_110_47#_M1037_g N_VGND_c_905_n 0.00691049f $X=8.64 $Y=0.445 $X2=0
+ $Y2=0
cc_422 N_A_110_47#_c_226_n N_VGND_c_905_n 0.00950576f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_423 N_A_110_47#_c_227_n N_VGND_c_905_n 0.00950576f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_497_n N_X_M1000_d 0.00301352f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_425 N_VPWR_c_497_n N_X_M1005_d 0.00301352f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_497_n N_X_M1010_d 0.00301352f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_497_n N_X_M1013_d 0.00301352f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_497_n N_X_M1016_d 0.00297078f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_c_497_n N_X_M1025_d 0.00297078f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_430 N_VPWR_c_497_n N_X_M1028_d 0.00297078f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_c_497_n N_X_M1034_d 0.00263171f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_M1001_s N_X_c_678_n 0.00334014f $X=2.7 $Y=1.485 $X2=0 $Y2=0
cc_433 N_VPWR_c_502_n N_X_c_678_n 0.0138265f $X=2.84 $Y=2.22 $X2=0 $Y2=0
cc_434 N_VPWR_M1006_s N_X_c_688_n 0.00334014f $X=3.56 $Y=1.485 $X2=0 $Y2=0
cc_435 N_VPWR_c_503_n N_X_c_688_n 0.0138265f $X=3.7 $Y=2.22 $X2=0 $Y2=0
cc_436 N_VPWR_M1011_s N_X_c_698_n 0.00334014f $X=4.42 $Y=1.485 $X2=0 $Y2=0
cc_437 N_VPWR_c_504_n N_X_c_698_n 0.0138265f $X=4.56 $Y=2.22 $X2=0 $Y2=0
cc_438 N_VPWR_M1014_s N_X_c_709_n 0.00324413f $X=5.28 $Y=1.485 $X2=0 $Y2=0
cc_439 N_VPWR_c_506_n N_X_c_709_n 0.0134101f $X=5.42 $Y=2.22 $X2=0 $Y2=0
cc_440 N_VPWR_M1024_s N_X_c_719_n 0.00334014f $X=6.135 $Y=1.485 $X2=0 $Y2=0
cc_441 N_VPWR_c_508_n N_X_c_719_n 0.0138265f $X=6.275 $Y=2.22 $X2=0 $Y2=0
cc_442 N_VPWR_M1027_s N_X_c_729_n 0.00334014f $X=6.995 $Y=1.485 $X2=0 $Y2=0
cc_443 N_VPWR_c_509_n N_X_c_729_n 0.0138265f $X=7.135 $Y=2.22 $X2=0 $Y2=0
cc_444 N_VPWR_c_515_n N_X_c_739_n 0.0149478f $X=2.71 $Y=2.717 $X2=0 $Y2=0
cc_445 N_VPWR_c_497_n N_X_c_739_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_517_n N_X_c_743_n 0.0149478f $X=3.57 $Y=2.717 $X2=0 $Y2=0
cc_447 N_VPWR_c_497_n N_X_c_743_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_519_n N_X_c_747_n 0.0149478f $X=4.43 $Y=2.717 $X2=0 $Y2=0
cc_449 N_VPWR_c_497_n N_X_c_747_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_505_n N_X_c_752_n 0.0149478f $X=5.29 $Y=2.717 $X2=0 $Y2=0
cc_451 N_VPWR_c_497_n N_X_c_752_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_452 N_VPWR_c_507_n N_X_c_757_n 0.0149478f $X=6.15 $Y=2.717 $X2=0 $Y2=0
cc_453 N_VPWR_c_497_n N_X_c_757_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_c_524_n N_X_c_762_n 0.0149478f $X=7.01 $Y=2.717 $X2=0 $Y2=0
cc_455 N_VPWR_c_497_n N_X_c_762_n 0.00987681f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_M1030_s N_X_c_666_n 0.00190439f $X=7.855 $Y=1.485 $X2=0 $Y2=0
cc_457 N_VPWR_M1035_s N_X_c_666_n 0.00336035f $X=8.715 $Y=1.485 $X2=0 $Y2=0
cc_458 N_VPWR_c_510_n N_X_c_666_n 0.014045f $X=7.995 $Y=2.22 $X2=0 $Y2=0
cc_459 N_VPWR_c_512_n N_X_c_666_n 0.0228763f $X=8.855 $Y=2.22 $X2=0 $Y2=0
cc_460 N_VPWR_c_521_n N_X_c_666_n 0.0149478f $X=7.87 $Y=2.717 $X2=0 $Y2=0
cc_461 N_VPWR_c_525_n N_X_c_666_n 0.0161141f $X=8.755 $Y=2.72 $X2=0 $Y2=0
cc_462 N_VPWR_c_497_n N_X_c_666_n 0.020855f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_463 N_X_c_643_n N_VGND_c_877_n 0.0164628f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_464 N_X_c_646_n N_VGND_c_878_n 0.0164628f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_465 N_X_c_648_n N_VGND_c_879_n 0.015936f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_466 N_X_c_648_n N_VGND_c_880_n 0.00226107f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_467 N_X_c_649_n N_VGND_c_880_n 0.0133875f $X=4.99 $Y=0.445 $X2=0 $Y2=0
cc_468 N_X_c_650_n N_VGND_c_880_n 0.00224999f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_469 N_X_c_650_n N_VGND_c_881_n 0.015713f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_470 N_X_c_650_n N_VGND_c_882_n 0.00225184f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_471 N_X_c_651_n N_VGND_c_882_n 0.0128416f $X=5.845 $Y=0.445 $X2=0 $Y2=0
cc_472 N_X_c_652_n N_VGND_c_882_n 0.00239951f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_473 N_X_c_652_n N_VGND_c_883_n 0.0161116f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_474 N_X_c_654_n N_VGND_c_884_n 0.0161116f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_475 X N_VGND_c_885_n 0.0186728f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_476 X N_VGND_c_887_n 0.0243436f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_477 N_X_c_642_n N_VGND_c_890_n 0.0128416f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_478 N_X_c_643_n N_VGND_c_890_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_479 N_X_c_643_n N_VGND_c_892_n 0.00224999f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_480 N_X_c_645_n N_VGND_c_892_n 0.0128416f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_481 N_X_c_646_n N_VGND_c_892_n 0.00224999f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_482 N_X_c_646_n N_VGND_c_894_n 0.00224999f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_483 N_X_c_647_n N_VGND_c_894_n 0.0128416f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_484 N_X_c_648_n N_VGND_c_894_n 0.00224999f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_485 N_X_c_654_n N_VGND_c_896_n 0.00225184f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_486 N_X_c_655_n N_VGND_c_896_n 0.0128416f $X=7.565 $Y=0.445 $X2=0 $Y2=0
cc_487 N_X_c_656_n N_VGND_c_896_n 0.00232492f $X=7.86 $Y=0.82 $X2=0 $Y2=0
cc_488 N_X_c_652_n N_VGND_c_899_n 0.00225184f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_489 N_X_c_653_n N_VGND_c_899_n 0.0128416f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_490 N_X_c_654_n N_VGND_c_899_n 0.00239951f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_491 N_X_c_657_n N_VGND_c_900_n 0.0129027f $X=8.425 $Y=0.445 $X2=0 $Y2=0
cc_492 X N_VGND_c_900_n 0.00498855f $X=7.965 $Y=0.765 $X2=0 $Y2=0
cc_493 N_X_M1002_s N_VGND_c_905_n 0.00268444f $X=2.27 $Y=0.235 $X2=0 $Y2=0
cc_494 N_X_M1004_s N_VGND_c_905_n 0.00234574f $X=3.13 $Y=0.235 $X2=0 $Y2=0
cc_495 N_X_M1008_s N_VGND_c_905_n 0.00234574f $X=3.99 $Y=0.235 $X2=0 $Y2=0
cc_496 N_X_M1017_s N_VGND_c_905_n 0.00230304f $X=4.85 $Y=0.235 $X2=0 $Y2=0
cc_497 N_X_M1020_s N_VGND_c_905_n 0.00234574f $X=5.705 $Y=0.235 $X2=0 $Y2=0
cc_498 N_X_M1029_s N_VGND_c_905_n 0.00234574f $X=6.565 $Y=0.235 $X2=0 $Y2=0
cc_499 N_X_M1032_s N_VGND_c_905_n 0.00234574f $X=7.425 $Y=0.235 $X2=0 $Y2=0
cc_500 N_X_M1036_s N_VGND_c_905_n 0.00234544f $X=8.285 $Y=0.235 $X2=0 $Y2=0
cc_501 N_X_c_642_n N_VGND_c_905_n 0.00979224f $X=2.41 $Y=0.445 $X2=0 $Y2=0
cc_502 N_X_c_643_n N_VGND_c_905_n 0.00829353f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_503 N_X_c_645_n N_VGND_c_905_n 0.00979224f $X=3.27 $Y=0.445 $X2=0 $Y2=0
cc_504 N_X_c_646_n N_VGND_c_905_n 0.00829353f $X=4 $Y=0.82 $X2=0 $Y2=0
cc_505 N_X_c_647_n N_VGND_c_905_n 0.00979224f $X=4.13 $Y=0.445 $X2=0 $Y2=0
cc_506 N_X_c_648_n N_VGND_c_905_n 0.0082634f $X=4.845 $Y=0.82 $X2=0 $Y2=0
cc_507 N_X_c_649_n N_VGND_c_905_n 0.0103326f $X=4.99 $Y=0.445 $X2=0 $Y2=0
cc_508 N_X_c_650_n N_VGND_c_905_n 0.00823851f $X=5.705 $Y=0.82 $X2=0 $Y2=0
cc_509 N_X_c_651_n N_VGND_c_905_n 0.00979224f $X=5.845 $Y=0.445 $X2=0 $Y2=0
cc_510 N_X_c_652_n N_VGND_c_905_n 0.00851943f $X=6.565 $Y=0.82 $X2=0 $Y2=0
cc_511 N_X_c_653_n N_VGND_c_905_n 0.00979224f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_512 N_X_c_654_n N_VGND_c_905_n 0.00851943f $X=7.425 $Y=0.82 $X2=0 $Y2=0
cc_513 N_X_c_655_n N_VGND_c_905_n 0.00979224f $X=7.565 $Y=0.445 $X2=0 $Y2=0
cc_514 N_X_c_656_n N_VGND_c_905_n 0.00379347f $X=7.86 $Y=0.82 $X2=0 $Y2=0
cc_515 N_X_c_657_n N_VGND_c_905_n 0.00981584f $X=8.425 $Y=0.445 $X2=0 $Y2=0
cc_516 X N_VGND_c_905_n 0.0103915f $X=7.965 $Y=0.765 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__clkbuf_16.pex.spice
* Created: Tue Sep  1 18:59:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__CLKBUF_16%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 40
r64 39 40 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.765 $Y2=1.155
r65 38 39 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=1.155
+ $X2=1.335 $Y2=1.155
r66 37 38 45.1103 $w=5.1e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.155
+ $X2=0.905 $Y2=1.155
r67 34 37 21.5061 $w=5.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.475 $Y2=1.155
r68 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r69 29 30 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r70 26 40 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.765 $Y=1.41
+ $X2=1.765 $Y2=1.155
r71 26 28 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.765 $Y=1.41
+ $X2=1.765 $Y2=1.985
r72 22 40 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.765 $Y=0.9
+ $X2=1.765 $Y2=1.155
r73 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.765 $Y=0.9
+ $X2=1.765 $Y2=0.445
r74 19 39 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.335 $Y=1.41
+ $X2=1.335 $Y2=1.155
r75 19 21 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.335 $Y=1.41
+ $X2=1.335 $Y2=1.985
r76 15 39 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.335 $Y=0.9
+ $X2=1.335 $Y2=1.155
r77 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.335 $Y=0.9
+ $X2=1.335 $Y2=0.445
r78 12 38 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.155
r79 12 14 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
r80 8 38 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.155
r81 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r82 5 37 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.155
r83 5 7 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.475 $Y=1.41
+ $X2=0.475 $Y2=1.985
r84 1 37 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.155
r85 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_16%A_110_47# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 133
+ 135 139 143 147 149 153 157 164 167 168
r288 164 165 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=7.505
+ $Y=1.16 $X2=7.505 $Y2=1.16
r289 161 164 235.098 $w=2.48e-07 $l=5.1e-06 $layer=LI1_cond $X=2.405 $Y=1.2
+ $X2=7.505 $Y2=1.2
r290 161 162 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=2.405
+ $Y=1.16 $X2=2.405 $Y2=1.16
r291 159 168 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=1.2 $X2=1.555
+ $Y2=1.2
r292 159 161 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=1.68 $Y=1.2
+ $X2=2.405 $Y2=1.2
r293 155 168 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.325
+ $X2=1.555 $Y2=1.2
r294 155 157 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.555 $Y=1.325
+ $X2=1.555 $Y2=1.92
r295 151 168 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.075
+ $X2=1.555 $Y2=1.2
r296 151 153 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=1.555 $Y=1.075
+ $X2=1.555 $Y2=0.445
r297 150 167 1.3064 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=1.2
+ $X2=0.695 $Y2=1.2
r298 149 168 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.43 $Y=1.2 $X2=1.555
+ $Y2=1.2
r299 149 150 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=1.43 $Y=1.2
+ $X2=0.82 $Y2=1.2
r300 145 167 5.20938 $w=2.47e-07 $l=1.26491e-07 $layer=LI1_cond $X=0.692
+ $Y=1.325 $X2=0.695 $Y2=1.2
r301 145 147 29.8694 $w=2.43e-07 $l=6.35e-07 $layer=LI1_cond $X=0.692 $Y=1.325
+ $X2=0.692 $Y2=1.96
r302 141 167 5.20938 $w=2.47e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=1.2
r303 141 143 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.695 $Y=1.075
+ $X2=0.695 $Y2=0.445
r304 137 139 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.64 $Y=1.325
+ $X2=8.64 $Y2=1.985
r305 133 137 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.64 $Y=1.137
+ $X2=8.64 $Y2=1.325
r306 133 135 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.64 $Y=0.95
+ $X2=8.64 $Y2=0.445
r307 129 131 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.21 $Y=1.325
+ $X2=8.21 $Y2=1.985
r308 125 133 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=8.21 $Y=1.137
+ $X2=8.64 $Y2=1.137
r309 125 129 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=8.21 $Y=1.137
+ $X2=8.21 $Y2=1.325
r310 125 127 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.21 $Y=0.95
+ $X2=8.21 $Y2=0.445
r311 121 123 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.78 $Y=1.325
+ $X2=7.78 $Y2=1.985
r312 117 125 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=8.21 $Y2=1.137
r313 117 121 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=7.78 $Y2=1.325
r314 117 165 40.7846 $w=3.75e-07 $l=2.75e-07 $layer=POLY_cond $X=7.78 $Y=1.137
+ $X2=7.505 $Y2=1.137
r315 117 119 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.78 $Y=0.95
+ $X2=7.78 $Y2=0.445
r316 113 115 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.325
+ $X2=7.35 $Y2=1.985
r317 109 165 22.9877 $w=3.75e-07 $l=1.55e-07 $layer=POLY_cond $X=7.35 $Y=1.137
+ $X2=7.505 $Y2=1.137
r318 109 113 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=7.35 $Y=1.137
+ $X2=7.35 $Y2=1.325
r319 109 111 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.35 $Y=0.95
+ $X2=7.35 $Y2=0.445
r320 105 107 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.92 $Y=1.325
+ $X2=6.92 $Y2=1.985
r321 101 109 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.92 $Y=1.137
+ $X2=7.35 $Y2=1.137
r322 101 105 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.92 $Y=1.137
+ $X2=6.92 $Y2=1.325
r323 101 103 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.92 $Y=0.95
+ $X2=6.92 $Y2=0.445
r324 97 99 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.49 $Y=1.325
+ $X2=6.49 $Y2=1.985
r325 93 101 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.49 $Y=1.137
+ $X2=6.92 $Y2=1.137
r326 93 97 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.49 $Y=1.137
+ $X2=6.49 $Y2=1.325
r327 93 95 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.49 $Y=0.95
+ $X2=6.49 $Y2=0.445
r328 89 91 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.06 $Y=1.325
+ $X2=6.06 $Y2=1.985
r329 85 93 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=6.06 $Y=1.137
+ $X2=6.49 $Y2=1.137
r330 85 89 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.06 $Y=1.137
+ $X2=6.06 $Y2=1.325
r331 85 87 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.06 $Y=0.95
+ $X2=6.06 $Y2=0.445
r332 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r333 77 85 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=5.63 $Y=1.137
+ $X2=6.06 $Y2=1.137
r334 77 81 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=5.63 $Y=1.137
+ $X2=5.63 $Y2=1.325
r335 77 79 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.63 $Y=0.95
+ $X2=5.63 $Y2=0.445
r336 73 75 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.205 $Y=1.325
+ $X2=5.205 $Y2=1.985
r337 69 77 63.0308 $w=3.75e-07 $l=4.25e-07 $layer=POLY_cond $X=5.205 $Y=1.137
+ $X2=5.63 $Y2=1.137
r338 69 73 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=5.205 $Y=1.137
+ $X2=5.205 $Y2=1.325
r339 69 71 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.205 $Y=0.95
+ $X2=5.205 $Y2=0.445
r340 65 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.775 $Y=1.325
+ $X2=4.775 $Y2=1.985
r341 61 69 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.775 $Y=1.137
+ $X2=5.205 $Y2=1.137
r342 61 65 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.775 $Y=1.137
+ $X2=4.775 $Y2=1.325
r343 61 63 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.775 $Y=0.95
+ $X2=4.775 $Y2=0.445
r344 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.345 $Y=1.325
+ $X2=4.345 $Y2=1.985
r345 53 61 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.775 $Y2=1.137
r346 53 57 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=4.345 $Y=1.137
+ $X2=4.345 $Y2=1.325
r347 53 55 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.345 $Y=0.95
+ $X2=4.345 $Y2=0.445
r348 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.915 $Y=1.325
+ $X2=3.915 $Y2=1.985
r349 45 53 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=4.345 $Y2=1.137
r350 45 49 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.915 $Y=1.137
+ $X2=3.915 $Y2=1.325
r351 45 47 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.915 $Y=0.95
+ $X2=3.915 $Y2=0.445
r352 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.325
+ $X2=3.485 $Y2=1.985
r353 37 45 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.915 $Y2=1.137
r354 37 41 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.485 $Y=1.137
+ $X2=3.485 $Y2=1.325
r355 37 39 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.485 $Y=0.95
+ $X2=3.485 $Y2=0.445
r356 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.985
r357 29 37 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.485 $Y2=1.137
r358 29 33 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.055 $Y=1.137
+ $X2=3.055 $Y2=1.325
r359 29 31 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.055 $Y=0.95
+ $X2=3.055 $Y2=0.445
r360 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=1.325
+ $X2=2.625 $Y2=1.985
r361 21 29 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=3.055 $Y2=1.137
r362 21 25 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.625 $Y2=1.325
r363 21 162 32.6277 $w=3.75e-07 $l=2.2e-07 $layer=POLY_cond $X=2.625 $Y=1.137
+ $X2=2.405 $Y2=1.137
r364 21 23 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.625 $Y=0.95
+ $X2=2.625 $Y2=0.445
r365 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.195 $Y=1.325
+ $X2=2.195 $Y2=1.985
r366 13 162 31.1446 $w=3.75e-07 $l=2.1e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.405 $Y2=1.137
r367 13 17 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=2.195 $Y=1.137
+ $X2=2.195 $Y2=1.325
r368 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.195 $Y=0.95
+ $X2=2.195 $Y2=0.445
r369 4 157 300 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.485 $X2=1.55 $Y2=1.92
r370 3 147 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.485 $X2=0.69 $Y2=1.96
r371 2 153 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
r372 1 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 52 56 58 62 64 68 72 76 78 80 83 84 86 87 89 90 91 92 94 95 96 98 116 125
+ 133 136 139 142 146
c145 11 0 4.2343e-20 $X=8.715 $Y=1.485
r146 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r147 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r148 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r149 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r150 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r151 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r152 128 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r153 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r154 125 145 4.10457 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.755 $Y=2.72
+ $X2=8.977 $Y2=2.72
r155 125 127 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.755 $Y=2.72
+ $X2=8.51 $Y2=2.72
r156 124 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r157 124 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r158 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r159 121 142 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=7.255 $Y=2.717
+ $X2=7.132 $Y2=2.717
r160 121 123 21.2312 $w=1.73e-07 $l=3.35e-07 $layer=LI1_cond $X=7.255 $Y=2.717
+ $X2=7.59 $Y2=2.717
r161 120 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r162 120 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r163 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 117 139 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=6.395 $Y=2.717
+ $X2=6.272 $Y2=2.717
r165 117 119 17.4286 $w=1.73e-07 $l=2.75e-07 $layer=LI1_cond $X=6.395 $Y=2.717
+ $X2=6.67 $Y2=2.717
r166 116 142 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=7.01 $Y=2.717
+ $X2=7.132 $Y2=2.717
r167 116 119 21.5481 $w=1.73e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.717
+ $X2=6.67 $Y2=2.717
r168 115 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r169 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r170 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r171 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r172 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r173 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r174 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r175 106 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r176 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r177 103 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.12 $Y2=2.72
r178 103 105 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.61 $Y2=2.72
r179 102 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r180 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r181 99 130 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r182 99 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.69 $Y2=2.72
r183 98 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=1.12 $Y2=2.72
r184 98 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 96 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r186 96 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r187 94 123 17.7455 $w=1.73e-07 $l=2.8e-07 $layer=LI1_cond $X=7.87 $Y=2.717
+ $X2=7.59 $Y2=2.717
r188 94 95 7.05609 $w=1.72e-07 $l=1.27e-07 $layer=LI1_cond $X=7.87 $Y=2.717
+ $X2=7.997 $Y2=2.717
r189 93 127 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.125 $Y=2.72
+ $X2=8.51 $Y2=2.72
r190 93 95 7.05609 $w=1.72e-07 $l=1.29491e-07 $layer=LI1_cond $X=8.125 $Y=2.72
+ $X2=7.997 $Y2=2.717
r191 91 114 3.8026 $w=1.73e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=2.717
+ $X2=4.37 $Y2=2.717
r192 91 92 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.43 $Y=2.717
+ $X2=4.56 $Y2=2.717
r193 89 111 7.60519 $w=1.73e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=2.717
+ $X2=3.45 $Y2=2.717
r194 89 90 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=2.717
+ $X2=3.7 $Y2=2.717
r195 88 114 34.2234 $w=1.73e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=2.717
+ $X2=4.37 $Y2=2.717
r196 88 90 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=2.717
+ $X2=3.7 $Y2=2.717
r197 86 108 11.4078 $w=1.73e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=2.717
+ $X2=2.53 $Y2=2.717
r198 86 87 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=2.717
+ $X2=2.84 $Y2=2.717
r199 85 111 30.4208 $w=1.73e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=2.717
+ $X2=3.45 $Y2=2.717
r200 85 87 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=2.717
+ $X2=2.84 $Y2=2.717
r201 83 105 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.61 $Y2=2.72
r202 83 84 7.16073 $w=1.72e-07 $l=1.31491e-07 $layer=LI1_cond $X=1.85 $Y=2.72
+ $X2=1.98 $Y2=2.717
r203 82 108 26.6182 $w=1.73e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=2.717
+ $X2=2.53 $Y2=2.717
r204 82 84 7.16073 $w=1.72e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=2.717
+ $X2=1.98 $Y2=2.717
r205 78 145 3.18012 $w=2.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=8.89 $Y=2.635
+ $X2=8.977 $Y2=2.72
r206 78 80 17.7135 $w=2.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.89 $Y=2.635
+ $X2=8.89 $Y2=2.22
r207 74 95 0.0190999 $w=2.55e-07 $l=8.7e-08 $layer=LI1_cond $X=7.997 $Y=2.63
+ $X2=7.997 $Y2=2.717
r208 74 76 18.5295 $w=2.53e-07 $l=4.1e-07 $layer=LI1_cond $X=7.997 $Y=2.63
+ $X2=7.997 $Y2=2.22
r209 70 142 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=7.132 $Y=2.63
+ $X2=7.132 $Y2=2.717
r210 70 72 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=7.132 $Y=2.63
+ $X2=7.132 $Y2=2.22
r211 66 139 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=6.272 $Y=2.63
+ $X2=6.272 $Y2=2.717
r212 66 68 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=6.272 $Y=2.63
+ $X2=6.272 $Y2=2.22
r213 65 136 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=5.535 $Y=2.717
+ $X2=5.412 $Y2=2.717
r214 64 139 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=6.15 $Y=2.717
+ $X2=6.272 $Y2=2.717
r215 64 65 38.9766 $w=1.73e-07 $l=6.15e-07 $layer=LI1_cond $X=6.15 $Y=2.717
+ $X2=5.535 $Y2=2.717
r216 60 136 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=5.412 $Y=2.63
+ $X2=5.412 $Y2=2.717
r217 60 62 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=5.412 $Y=2.63
+ $X2=5.412 $Y2=2.22
r218 59 92 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.69 $Y=2.717
+ $X2=4.56 $Y2=2.717
r219 58 136 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=5.29 $Y=2.717
+ $X2=5.412 $Y2=2.717
r220 58 59 38.026 $w=1.73e-07 $l=6e-07 $layer=LI1_cond $X=5.29 $Y=2.717 $X2=4.69
+ $Y2=2.717
r221 54 92 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=4.56 $Y=2.63
+ $X2=4.56 $Y2=2.717
r222 54 56 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=4.56 $Y=2.63
+ $X2=4.56 $Y2=2.22
r223 50 90 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=3.7 $Y=2.63
+ $X2=3.7 $Y2=2.717
r224 50 52 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=3.7 $Y=2.63 $X2=3.7
+ $Y2=2.22
r225 46 87 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=2.84 $Y=2.63
+ $X2=2.84 $Y2=2.717
r226 46 48 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=2.84 $Y=2.63
+ $X2=2.84 $Y2=2.22
r227 42 84 0.0838798 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=1.98 $Y=2.63
+ $X2=1.98 $Y2=2.717
r228 42 44 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=1.98 $Y=2.63
+ $X2=1.98 $Y2=2
r229 38 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r230 38 40 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2
r231 34 130 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.195 $Y2=2.72
r232 34 36 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=2
r233 11 80 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.485 $X2=8.855 $Y2=2.22
r234 10 76 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.485 $X2=7.995 $Y2=2.22
r235 9 72 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=6.995
+ $Y=1.485 $X2=7.135 $Y2=2.22
r236 8 68 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=6.135
+ $Y=1.485 $X2=6.275 $Y2=2.22
r237 7 62 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.485 $X2=5.42 $Y2=2.22
r238 6 56 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.485 $X2=4.56 $Y2=2.22
r239 5 52 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.7 $Y2=2.22
r240 4 48 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.485 $X2=2.84 $Y2=2.22
r241 3 44 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=1.485 $X2=1.98 $Y2=2
r242 2 40 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.485 $X2=1.12 $Y2=2
r243 1 36 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 56 57 61 65 67 71 75 77 81 85 87 91 95 97 101 105 107 111 115 119 124
+ 125 127 128 130 131 133 134 136 137 139 140 141 142 143 168 173
c231 141 0 1.18325e-19 $X=8.51 $Y=0.85
r232 171 173 0.603562 $w=1.516e-06 $l=7.5e-08 $layer=LI1_cond $X=8.225 $Y=1.615
+ $X2=8.225 $Y2=1.69
r233 158 168 0.966712 $w=1.516e-06 $l=2.33846e-07 $layer=LI1_cond $X=8.442
+ $Y=1.495 $X2=8.225 $Y2=1.53
r234 143 171 0.48285 $w=1.516e-06 $l=6e-08 $layer=LI1_cond $X=8.225 $Y=1.555
+ $X2=8.225 $Y2=1.615
r235 143 168 0.201187 $w=1.516e-06 $l=2.5e-08 $layer=LI1_cond $X=8.225 $Y=1.555
+ $X2=8.225 $Y2=1.53
r236 143 158 0.261803 $w=1.163e-06 $l=2.5e-08 $layer=LI1_cond $X=8.442 $Y=1.47
+ $X2=8.442 $Y2=1.495
r237 142 143 2.93219 $w=1.163e-06 $l=2.8e-07 $layer=LI1_cond $X=8.442 $Y=1.19
+ $X2=8.442 $Y2=1.47
r238 141 157 1.4003 $w=7.12e-07 $l=8.5e-08 $layer=LI1_cond $X=8.442 $Y=0.82
+ $X2=8.442 $Y2=0.905
r239 141 142 2.82747 $w=1.163e-06 $l=2.7e-07 $layer=LI1_cond $X=8.442 $Y=0.92
+ $X2=8.442 $Y2=1.19
r240 141 157 0.157082 $w=1.163e-06 $l=1.5e-08 $layer=LI1_cond $X=8.442 $Y=0.92
+ $X2=8.442 $Y2=0.905
r241 117 141 1.4003 $w=7.12e-07 $l=9.31128e-08 $layer=LI1_cond $X=8.425 $Y=0.735
+ $X2=8.442 $Y2=0.82
r242 117 119 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=8.425 $Y=0.735
+ $X2=8.425 $Y2=0.445
r243 116 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.685 $Y=0.82
+ $X2=7.555 $Y2=0.82
r244 115 141 6.76561 $w=1.7e-07 $l=5.82e-07 $layer=LI1_cond $X=7.86 $Y=0.82
+ $X2=8.442 $Y2=0.82
r245 115 116 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.86 $Y=0.82
+ $X2=7.685 $Y2=0.82
r246 109 140 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0.735
+ $X2=7.555 $Y2=0.82
r247 109 111 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=7.555 $Y=0.735
+ $X2=7.555 $Y2=0.445
r248 108 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=1.615
+ $X2=6.695 $Y2=1.615
r249 107 171 12.2163 $w=2.4e-07 $l=8e-07 $layer=LI1_cond $X=7.425 $Y=1.615
+ $X2=8.225 $Y2=1.615
r250 107 108 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=7.425 $Y=1.615
+ $X2=6.825 $Y2=1.615
r251 106 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=0.82
+ $X2=6.695 $Y2=0.82
r252 105 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.425 $Y=0.82
+ $X2=7.555 $Y2=0.82
r253 105 106 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.425 $Y=0.82
+ $X2=6.825 $Y2=0.82
r254 99 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=0.735
+ $X2=6.695 $Y2=0.82
r255 99 101 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=6.695 $Y=0.735
+ $X2=6.695 $Y2=0.445
r256 98 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.965 $Y=1.615
+ $X2=5.835 $Y2=1.615
r257 97 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.565 $Y=1.615
+ $X2=6.695 $Y2=1.615
r258 97 98 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=6.565 $Y=1.615
+ $X2=5.965 $Y2=1.615
r259 96 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.965 $Y=0.82
+ $X2=5.835 $Y2=0.82
r260 95 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.565 $Y=0.82
+ $X2=6.695 $Y2=0.82
r261 95 96 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.565 $Y=0.82
+ $X2=5.965 $Y2=0.82
r262 89 134 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0.735
+ $X2=5.835 $Y2=0.82
r263 89 91 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=5.835 $Y=0.735
+ $X2=5.835 $Y2=0.445
r264 88 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.12 $Y=1.615
+ $X2=4.99 $Y2=1.615
r265 87 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.705 $Y=1.615
+ $X2=5.835 $Y2=1.615
r266 87 88 28.0908 $w=2.38e-07 $l=5.85e-07 $layer=LI1_cond $X=5.705 $Y=1.615
+ $X2=5.12 $Y2=1.615
r267 86 131 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.12 $Y=0.82
+ $X2=4.982 $Y2=0.82
r268 85 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.705 $Y=0.82
+ $X2=5.835 $Y2=0.82
r269 85 86 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=5.705 $Y=0.82
+ $X2=5.12 $Y2=0.82
r270 79 131 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.982 $Y=0.735
+ $X2=4.982 $Y2=0.82
r271 79 81 12.153 $w=2.73e-07 $l=2.9e-07 $layer=LI1_cond $X=4.982 $Y=0.735
+ $X2=4.982 $Y2=0.445
r272 78 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=1.615
+ $X2=4.13 $Y2=1.615
r273 77 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.86 $Y=1.615
+ $X2=4.99 $Y2=1.615
r274 77 78 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=4.86 $Y=1.615
+ $X2=4.26 $Y2=1.615
r275 76 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=0.82
+ $X2=4.13 $Y2=0.82
r276 75 131 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.845 $Y=0.82
+ $X2=4.982 $Y2=0.82
r277 75 76 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.845 $Y=0.82
+ $X2=4.26 $Y2=0.82
r278 69 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.82
r279 69 71 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r280 68 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.615
+ $X2=3.27 $Y2=1.615
r281 67 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=1.615 $X2=4.13
+ $Y2=1.615
r282 67 68 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=1.615 $X2=3.4
+ $Y2=1.615
r283 66 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.82
+ $X2=3.27 $Y2=0.82
r284 65 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=0.82 $X2=4.13
+ $Y2=0.82
r285 65 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=0.82 $X2=3.4
+ $Y2=0.82
r286 59 125 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.82
r287 59 61 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r288 58 124 3.55196 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.615
+ $X2=2.41 $Y2=1.615
r289 57 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=3.27 $Y2=1.615
r290 57 58 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.615
+ $X2=2.54 $Y2=1.615
r291 55 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.82
+ $X2=3.27 $Y2=0.82
r292 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.82 $X2=2.54
+ $Y2=0.82
r293 49 56 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.54 $Y2=0.82
r294 49 51 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r295 16 173 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=8.285
+ $Y=1.485 $X2=8.425 $Y2=1.69
r296 15 173 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=7.425
+ $Y=1.485 $X2=7.565 $Y2=1.69
r297 14 139 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=6.565
+ $Y=1.485 $X2=6.705 $Y2=1.69
r298 13 136 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=5.705
+ $Y=1.485 $X2=5.845 $Y2=1.69
r299 12 133 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=4.85
+ $Y=1.485 $X2=4.99 $Y2=1.69
r300 11 130 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.485 $X2=4.13 $Y2=1.69
r301 10 127 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.485 $X2=3.27 $Y2=1.69
r302 9 124 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.485 $X2=2.41 $Y2=1.69
r303 8 119 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.285
+ $Y=0.235 $X2=8.425 $Y2=0.445
r304 7 111 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.565 $Y2=0.445
r305 6 101 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.565
+ $Y=0.235 $X2=6.705 $Y2=0.445
r306 5 91 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.845 $Y2=0.445
r307 4 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.235 $X2=4.99 $Y2=0.445
r308 3 71 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r309 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r310 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__CLKBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 52 56 58 62 64 68 72 76 78 80 83 84 86 87 89 90 91 92 94 95 96 98 116 125
+ 133 136 139 142 146
c160 94 0 7.59816e-20 $X=7.865 $Y=0
r161 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r162 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r163 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r164 137 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r165 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r166 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r167 128 146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r168 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r169 125 145 4.35621 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.962 $Y2=0
r170 125 127 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.725 $Y=0
+ $X2=8.51 $Y2=0
r171 124 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r172 124 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r173 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r174 121 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.13 $Y2=0
r175 121 123 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.59 $Y2=0
r176 120 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r177 120 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r178 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r179 117 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.395 $Y=0
+ $X2=6.27 $Y2=0
r180 117 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.395 $Y=0
+ $X2=6.67 $Y2=0
r181 116 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.13 $Y2=0
r182 116 119 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.67 $Y2=0
r183 115 137 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r184 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r185 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r186 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r187 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r188 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r189 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r190 106 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r191 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r192 103 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r193 103 105 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=0
+ $X2=1.61 $Y2=0
r194 102 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r195 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r196 99 130 4.57719 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0
+ $X2=0.195 $Y2=0
r197 99 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r198 98 133 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r199 98 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.69
+ $Y2=0
r200 96 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r201 96 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r202 94 123 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.865 $Y=0
+ $X2=7.59 $Y2=0
r203 94 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.865 $Y=0 $X2=7.995
+ $Y2=0
r204 93 127 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.125 $Y=0
+ $X2=8.51 $Y2=0
r205 93 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.125 $Y=0 $X2=7.995
+ $Y2=0
r206 91 114 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.37
+ $Y2=0
r207 91 92 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.552
+ $Y2=0
r208 89 111 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r209 89 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r210 88 114 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.37
+ $Y2=0
r211 88 90 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r212 86 108 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.53
+ $Y2=0
r213 86 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r214 85 111 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=3.45
+ $Y2=0
r215 85 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r216 83 105 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.61
+ $Y2=0
r217 83 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r218 82 108 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.53
+ $Y2=0
r219 82 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r220 78 145 3.16147 $w=3e-07 $l=1.22327e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.962 $Y2=0
r221 78 80 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0.4
r222 74 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=0.085
+ $X2=7.995 $Y2=0
r223 74 76 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.995 $Y=0.085
+ $X2=7.995 $Y2=0.4
r224 70 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0
r225 70 72 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0.4
r226 66 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0
r227 66 68 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.27 $Y=0.085
+ $X2=6.27 $Y2=0.4
r228 65 136 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=5.535 $Y=0
+ $X2=5.412 $Y2=0
r229 64 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=6.27 $Y2=0
r230 64 65 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.145 $Y=0
+ $X2=5.535 $Y2=0
r231 60 136 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.412 $Y=0.085
+ $X2=5.412 $Y2=0
r232 60 62 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=5.412 $Y=0.085
+ $X2=5.412 $Y2=0.4
r233 59 92 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=4.552 $Y2=0
r234 58 136 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.412 $Y2=0
r235 58 59 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.29 $Y=0 $X2=4.675
+ $Y2=0
r236 54 92 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.552 $Y2=0
r237 54 56 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=4.552 $Y=0.085
+ $X2=4.552 $Y2=0.4
r238 50 90 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r239 50 52 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r240 46 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r241 46 48 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r242 42 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r243 42 44 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.445
r244 38 133 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r245 38 40 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r246 34 130 2.98104 $w=3.05e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.195 $Y2=0
r247 34 36 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.38
r248 11 80 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.715
+ $Y=0.235 $X2=8.855 $Y2=0.4
r249 10 76 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.235 $X2=7.995 $Y2=0.4
r250 9 72 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=0.235 $X2=7.135 $Y2=0.4
r251 8 68 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.135
+ $Y=0.235 $X2=6.275 $Y2=0.4
r252 7 62 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.28
+ $Y=0.235 $X2=5.42 $Y2=0.4
r253 6 56 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.56 $Y2=0.4
r254 5 52 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r255 4 48 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r256 3 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.445
r257 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r258 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__or4b_1.pex.spice
* Created: Thu Aug 27 14:44:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR4B_1%D_N 3 7 9 10 17
r26 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r27 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r28 9 10 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.255 $Y=0.85
+ $X2=0.255 $Y2=1.16
r29 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r30 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r31 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r32 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%A_109_53# 1 2 9 13 17 21 27 32
r40 28 32 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.165 $Y=1.16
+ $X2=1.41 $Y2=1.16
r41 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.16 $X2=1.165 $Y2=1.16
r42 25 27 15.6453 $w=3.28e-07 $l=4.48e-07 $layer=LI1_cond $X=0.717 $Y=1.16
+ $X2=1.165 $Y2=1.16
r43 23 25 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=0.715 $Y=1.16
+ $X2=0.717 $Y2=1.16
r44 19 23 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=1.325
+ $X2=0.715 $Y2=1.16
r45 19 21 18.9673 $w=2.38e-07 $l=3.95e-07 $layer=LI1_cond $X=0.715 $Y=1.325
+ $X2=0.715 $Y2=1.72
r46 15 25 2.50173 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=0.717 $Y=0.995
+ $X2=0.717 $Y2=1.16
r47 15 17 23.2841 $w=2.43e-07 $l=4.95e-07 $layer=LI1_cond $X=0.717 $Y=0.995
+ $X2=0.717 $Y2=0.5
r48 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.16
r49 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.41 $Y=1.325
+ $X2=1.41 $Y2=1.695
r50 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.16
r51 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.475
r52 2 21 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.72
r53 1 17 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.265 $X2=0.68 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%C 3 7 9 11 18
r37 18 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=1.83 $Y2=1.325
r38 18 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.16
+ $X2=1.83 $Y2=0.995
r39 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.16 $X2=1.83 $Y2=1.16
r40 11 19 4.62998 $w=6.18e-07 $l=2.4e-07 $layer=LI1_cond $X=2.07 $Y=1.305
+ $X2=1.83 $Y2=1.305
r41 9 19 4.24415 $w=6.18e-07 $l=2.2e-07 $layer=LI1_cond $X=1.61 $Y=1.305
+ $X2=1.83 $Y2=1.305
r42 7 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.885 $Y=1.695
+ $X2=1.885 $Y2=1.325
r43 3 20 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.865 $Y=0.475
+ $X2=1.865 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%B 2 4 7 8 9 10 11 12 13 20
r40 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=2.28 $X2=2.295 $Y2=2.28
r41 13 20 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.07 $Y=2.27
+ $X2=2.295 $Y2=2.27
r42 12 13 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=1.61 $Y=2.27
+ $X2=2.07 $Y2=2.27
r43 11 12 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=2.27
+ $X2=1.61 $Y2=2.27
r44 10 11 18.0814 $w=2.88e-07 $l=4.55e-07 $layer=LI1_cond $X=0.695 $Y=2.27
+ $X2=1.15 $Y2=2.27
r45 8 9 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=2.267 $Y=0.76
+ $X2=2.267 $Y2=0.91
r46 7 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.285 $Y=0.475
+ $X2=2.285 $Y2=0.76
r47 4 9 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.25 $Y=1.695
+ $X2=2.25 $Y2=0.91
r48 2 19 34.1791 $w=3.28e-07 $l=1.55885e-07 $layer=POLY_cond $X=2.25 $Y=2.145
+ $X2=2.295 $Y2=2.28
r49 2 4 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.25 $Y=2.145 $X2=2.25
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%A 3 7 9 12 13
r42 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=1.325
r43 12 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.69 $Y2=0.995
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.16 $X2=2.69 $Y2=1.16
r45 9 13 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=1.16 $X2=2.69
+ $Y2=1.16
r46 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.705 $Y=1.695
+ $X2=2.705 $Y2=1.325
r47 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.705 $Y=0.475
+ $X2=2.705 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%A_215_297# 1 2 3 12 15 17 21 23 24 27 29 31
+ 36 38 42 43 48 49 50 53
c98 48 0 1.14153e-19 $X=3.17 $Y=1.16
c99 36 0 1.06604e-19 $X=3.065 $Y=1.495
r100 49 54 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.17 $Y2=1.325
r101 49 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.16
+ $X2=3.17 $Y2=0.995
r102 48 51 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.117 $Y=1.16
+ $X2=3.117 $Y2=1.325
r103 48 50 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.117 $Y=1.16
+ $X2=3.117 $Y2=0.995
r104 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.16 $X2=3.17 $Y2=1.16
r105 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.575 $Y=1.58
+ $X2=2.575 $Y2=1.87
r106 38 40 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=1.19 $Y=1.685
+ $X2=1.19 $Y2=1.87
r107 36 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.065 $Y=1.495
+ $X2=3.065 $Y2=1.325
r108 33 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.065 $Y=0.825
+ $X2=3.065 $Y2=0.995
r109 32 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.58
+ $X2=2.575 $Y2=1.58
r110 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.98 $Y=1.58
+ $X2=3.065 $Y2=1.495
r111 31 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.98 $Y=1.58
+ $X2=2.66 $Y2=1.58
r112 30 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.74
+ $X2=2.495 $Y2=0.74
r113 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.98 $Y=0.74
+ $X2=3.065 $Y2=0.825
r114 29 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.98 $Y=0.74 $X2=2.58
+ $Y2=0.74
r115 25 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.655
+ $X2=2.495 $Y2=0.74
r116 25 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.495 $Y=0.655
+ $X2=2.495 $Y2=0.47
r117 23 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.74
+ $X2=2.495 $Y2=0.74
r118 23 24 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.41 $Y=0.74
+ $X2=1.735 $Y2=0.74
r119 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=0.655
+ $X2=1.735 $Y2=0.74
r120 19 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.65 $Y=0.655
+ $X2=1.65 $Y2=0.47
r121 18 40 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.35 $Y=1.87
+ $X2=1.19 $Y2=1.87
r122 17 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=1.87
+ $X2=2.575 $Y2=1.87
r123 17 18 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.49 $Y=1.87
+ $X2=1.35 $Y2=1.87
r124 15 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.195 $Y=1.985
+ $X2=3.195 $Y2=1.325
r125 12 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.195 $Y=0.56
+ $X2=3.195 $Y2=0.995
r126 3 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.2 $Y2=1.685
r127 2 27 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.265 $X2=2.495 $Y2=0.47
r128 1 21 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.265 $X2=1.65 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%VPWR 1 2 7 9 13 15 17 27 28 34
c37 2 0 1.06604e-19 $X=2.78 $Y=1.485
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r41 25 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.11 $Y=2.72 $X2=2.97
+ $Y2=2.72
r42 25 27 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 21 24 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 20 23 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 18 31 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r49 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 17 34 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.83 $Y=2.72 $X2=2.97
+ $Y2=2.72
r51 17 23 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.83 $Y=2.72 $X2=2.53
+ $Y2=2.72
r52 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r53 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 11 34 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2.72
r55 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.97 $Y=2.635
+ $X2=2.97 $Y2=2
r56 7 31 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.212 $Y2=2.72
r57 7 9 31.0143 $w=3.38e-07 $l=9.15e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=1.72
r58 2 13 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=1.485 $X2=2.98 $Y2=2
r59 1 9 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.72
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%X 1 2 12 14 15 16
r18 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=3.457 $Y=1.632
+ $X2=3.457 $Y2=1.845
r19 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=3.457 $Y=1.632
+ $X2=3.457 $Y2=1.495
r20 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=3.405 $Y=0.587
+ $X2=3.51 $Y2=0.587
r21 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.51 $Y=0.76 $X2=3.51
+ $Y2=0.587
r22 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.51 $Y=0.76
+ $X2=3.51 $Y2=1.495
r23 2 16 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=1.485 $X2=3.405 $Y2=1.845
r24 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.235 $X2=3.405 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR4B_1%VGND 1 2 3 4 13 15 19 23 27 29 31 36 41 48 49
+ 55 58 61
r64 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r65 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r66 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r67 49 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r68 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r69 46 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=2.94
+ $Y2=0
r70 46 48 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.45
+ $Y2=0
r71 45 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r72 45 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r73 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r74 42 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.075
+ $Y2=0
r75 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.53
+ $Y2=0
r76 41 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.94
+ $Y2=0
r77 41 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.53
+ $Y2=0
r78 40 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r79 40 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r80 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r81 37 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.2
+ $Y2=0
r82 37 39 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.61
+ $Y2=0
r83 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=2.075
+ $Y2=0
r84 36 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=1.61
+ $Y2=0
r85 35 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r86 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r87 32 52 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r88 32 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r89 31 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r90 31 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.69
+ $Y2=0
r91 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r92 29 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r93 25 61 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r94 25 27 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.4
r95 21 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r96 21 23 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.4
r97 17 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085 $X2=1.2
+ $Y2=0
r98 17 19 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.5
r99 13 52 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.212 $Y2=0
r100 13 15 14.0666 $w=3.38e-07 $l=4.15e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.5
r101 4 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.265 $X2=2.965 $Y2=0.4
r102 3 23 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.265 $X2=2.075 $Y2=0.4
r103 2 19 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.265 $X2=1.2 $Y2=0.5
r104 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends


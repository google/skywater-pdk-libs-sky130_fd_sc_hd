* File: sky130_fd_sc_hd__o31a_1.spice.pex
* Created: Thu Aug 27 14:39:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O31A_1%A_103_199# 1 2 7 9 12 16 17 19 20 22 23 24 25
+ 26 27 30 34
c82 30 0 1.67937e-19 $X=3.05 $Y=1.495
c83 17 0 1.97172e-19 $X=0.65 $Y=1.16
r84 34 36 16.7792 $w=4.88e-07 $l=4.65e-07 $layer=LI1_cond $X=2.89 $Y=0.36
+ $X2=2.89 $Y2=0.825
r85 30 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=1.495
+ $X2=3.05 $Y2=0.825
r86 28 32 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.615 $Y=1.58
+ $X2=2.49 $Y2=1.58
r87 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.965 $Y=1.58
+ $X2=3.05 $Y2=1.495
r88 27 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.965 $Y=1.58
+ $X2=2.615 $Y2=1.58
r89 25 32 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=1.665
+ $X2=2.49 $Y2=1.58
r90 25 26 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=2.49 $Y=1.665
+ $X2=2.49 $Y2=2.295
r91 23 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.365 $Y=2.38
+ $X2=2.49 $Y2=2.295
r92 23 24 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.365 $Y=2.38
+ $X2=1.355 $Y2=2.38
r93 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.27 $Y=2.295
+ $X2=1.355 $Y2=2.38
r94 21 22 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.27 $Y=1.615
+ $X2=1.27 $Y2=2.295
r95 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.185 $Y=1.53
+ $X2=1.27 $Y2=1.615
r96 19 20 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.185 $Y=1.53
+ $X2=0.735 $Y2=1.53
r97 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.65
+ $Y=1.16 $X2=0.65 $Y2=1.16
r98 14 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.65 $Y=1.445
+ $X2=0.735 $Y2=1.53
r99 14 16 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.65 $Y=1.445
+ $X2=0.65 $Y2=1.16
r100 10 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.325
+ $X2=0.65 $Y2=1.16
r101 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.65 $Y=1.325
+ $X2=0.65 $Y2=1.985
r102 7 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=0.995
+ $X2=0.65 $Y2=1.16
r103 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.65 $Y=0.995
+ $X2=0.65 $Y2=0.56
r104 2 32 300 $w=1.7e-07 $l=3.62077e-07 $layer=licon1_PDIFF $count=2 $X=2.165
+ $Y=1.485 $X2=2.45 $Y2=1.66
r105 1 34 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=2.645
+ $Y=0.235 $X2=2.81 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%A1 3 6 8 11 13
r33 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.16
+ $X2=1.13 $Y2=1.325
r34 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.16
+ $X2=1.13 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.16 $X2=1.13 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.19 $Y=1.985
+ $X2=1.19 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.19 $Y=0.56 $X2=1.19
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%A2 1 3 6 8 9 10 15
c36 15 0 1.90303e-19 $X=1.61 $Y=1.16
r37 9 10 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.625 $Y=1.53
+ $X2=1.625 $Y2=1.87
r38 9 26 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.625 $Y=1.53
+ $X2=1.625 $Y2=1.325
r39 8 26 8.18414 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.602 $Y=1.16
+ $X2=1.602 $Y2=1.325
r40 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r41 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.325
+ $X2=1.61 $Y2=1.16
r42 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.61 $Y=1.325 $X2=1.61
+ $Y2=1.985
r43 1 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=0.995
+ $X2=1.61 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.61 $Y=0.995 $X2=1.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%A3 1 3 6 8 11
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.16 $X2=2.09 $Y2=1.16
r36 4 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.325
+ $X2=2.09 $Y2=1.16
r37 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.09 $Y=1.325 $X2=2.09
+ $Y2=1.985
r38 1 11 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=0.995
+ $X2=2.09 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.09 $Y=0.995 $X2=2.09
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%B1 3 6 8 11 13
r33 11 14 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.587 $Y=1.16
+ $X2=2.587 $Y2=1.325
r34 11 13 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=2.587 $Y=1.16
+ $X2=2.587 $Y2=0.995
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.57
+ $Y=1.16 $X2=2.57 $Y2=1.16
r36 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.665 $Y=1.985
+ $X2=2.665 $Y2=1.325
r37 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.56 $X2=2.57
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%X 1 2 7 8 9 10 11 12 24 32 39
c16 39 0 1.76926e-19 $X=0.23 $Y=1.87
r17 39 40 1.93707 $w=4.38e-07 $l=3.5e-08 $layer=LI1_cond $X=0.305 $Y=1.87
+ $X2=0.305 $Y2=1.835
r18 24 37 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=0.85
+ $X2=0.24 $Y2=0.825
r19 12 43 6.54797 $w=4.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.305 $Y=2.21
+ $X2=0.305 $Y2=1.96
r20 11 43 1.70247 $w=4.38e-07 $l=6.5e-08 $layer=LI1_cond $X=0.305 $Y=1.895
+ $X2=0.305 $Y2=1.96
r21 11 39 0.654797 $w=4.38e-07 $l=2.5e-08 $layer=LI1_cond $X=0.305 $Y=1.895
+ $X2=0.305 $Y2=1.87
r22 11 40 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=1.81
+ $X2=0.24 $Y2=1.835
r23 10 11 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=1.53
+ $X2=0.24 $Y2=1.81
r24 9 10 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=1.19 $X2=0.24
+ $Y2=1.53
r25 8 37 1.80611 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=0.305 $Y=0.795
+ $X2=0.305 $Y2=0.825
r26 8 9 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=0.88 $X2=0.24
+ $Y2=1.19
r27 8 24 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.88 $X2=0.24
+ $Y2=0.85
r28 7 8 7.46469 $w=4.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.305 $Y=0.51
+ $X2=0.305 $Y2=0.795
r29 7 32 3.92878 $w=4.38e-07 $l=1.5e-07 $layer=LI1_cond $X=0.305 $Y=0.51
+ $X2=0.305 $Y2=0.36
r30 2 43 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=1.485 $X2=0.36 $Y2=1.96
r31 1 32 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.235 $X2=0.36 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%VPWR 1 2 9 11 13 16 17 18 24 33
c38 9 0 2.02454e-20 $X=0.92 $Y=1.96
c39 2 0 1.67937e-19 $X=2.74 $Y=1.485
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r42 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 24 32 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.007 $Y2=2.72
r47 24 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 22 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 16 21 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.7 $Y=2.72 $X2=0.69
+ $Y2=2.72
r52 16 17 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=0.7 $Y=2.72
+ $X2=0.857 $Y2=2.72
r53 15 26 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 15 17 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.857 $Y2=2.72
r55 11 32 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=3.007 $Y2=2.72
r56 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=1.96
r57 7 17 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.857 $Y=2.635
+ $X2=0.857 $Y2=2.72
r58 7 9 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=0.857 $Y=2.635
+ $X2=0.857 $Y2=1.96
r59 2 13 300 $w=1.7e-07 $l=5.74565e-07 $layer=licon1_PDIFF $count=2 $X=2.74
+ $Y=1.485 $X2=2.96 $Y2=1.96
r60 1 9 300 $w=1.7e-07 $l=5.64137e-07 $layer=licon1_PDIFF $count=2 $X=0.725
+ $Y=1.485 $X2=0.92 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%VGND 1 2 9 12 13 14 20 26 27 31
r47 31 34 9.87808 $w=4.18e-07 $l=3.6e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.865
+ $Y2=0.36
r48 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 27 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r50 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r51 24 31 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.865
+ $Y2=0
r52 24 26 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.99
+ $Y2=0
r53 23 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r54 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r55 20 31 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.865
+ $Y2=0
r56 20 22 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.61
+ $Y2=0
r57 18 23 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r58 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r59 14 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r60 12 17 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.695 $Y=0 $X2=0.69
+ $Y2=0
r61 12 13 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.695 $Y=0 $X2=0.92
+ $Y2=0
r62 11 22 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.61
+ $Y2=0
r63 11 13 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.145 $Y=0 $X2=0.92
+ $Y2=0
r64 7 13 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=0.085 $X2=0.92
+ $Y2=0
r65 7 9 7.30937 $w=4.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.92 $Y=0.085
+ $X2=0.92 $Y2=0.36
r66 2 34 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.685
+ $Y=0.235 $X2=1.85 $Y2=0.36
r67 1 9 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=0.725
+ $Y=0.235 $X2=0.92 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HD__O31A_1%A_253_47# 1 2 7 10 11 12
c23 11 0 1.90303e-19 $X=1.485 $Y=0.74
r24 12 14 5.03913 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.36 $Y=0.655
+ $X2=2.36 $Y2=0.56
r25 10 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.245 $Y=0.74
+ $X2=2.36 $Y2=0.655
r26 10 11 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.245 $Y=0.74
+ $X2=1.485 $Y2=0.74
r27 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.4 $Y=0.655
+ $X2=1.485 $Y2=0.74
r28 7 9 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.4 $Y=0.655 $X2=1.4
+ $Y2=0.56
r29 2 14 182 $w=1.7e-07 $l=3.99061e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.235 $X2=2.33 $Y2=0.56
r30 1 9 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.265
+ $Y=0.235 $X2=1.4 $Y2=0.56
.ends


* File: sky130_fd_sc_hd__and4_2.spice
* Created: Tue Sep  1 18:58:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__and4_2.pex.spice"
.subckt sky130_fd_sc_hd__and4_2  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1010 A_109_47# N_A_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1092 PD=0.715 PS=1.36 NRD=26.424 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1000 A_198_47# N_B_M1000_g A_109_47# VNB NSHORT L=0.15 W=0.42 AD=0.0798
+ AS=0.06195 PD=0.8 PS=0.715 NRD=38.568 NRS=26.424 M=1 R=2.8 SA=75000.6
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1009 A_304_47# N_C_M1009_g A_198_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0798 PD=0.75 PS=0.8 NRD=31.428 NRS=38.568 M=1 R=2.8 SA=75001.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_D_M1011_g A_304_47# VNB NSHORT L=0.15 W=0.42 AD=0.137501
+ AS=0.0693 PD=0.993084 PS=0.75 NRD=94.992 NRS=31.428 M=1 R=2.8 SA=75001.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_47#_M1002_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.212799 PD=0.98 PS=1.53692 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75001.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1002_d N_A_27_47#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.195 PD=0.98 PS=1.9 NRD=10.152 NRS=6.456 M=1 R=4.33333
+ SA=75002.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_27_47#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07455 AS=0.1092 PD=0.775 PS=1.36 NRD=18.7544 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_27_47#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0777 AS=0.07455 PD=0.79 PS=0.775 NRD=21.0987 NRS=16.4101 M=1 R=2.8
+ SA=75000.7 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1001 N_A_27_47#_M1001_d N_C_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0777 PD=0.7 PS=0.79 NRD=0 NRS=21.0987 M=1 R=2.8 SA=75001.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_A_27_47#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.165604 AS=0.0588 PD=0.955352 PS=0.7 NRD=123.105 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.394296 PD=1.33 PS=2.27465 NRD=0 NRS=14.7553 M=1 R=6.66667
+ SA=75001.3 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1008 N_X_M1003_d N_A_27_47#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.3 PD=1.33 PS=2.6 NRD=10.8153 NRS=4.9053 M=1 R=6.66667 SA=75001.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__and4_2.pxi.spice"
*
.ends
*
*

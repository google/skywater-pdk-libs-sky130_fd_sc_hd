* File: sky130_fd_sc_hd__o21ba_1.spice
* Created: Tue Sep  1 19:21:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o21ba_1.pex.spice"
.subckt sky130_fd_sc_hd__o21ba_1  VNB VPB B1_N A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_79_199#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121799 AS=0.169 PD=1.19673 PS=1.82 NRD=5.532 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1002 N_A_222_93#_M1002_d N_B1_N_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0787009 PD=1.36 PS=0.773271 NRD=0 NRS=7.14 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_448_47#_M1009_d N_A_222_93#_M1009_g N_A_79_199#_M1009_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.10725 AS=0.169 PD=0.98 PS=1.82 NRD=10.152 NRS=0 M=1
+ R=4.33333 SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_448_47#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.10725 PD=0.92 PS=0.98 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1008 N_A_448_47#_M1008_d N_A1_M1008_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.08775 PD=1.83 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_79_199#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26162 AS=0.26 PD=1.99296 PS=2.52 NRD=14.7553 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1003 N_A_222_93#_M1003_d N_B1_N_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1176 AS=0.10988 PD=1.4 PS=0.837042 NRD=0 NRS=96.9043 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_79_199#_M1004_d N_A_222_93#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1 AD=0.165 AS=0.3 PD=1.33 PS=2.6 NRD=10.8153 NRS=6.8753 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1001 A_544_297# N_A2_M1001_g N_A_79_199#_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.165 PD=1.21 PS=1.33 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_544_297# VPB PHIGHVT L=0.15 W=1 AD=0.28
+ AS=0.105 PD=2.56 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75001.1 SB=75000.2
+ A=0.15 P=2.3 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__o21ba_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor2b_1.pxi.spice
* Created: Tue Sep  1 19:17:59 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2B_1%B_N N_B_N_M1003_g N_B_N_M1005_g N_B_N_c_44_n
+ N_B_N_c_45_n B_N B_N PM_SKY130_FD_SC_HD__NOR2B_1%B_N
x_PM_SKY130_FD_SC_HD__NOR2B_1%A N_A_M1001_g N_A_M1000_g A N_A_c_74_n N_A_c_75_n
+ PM_SKY130_FD_SC_HD__NOR2B_1%A
x_PM_SKY130_FD_SC_HD__NOR2B_1%A_74_47# N_A_74_47#_M1003_s N_A_74_47#_M1005_s
+ N_A_74_47#_M1004_g N_A_74_47#_M1002_g N_A_74_47#_c_122_n N_A_74_47#_c_118_n
+ N_A_74_47#_c_112_n N_A_74_47#_c_119_n N_A_74_47#_c_113_n N_A_74_47#_c_114_n
+ N_A_74_47#_c_115_n N_A_74_47#_c_116_n PM_SKY130_FD_SC_HD__NOR2B_1%A_74_47#
x_PM_SKY130_FD_SC_HD__NOR2B_1%VPWR N_VPWR_M1005_d N_VPWR_c_182_n VPWR
+ N_VPWR_c_183_n N_VPWR_c_184_n N_VPWR_c_181_n N_VPWR_c_186_n
+ PM_SKY130_FD_SC_HD__NOR2B_1%VPWR
x_PM_SKY130_FD_SC_HD__NOR2B_1%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_212_n N_Y_c_207_n
+ N_Y_c_208_n Y N_Y_c_210_n N_Y_c_209_n PM_SKY130_FD_SC_HD__NOR2B_1%Y
x_PM_SKY130_FD_SC_HD__NOR2B_1%VGND N_VGND_M1003_d N_VGND_M1004_d N_VGND_c_246_n
+ N_VGND_c_247_n N_VGND_c_248_n N_VGND_c_249_n N_VGND_c_250_n VGND
+ N_VGND_c_251_n N_VGND_c_252_n PM_SKY130_FD_SC_HD__NOR2B_1%VGND
cc_1 VNB N_B_N_M1003_g 0.0357768f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.445
cc_2 VNB N_B_N_c_44_n 0.0413585f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_3 VNB N_B_N_c_45_n 0.0106322f $X=-0.19 $Y=-0.24 $X2=0.707 $Y2=1.16
cc_4 VNB B_N 0.0263972f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB A 0.00205316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_c_74_n 0.0253382f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_A_c_75_n 0.0169902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_74_47#_c_112_n 0.00758253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_74_47#_c_113_n 0.00490456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_74_47#_c_114_n 0.00266793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_74_47#_c_115_n 0.0273743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_74_47#_c_116_n 0.0197371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_181_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_207_n 0.0183975f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_15 VNB N_Y_c_208_n 0.00383112f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_Y_c_209_n 0.0200631f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_17 VNB N_VGND_c_246_n 0.00697301f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_18 VNB N_VGND_c_247_n 0.0149623f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_19 VNB N_VGND_c_248_n 0.0210804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_249_n 0.0259297f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_21 VNB N_VGND_c_250_n 0.00403597f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_22 VNB N_VGND_c_251_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_252_n 0.146507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_B_N_M1005_g 0.0270962f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.695
cc_25 VPB N_B_N_c_44_n 0.0183666f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_26 VPB N_B_N_c_45_n 8.10111e-19 $X=-0.19 $Y=1.305 $X2=0.707 $Y2=1.16
cc_27 VPB B_N 0.00949562f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_28 VPB N_A_M1000_g 0.0208466f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.695
cc_29 VPB A 0.00217973f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_c_74_n 0.00637895f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_31 VPB N_A_74_47#_M1002_g 0.0225996f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_A_74_47#_c_118_n 0.00189339f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_33 VPB N_A_74_47#_c_119_n 0.00314759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_74_47#_c_113_n 0.00553539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_74_47#_c_115_n 0.00706905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_182_n 0.0215995f $X=-0.19 $Y=1.305 $X2=0.71 $Y2=1.695
cc_37 VPB N_VPWR_c_183_n 0.0299875f $X=-0.19 $Y=1.305 $X2=0.707 $Y2=1.16
cc_38 VPB N_VPWR_c_184_n 0.0305629f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_39 VPB N_VPWR_c_181_n 0.0676679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_186_n 0.00507883f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_41 VPB N_Y_c_210_n 0.0361418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_Y_c_209_n 0.027368f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_43 N_B_N_M1005_g N_A_M1000_g 0.01777f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_44 N_B_N_c_45_n A 0.00201034f $X=0.707 $Y=1.16 $X2=0 $Y2=0
cc_45 N_B_N_c_45_n N_A_c_74_n 0.0222918f $X=0.707 $Y=1.16 $X2=0 $Y2=0
cc_46 N_B_N_M1003_g N_A_c_75_n 0.0181749f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_47 N_B_N_M1005_g N_A_74_47#_c_122_n 0.0141126f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_48 N_B_N_M1003_g N_A_74_47#_c_112_n 0.00277988f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_49 N_B_N_c_44_n N_A_74_47#_c_112_n 0.00498936f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_50 N_B_N_M1005_g N_A_74_47#_c_119_n 0.00671406f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_51 N_B_N_c_44_n N_A_74_47#_c_119_n 0.00321379f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_52 N_B_N_M1003_g N_A_74_47#_c_113_n 0.0121975f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_53 N_B_N_M1005_g N_A_74_47#_c_113_n 0.00677654f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_54 N_B_N_c_44_n N_A_74_47#_c_113_n 0.0146708f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_55 N_B_N_c_45_n N_A_74_47#_c_113_n 0.00504081f $X=0.707 $Y=1.16 $X2=0 $Y2=0
cc_56 B_N N_A_74_47#_c_113_n 0.0438196f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B_N_M1005_g N_VPWR_c_182_n 0.00397807f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_58 N_B_N_M1005_g N_VPWR_c_183_n 0.00327927f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_59 N_B_N_M1005_g N_VPWR_c_181_n 0.00417489f $X=0.71 $Y=1.695 $X2=0 $Y2=0
cc_60 N_B_N_M1003_g N_VGND_c_246_n 0.0100744f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_61 N_B_N_M1003_g N_VGND_c_249_n 0.00523996f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_62 B_N N_VGND_c_249_n 0.00375784f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_B_N_M1003_g N_VGND_c_252_n 0.0104475f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_64 B_N N_VGND_c_252_n 0.00623997f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_M1000_g N_A_74_47#_M1002_g 0.0498482f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1000_g N_A_74_47#_c_122_n 0.0142825f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_67 A N_A_74_47#_c_122_n 0.0225917f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_c_74_n N_A_74_47#_c_122_n 0.00110992f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_69 A N_A_74_47#_c_118_n 0.00486391f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_74_n N_A_74_47#_c_118_n 0.00151515f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1000_g N_A_74_47#_c_119_n 7.96426e-19 $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_A_74_47#_c_113_n 8.8363e-19 $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_73 A N_A_74_47#_c_113_n 0.0135485f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_74_n N_A_74_47#_c_113_n 6.58322e-19 $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_c_75_n N_A_74_47#_c_113_n 5.88788e-19 $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_76 A N_A_74_47#_c_114_n 0.0107754f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_c_74_n N_A_74_47#_c_114_n 5.85984e-19 $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_78 A N_A_74_47#_c_115_n 5.75929e-19 $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_74_n N_A_74_47#_c_115_n 0.0498482f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_75_n N_A_74_47#_c_116_n 0.0124776f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VPWR_c_182_n 0.0165696f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_VPWR_c_184_n 0.0046653f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_VPWR_c_181_n 0.00783311f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_84 N_A_c_75_n N_Y_c_212_n 0.00517383f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_85 A N_Y_c_208_n 0.00725012f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_74_n N_Y_c_208_n 0.00177728f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_c_75_n N_Y_c_208_n 0.00231966f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_Y_c_210_n 0.00168712f $X=1.25 $Y=1.985 $X2=0 $Y2=0
cc_89 A N_VGND_c_246_n 0.00872494f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_74_n N_VGND_c_246_n 0.00174866f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_c_75_n N_VGND_c_246_n 0.00166284f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_c_75_n N_VGND_c_251_n 0.00541359f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_75_n N_VGND_c_252_n 0.00970758f $X=1.16 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_74_47#_c_122_n N_VPWR_M1005_d 0.00827116f $X=1.535 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_74_47#_M1002_g N_VPWR_c_182_n 0.00289549f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_74_47#_c_122_n N_VPWR_c_182_n 0.0213829f $X=1.535 $Y=1.595 $X2=0 $Y2=0
cc_97 N_A_74_47#_c_119_n N_VPWR_c_182_n 0.00336569f $X=0.545 $Y=1.595 $X2=0
+ $Y2=0
cc_98 N_A_74_47#_M1002_g N_VPWR_c_184_n 0.00541359f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_74_47#_M1002_g N_VPWR_c_181_n 0.0106743f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_74_47#_c_119_n N_VPWR_c_181_n 0.00997842f $X=0.545 $Y=1.595 $X2=0
+ $Y2=0
cc_101 N_A_74_47#_c_122_n A_265_297# 0.00559765f $X=1.535 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_74_47#_c_116_n N_Y_c_212_n 0.0109314f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_74_47#_c_114_n N_Y_c_207_n 0.0200688f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_74_47#_c_115_n N_Y_c_207_n 0.00440824f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_74_47#_c_116_n N_Y_c_207_n 0.0104021f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_74_47#_c_122_n N_Y_c_208_n 0.00531927f $X=1.535 $Y=1.595 $X2=0 $Y2=0
cc_107 N_A_74_47#_c_114_n N_Y_c_208_n 0.00217156f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_74_47#_c_116_n N_Y_c_208_n 9.83966e-19 $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_74_47#_M1002_g N_Y_c_210_n 0.0105468f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_74_47#_c_122_n N_Y_c_210_n 0.0023139f $X=1.535 $Y=1.595 $X2=0 $Y2=0
cc_111 N_A_74_47#_c_114_n N_Y_c_210_n 0.00400794f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_74_47#_c_115_n N_Y_c_210_n 0.00283915f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_74_47#_M1002_g N_Y_c_209_n 0.00632756f $X=1.61 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_74_47#_c_118_n N_Y_c_209_n 0.0117284f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_115 N_A_74_47#_c_114_n N_Y_c_209_n 0.012744f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_74_47#_c_115_n N_Y_c_209_n 0.00622964f $X=1.7 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_74_47#_c_116_n N_Y_c_209_n 0.00281769f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_74_47#_c_122_n N_VGND_c_246_n 0.00345418f $X=1.535 $Y=1.595 $X2=0
+ $Y2=0
cc_119 N_A_74_47#_c_112_n N_VGND_c_246_n 0.0125167f $X=0.585 $Y=0.457 $X2=0
+ $Y2=0
cc_120 N_A_74_47#_c_113_n N_VGND_c_246_n 0.0240171f $X=0.545 $Y=1.51 $X2=0 $Y2=0
cc_121 N_A_74_47#_c_116_n N_VGND_c_248_n 0.00327039f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_74_47#_c_112_n N_VGND_c_249_n 0.011702f $X=0.585 $Y=0.457 $X2=0 $Y2=0
cc_123 N_A_74_47#_c_116_n N_VGND_c_251_n 0.00423334f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_74_47#_M1003_s N_VGND_c_252_n 0.00223287f $X=0.37 $Y=0.235 $X2=0
+ $Y2=0
cc_125 N_A_74_47#_c_112_n N_VGND_c_252_n 0.0117059f $X=0.585 $Y=0.457 $X2=0
+ $Y2=0
cc_126 N_A_74_47#_c_116_n N_VGND_c_252_n 0.00685219f $X=1.7 $Y=0.995 $X2=0 $Y2=0
cc_127 N_VPWR_c_181_n A_265_297# 0.00897657f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_128 N_VPWR_c_181_n N_Y_M1002_d 0.00209319f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_182_n N_Y_c_210_n 0.0216723f $X=1.04 $Y=2 $X2=0 $Y2=0
cc_130 N_VPWR_c_184_n N_Y_c_210_n 0.0373607f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_131 N_VPWR_c_181_n N_Y_c_210_n 0.0212464f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_132 N_Y_c_207_n N_VGND_M1004_d 0.00280958f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_133 N_Y_c_208_n N_VGND_c_246_n 0.00751224f $X=1.565 $Y=0.81 $X2=0 $Y2=0
cc_134 N_Y_c_207_n N_VGND_c_247_n 0.00162138f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_135 N_Y_c_207_n N_VGND_c_248_n 0.030716f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_136 N_Y_c_212_n N_VGND_c_251_n 0.0188385f $X=1.4 $Y=0.39 $X2=0 $Y2=0
cc_137 N_Y_c_207_n N_VGND_c_251_n 0.00198102f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_138 N_Y_M1001_d N_VGND_c_252_n 0.00215201f $X=1.265 $Y=0.235 $X2=0 $Y2=0
cc_139 N_Y_c_212_n N_VGND_c_252_n 0.0122019f $X=1.4 $Y=0.39 $X2=0 $Y2=0
cc_140 N_Y_c_207_n N_VGND_c_252_n 0.00806399f $X=2.035 $Y=0.81 $X2=0 $Y2=0

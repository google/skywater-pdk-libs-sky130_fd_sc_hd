* File: sky130_fd_sc_hd__buf_6.pxi.spice
* Created: Tue Sep  1 18:59:23 2020
* 
x_PM_SKY130_FD_SC_HD__BUF_6%A N_A_M1001_g N_A_M1006_g N_A_M1012_g N_A_M1008_g A
+ A N_A_c_81_n N_A_c_82_n PM_SKY130_FD_SC_HD__BUF_6%A
x_PM_SKY130_FD_SC_HD__BUF_6%A_161_47# N_A_161_47#_M1001_s N_A_161_47#_M1006_s
+ N_A_161_47#_M1002_g N_A_161_47#_M1000_g N_A_161_47#_M1004_g
+ N_A_161_47#_M1003_g N_A_161_47#_M1007_g N_A_161_47#_M1005_g
+ N_A_161_47#_M1013_g N_A_161_47#_M1009_g N_A_161_47#_M1014_g
+ N_A_161_47#_M1010_g N_A_161_47#_M1015_g N_A_161_47#_M1011_g
+ N_A_161_47#_c_155_n N_A_161_47#_c_151_n N_A_161_47#_c_161_n
+ N_A_161_47#_c_139_n N_A_161_47#_c_140_n N_A_161_47#_c_169_n
+ N_A_161_47#_c_141_n N_A_161_47#_c_142_n N_A_161_47#_c_214_p
+ N_A_161_47#_c_143_n N_A_161_47#_c_144_n PM_SKY130_FD_SC_HD__BUF_6%A_161_47#
x_PM_SKY130_FD_SC_HD__BUF_6%VPWR N_VPWR_M1006_d N_VPWR_M1008_d N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_M1011_d N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n VPWR VPWR N_VPWR_c_279_n
+ N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_267_n
+ PM_SKY130_FD_SC_HD__BUF_6%VPWR
x_PM_SKY130_FD_SC_HD__BUF_6%X N_X_M1002_d N_X_M1007_d N_X_M1014_d N_X_M1000_s
+ N_X_M1005_s N_X_M1010_s N_X_c_389_p N_X_c_374_n N_X_c_344_n N_X_c_345_n
+ N_X_c_346_n N_X_c_347_n N_X_c_338_n N_X_c_341_n X N_X_c_340_n
+ PM_SKY130_FD_SC_HD__BUF_6%X
x_PM_SKY130_FD_SC_HD__BUF_6%VGND N_VGND_M1001_d N_VGND_M1012_d N_VGND_M1004_s
+ N_VGND_M1013_s N_VGND_M1015_s N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n
+ N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n VGND VGND N_VGND_c_417_n
+ N_VGND_c_418_n N_VGND_c_419_n N_VGND_c_420_n N_VGND_c_421_n
+ PM_SKY130_FD_SC_HD__BUF_6%VGND
cc_1 VNB N_A_M1001_g 0.0242802f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.56
cc_2 VNB N_A_M1006_g 5.16789e-19 $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.985
cc_3 VNB N_A_M1012_g 0.0175136f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=0.56
cc_4 VNB N_A_M1008_g 4.2558e-19 $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.985
cc_5 VNB A 0.0109395f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.105
cc_6 VNB N_A_c_81_n 0.040848f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_7 VNB N_A_c_82_n 0.0262097f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.16
cc_8 VNB N_A_161_47#_M1002_g 0.0169536f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.025
cc_9 VNB N_A_161_47#_M1000_g 4.13034e-19 $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.295
cc_10 VNB N_A_161_47#_M1004_g 0.0170351f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.105
cc_11 VNB N_A_161_47#_M1003_g 4.47359e-19 $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_12 VNB N_A_161_47#_M1007_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_161_47#_M1005_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.16
cc_14 VNB N_A_161_47#_M1013_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_161_47#_M1009_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_161_47#_M1014_g 0.0160724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_161_47#_M1010_g 3.74796e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_161_47#_M1015_g 0.0233973f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_161_47#_M1011_g 7.17859e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_161_47#_c_139_n 0.00178841f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_161_47#_c_140_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_161_47#_c_141_n 0.00157323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_161_47#_c_142_n 3.48073e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_161_47#_c_143_n 0.00100657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_161_47#_c_144_n 0.107025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_267_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_338_n 0.00154078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB X 0.00226381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_340_n 0.00250845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_406_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.105
cc_31 VNB N_VGND_c_407_n 0.00354062f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_32 VNB N_VGND_c_408_n 0.0151681f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_33 VNB N_VGND_c_409_n 3.15634e-19 $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.16
cc_34 VNB N_VGND_c_410_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.195
cc_35 VNB N_VGND_c_411_n 0.0103361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_412_n 0.0317254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_413_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_414_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_415_n 0.0173211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_416_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_417_n 0.0112541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_418_n 0.01186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_419_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_420_n 0.00436716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_421_n 0.230426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_A_M1006_g 0.0274372f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.985
cc_47 VPB N_A_M1008_g 0.0197846f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.985
cc_48 VPB A 0.0118256f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.105
cc_49 VPB N_A_161_47#_M1000_g 0.0186264f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.295
cc_50 VPB N_A_161_47#_M1003_g 0.0189288f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_51 VPB N_A_161_47#_M1005_g 0.0177798f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.16
cc_52 VPB N_A_161_47#_M1009_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_161_47#_M1010_g 0.0177798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_161_47#_M1011_g 0.0266676f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_161_47#_c_151_n 0.00117749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_161_47#_c_142_n 0.00164506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_268_n 0.00516914f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.105
cc_58 VPB N_VPWR_c_269_n 0.00169924f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_59 VPB N_VPWR_c_270_n 0.0128097f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_60 VPB N_VPWR_c_271_n 3.03604e-19 $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.16
cc_61 VPB N_VPWR_c_272_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_273_n 0.0103102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_274_n 0.0452743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_275_n 0.0159859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_276_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_277_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_278_n 0.00340355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_279_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_280_n 0.0124787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_281_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_282_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_267_n 0.0555743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_341_n 0.00177728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB X 0.00226906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_X_c_340_n 0.00295437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 N_A_M1012_g N_A_161_47#_M1002_g 0.0225534f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_77 N_A_M1008_g N_A_161_47#_M1000_g 0.0225534f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1001_g N_A_161_47#_c_155_n 0.0110414f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_79 N_A_M1012_g N_A_161_47#_c_155_n 0.0066297f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_80 N_A_M1006_g N_A_161_47#_c_151_n 0.00229676f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_M1008_g N_A_161_47#_c_151_n 8.84614e-19 $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_82 A N_A_161_47#_c_151_n 0.0223559f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_c_82_n N_A_161_47#_c_151_n 6.77113e-19 $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_M1006_g N_A_161_47#_c_161_n 0.0091348f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_85 N_A_M1008_g N_A_161_47#_c_161_n 0.0101539f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_86 N_A_M1012_g N_A_161_47#_c_139_n 0.00895754f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_87 A N_A_161_47#_c_139_n 0.00553612f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_88 N_A_M1001_g N_A_161_47#_c_140_n 0.00871241f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_89 N_A_M1012_g N_A_161_47#_c_140_n 0.00110555f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_90 A N_A_161_47#_c_140_n 0.026868f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_91 N_A_c_82_n N_A_161_47#_c_140_n 0.00213429f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_A_161_47#_c_169_n 0.0111745f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_93 A N_A_161_47#_c_169_n 0.00553612f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A_M1012_g N_A_161_47#_c_141_n 0.0037087f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_95 A N_A_161_47#_c_142_n 0.00543401f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A_c_82_n N_A_161_47#_c_142_n 0.00415064f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_97 A N_A_161_47#_c_143_n 0.0146413f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A_c_82_n N_A_161_47#_c_143_n 0.00138162f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_99 A N_A_161_47#_c_144_n 2.21007e-19 $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_c_82_n N_A_161_47#_c_144_n 0.0225534f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_M1006_g N_VPWR_c_268_n 0.00316354f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_102 A N_VPWR_c_268_n 0.0139638f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_103 N_A_c_81_n N_VPWR_c_268_n 0.00124637f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_M1008_g N_VPWR_c_269_n 0.00150833f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_M1006_g N_VPWR_c_277_n 0.00541359f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_M1008_g N_VPWR_c_277_n 0.00541359f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_M1006_g N_VPWR_c_267_n 0.0106288f $X=0.73 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1008_g N_VPWR_c_267_n 0.00952874f $X=1.15 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_M1001_g N_VGND_c_406_n 0.00316354f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_110 A N_VGND_c_406_n 0.00564094f $X=0.89 $Y=1.105 $X2=0 $Y2=0
cc_111 N_A_c_81_n N_VGND_c_406_n 0.00315359f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_M1012_g N_VGND_c_407_n 0.00146448f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_M1001_g N_VGND_c_415_n 0.00541359f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_114 N_A_M1012_g N_VGND_c_415_n 0.00424416f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_VGND_c_421_n 0.0106288f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_M1012_g N_VGND_c_421_n 0.00576327f $X=1.15 $Y=0.56 $X2=0 $Y2=0
cc_117 N_A_161_47#_c_169_n N_VPWR_M1008_d 0.00304347f $X=1.355 $Y=1.57 $X2=0
+ $Y2=0
cc_118 N_A_161_47#_M1000_g N_VPWR_c_269_n 0.00997222f $X=1.57 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A_161_47#_M1003_g N_VPWR_c_269_n 6.64064e-19 $X=1.99 $Y=1.985 $X2=0
+ $Y2=0
cc_120 N_A_161_47#_c_169_n N_VPWR_c_269_n 0.014319f $X=1.355 $Y=1.57 $X2=0 $Y2=0
cc_121 N_A_161_47#_M1000_g N_VPWR_c_270_n 0.00505556f $X=1.57 $Y=1.985 $X2=0
+ $Y2=0
cc_122 N_A_161_47#_M1003_g N_VPWR_c_270_n 0.0046653f $X=1.99 $Y=1.985 $X2=0
+ $Y2=0
cc_123 N_A_161_47#_M1000_g N_VPWR_c_271_n 6.76314e-19 $X=1.57 $Y=1.985 $X2=0
+ $Y2=0
cc_124 N_A_161_47#_M1003_g N_VPWR_c_271_n 0.0111118f $X=1.99 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_161_47#_M1005_g N_VPWR_c_271_n 0.0110878f $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_126 N_A_161_47#_M1009_g N_VPWR_c_271_n 6.72101e-19 $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_161_47#_M1005_g N_VPWR_c_272_n 6.72101e-19 $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_161_47#_M1009_g N_VPWR_c_272_n 0.0110878f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_A_161_47#_M1010_g N_VPWR_c_272_n 0.0110878f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_161_47#_M1011_g N_VPWR_c_272_n 6.72101e-19 $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_161_47#_c_144_n N_VPWR_c_272_n 3.70191e-19 $X=3.67 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_161_47#_M1010_g N_VPWR_c_274_n 8.11858e-19 $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_161_47#_M1011_g N_VPWR_c_274_n 0.0161769f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_161_47#_c_161_n N_VPWR_c_277_n 0.0189039f $X=0.94 $Y=2.31 $X2=0 $Y2=0
cc_135 N_A_161_47#_M1005_g N_VPWR_c_279_n 0.0046653f $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_161_47#_M1009_g N_VPWR_c_279_n 0.0046653f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_161_47#_M1010_g N_VPWR_c_280_n 0.0046653f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_161_47#_M1011_g N_VPWR_c_280_n 0.0046653f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_161_47#_M1006_s N_VPWR_c_267_n 0.00215201f $X=0.805 $Y=1.485 $X2=0
+ $Y2=0
cc_140 N_A_161_47#_M1000_g N_VPWR_c_267_n 0.00858194f $X=1.57 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_161_47#_M1003_g N_VPWR_c_267_n 0.00796766f $X=1.99 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_161_47#_M1005_g N_VPWR_c_267_n 0.00796766f $X=2.41 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_161_47#_M1009_g N_VPWR_c_267_n 0.00796766f $X=2.83 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_161_47#_M1010_g N_VPWR_c_267_n 0.00796766f $X=3.25 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_161_47#_M1011_g N_VPWR_c_267_n 0.00796766f $X=3.67 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_161_47#_c_161_n N_VPWR_c_267_n 0.0122217f $X=0.94 $Y=2.31 $X2=0 $Y2=0
cc_147 N_A_161_47#_c_144_n N_X_c_344_n 3.16187e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_161_47#_c_144_n N_X_c_345_n 2.95142e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_161_47#_c_144_n N_X_c_346_n 3.16187e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_161_47#_c_144_n N_X_c_347_n 2.95142e-19 $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_161_47#_M1002_g N_X_c_338_n 6.92734e-19 $X=1.57 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_161_47#_c_139_n N_X_c_338_n 0.00808484f $X=1.355 $Y=0.82 $X2=0 $Y2=0
cc_153 N_A_161_47#_c_214_p N_X_c_338_n 0.0104485f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_161_47#_c_144_n N_X_c_338_n 0.00213429f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_161_47#_M1000_g N_X_c_341_n 6.26722e-19 $X=1.57 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_161_47#_c_142_n N_X_c_341_n 0.00314617f $X=1.44 $Y=1.485 $X2=0 $Y2=0
cc_157 N_A_161_47#_c_214_p N_X_c_341_n 0.00928852f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_161_47#_c_144_n N_X_c_341_n 0.00211055f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_161_47#_M1004_g X 0.0128214f $X=1.99 $Y=0.56 $X2=0 $Y2=0
cc_160 N_A_161_47#_M1003_g X 0.014825f $X=1.99 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_161_47#_c_144_n X 0.0029023f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_161_47#_M1004_g N_X_c_340_n 0.00200301f $X=1.99 $Y=0.56 $X2=0 $Y2=0
cc_163 N_A_161_47#_M1003_g N_X_c_340_n 0.00285078f $X=1.99 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_161_47#_M1007_g N_X_c_340_n 0.0135801f $X=2.41 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_161_47#_M1005_g N_X_c_340_n 0.0173868f $X=2.41 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A_161_47#_M1013_g N_X_c_340_n 0.013882f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_161_47#_M1009_g N_X_c_340_n 0.0178237f $X=2.83 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_161_47#_M1014_g N_X_c_340_n 0.0132046f $X=3.25 $Y=0.56 $X2=0 $Y2=0
cc_169 N_A_161_47#_M1010_g N_X_c_340_n 0.0171762f $X=3.25 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_161_47#_M1015_g N_X_c_340_n 0.00494338f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_171 N_A_161_47#_M1011_g N_X_c_340_n 0.00630163f $X=3.67 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_161_47#_c_214_p N_X_c_340_n 0.0071292f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_161_47#_c_144_n N_X_c_340_n 0.0677348f $X=3.67 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_161_47#_c_139_n N_VGND_M1012_d 0.00164499f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_175 N_A_161_47#_M1002_g N_VGND_c_407_n 0.00137415f $X=1.57 $Y=0.56 $X2=0
+ $Y2=0
cc_176 N_A_161_47#_c_139_n N_VGND_c_407_n 0.0128905f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_177 N_A_161_47#_M1002_g N_VGND_c_408_n 0.00556122f $X=1.57 $Y=0.56 $X2=0
+ $Y2=0
cc_178 N_A_161_47#_M1004_g N_VGND_c_408_n 0.00350562f $X=1.99 $Y=0.56 $X2=0
+ $Y2=0
cc_179 N_A_161_47#_c_139_n N_VGND_c_408_n 8.04923e-19 $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_180 N_A_161_47#_M1002_g N_VGND_c_409_n 6.10735e-19 $X=1.57 $Y=0.56 $X2=0
+ $Y2=0
cc_181 N_A_161_47#_M1004_g N_VGND_c_409_n 0.00787546f $X=1.99 $Y=0.56 $X2=0
+ $Y2=0
cc_182 N_A_161_47#_M1007_g N_VGND_c_409_n 0.00769005f $X=2.41 $Y=0.56 $X2=0
+ $Y2=0
cc_183 N_A_161_47#_M1013_g N_VGND_c_409_n 5.77787e-19 $X=2.83 $Y=0.56 $X2=0
+ $Y2=0
cc_184 N_A_161_47#_M1007_g N_VGND_c_410_n 5.77787e-19 $X=2.41 $Y=0.56 $X2=0
+ $Y2=0
cc_185 N_A_161_47#_M1013_g N_VGND_c_410_n 0.00769005f $X=2.83 $Y=0.56 $X2=0
+ $Y2=0
cc_186 N_A_161_47#_M1014_g N_VGND_c_410_n 0.00769005f $X=3.25 $Y=0.56 $X2=0
+ $Y2=0
cc_187 N_A_161_47#_M1015_g N_VGND_c_410_n 5.77787e-19 $X=3.67 $Y=0.56 $X2=0
+ $Y2=0
cc_188 N_A_161_47#_c_144_n N_VGND_c_410_n 3.77859e-19 $X=3.67 $Y=1.16 $X2=0
+ $Y2=0
cc_189 N_A_161_47#_M1014_g N_VGND_c_412_n 7.33828e-19 $X=3.25 $Y=0.56 $X2=0
+ $Y2=0
cc_190 N_A_161_47#_M1015_g N_VGND_c_412_n 0.0125262f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_161_47#_c_155_n N_VGND_c_415_n 0.0188551f $X=0.94 $Y=0.38 $X2=0 $Y2=0
cc_192 N_A_161_47#_c_139_n N_VGND_c_415_n 0.00193763f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_193 N_A_161_47#_M1007_g N_VGND_c_417_n 0.00350562f $X=2.41 $Y=0.56 $X2=0
+ $Y2=0
cc_194 N_A_161_47#_M1013_g N_VGND_c_417_n 0.00350562f $X=2.83 $Y=0.56 $X2=0
+ $Y2=0
cc_195 N_A_161_47#_M1014_g N_VGND_c_418_n 0.00350562f $X=3.25 $Y=0.56 $X2=0
+ $Y2=0
cc_196 N_A_161_47#_M1015_g N_VGND_c_418_n 0.0046653f $X=3.67 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_161_47#_M1001_s N_VGND_c_421_n 0.00215201f $X=0.805 $Y=0.235 $X2=0
+ $Y2=0
cc_198 N_A_161_47#_M1002_g N_VGND_c_421_n 0.00973329f $X=1.57 $Y=0.56 $X2=0
+ $Y2=0
cc_199 N_A_161_47#_M1004_g N_VGND_c_421_n 0.00418574f $X=1.99 $Y=0.56 $X2=0
+ $Y2=0
cc_200 N_A_161_47#_M1007_g N_VGND_c_421_n 0.00418574f $X=2.41 $Y=0.56 $X2=0
+ $Y2=0
cc_201 N_A_161_47#_M1013_g N_VGND_c_421_n 0.00418574f $X=2.83 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_161_47#_M1014_g N_VGND_c_421_n 0.00418574f $X=3.25 $Y=0.56 $X2=0
+ $Y2=0
cc_203 N_A_161_47#_M1015_g N_VGND_c_421_n 0.00796766f $X=3.67 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_161_47#_c_155_n N_VGND_c_421_n 0.0122069f $X=0.94 $Y=0.38 $X2=0 $Y2=0
cc_205 N_A_161_47#_c_139_n N_VGND_c_421_n 0.00653201f $X=1.355 $Y=0.82 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_267_n N_X_M1000_s 0.00570907f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_207 N_VPWR_c_267_n N_X_M1005_s 0.00570907f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_208 N_VPWR_c_267_n N_X_M1010_s 0.00570907f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_209 N_VPWR_c_270_n N_X_c_374_n 0.0113958f $X=2.035 $Y=2.72 $X2=0 $Y2=0
cc_210 N_VPWR_c_267_n N_X_c_374_n 0.00646998f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_211 N_VPWR_c_279_n N_X_c_345_n 0.0113958f $X=2.875 $Y=2.72 $X2=0 $Y2=0
cc_212 N_VPWR_c_267_n N_X_c_345_n 0.00646998f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_213 N_VPWR_c_280_n N_X_c_347_n 0.0113958f $X=3.715 $Y=2.72 $X2=0 $Y2=0
cc_214 N_VPWR_c_267_n N_X_c_347_n 0.00646998f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_215 N_VPWR_M1003_d X 0.00103514f $X=2.065 $Y=1.485 $X2=0 $Y2=0
cc_216 N_VPWR_c_271_n X 0.00764235f $X=2.2 $Y=2 $X2=0 $Y2=0
cc_217 N_VPWR_M1003_d N_X_c_340_n 8.43175e-19 $X=2.065 $Y=1.485 $X2=0 $Y2=0
cc_218 N_VPWR_M1009_d N_X_c_340_n 0.00193841f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_219 N_VPWR_c_271_n N_X_c_340_n 0.0070082f $X=2.2 $Y=2 $X2=0 $Y2=0
cc_220 N_VPWR_c_272_n N_X_c_340_n 0.0154647f $X=3.04 $Y=2 $X2=0 $Y2=0
cc_221 N_VPWR_c_274_n N_VGND_c_412_n 0.00942828f $X=3.88 $Y=1.66 $X2=0 $Y2=0
cc_222 X N_VGND_M1004_s 9.03495e-19 $X=2.21 $Y=0.765 $X2=0 $Y2=0
cc_223 N_X_c_340_n N_VGND_M1004_s 7.35111e-19 $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_224 N_X_c_340_n N_VGND_M1013_s 0.00169066f $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_225 N_X_c_389_p N_VGND_c_408_n 0.0113595f $X=1.78 $Y=0.56 $X2=0 $Y2=0
cc_226 X N_VGND_c_408_n 0.00193763f $X=2.21 $Y=0.765 $X2=0 $Y2=0
cc_227 X N_VGND_c_409_n 0.00896031f $X=2.21 $Y=0.765 $X2=0 $Y2=0
cc_228 N_X_c_340_n N_VGND_c_409_n 0.00820188f $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_229 N_X_c_340_n N_VGND_c_410_n 0.0180722f $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_230 N_X_c_344_n N_VGND_c_417_n 0.0111222f $X=2.62 $Y=0.56 $X2=0 $Y2=0
cc_231 N_X_c_340_n N_VGND_c_417_n 0.0042033f $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_232 N_X_c_346_n N_VGND_c_418_n 0.0111222f $X=3.46 $Y=0.56 $X2=0 $Y2=0
cc_233 N_X_c_340_n N_VGND_c_418_n 0.00210921f $X=3.46 $Y=1.175 $X2=0 $Y2=0
cc_234 N_X_M1002_d N_VGND_c_421_n 0.00418657f $X=1.645 $Y=0.235 $X2=0 $Y2=0
cc_235 N_X_M1007_d N_VGND_c_421_n 0.00269036f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_236 N_X_M1014_d N_VGND_c_421_n 0.00415697f $X=3.325 $Y=0.235 $X2=0 $Y2=0
cc_237 N_X_c_389_p N_VGND_c_421_n 0.0064623f $X=1.78 $Y=0.56 $X2=0 $Y2=0
cc_238 N_X_c_344_n N_VGND_c_421_n 0.00641247f $X=2.62 $Y=0.56 $X2=0 $Y2=0
cc_239 N_X_c_346_n N_VGND_c_421_n 0.00641247f $X=3.46 $Y=0.56 $X2=0 $Y2=0
cc_240 X N_VGND_c_421_n 0.00451514f $X=2.21 $Y=0.765 $X2=0 $Y2=0
cc_241 N_X_c_340_n N_VGND_c_421_n 0.0145912f $X=3.46 $Y=1.175 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a221oi_2.pex.spice
* Created: Tue Sep  1 18:52:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A221OI_2%C1 1 3 6 8 10 13 15 16 24
r38 23 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.48 $Y=1.16 $X2=0.9
+ $Y2=1.16
r39 20 23 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.255 $Y=1.16
+ $X2=0.48 $Y2=1.16
r40 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r41 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r42 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=1.325
+ $X2=0.9 $Y2=1.16
r43 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.9 $Y=1.325 $X2=0.9
+ $Y2=1.985
r44 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.9 $Y=0.995 $X2=0.9
+ $Y2=1.16
r45 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995 $X2=0.9
+ $Y2=0.56
r46 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.325
+ $X2=0.48 $Y2=1.16
r47 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.48 $Y=1.325 $X2=0.48
+ $Y2=1.985
r48 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995 $X2=0.48
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%B2 1 3 6 8 10 13 15 19 20 22 23 27 28
c81 28 0 1.81811e-19 $X=1.84 $Y=1.16
c82 27 0 2.75292e-19 $X=1.84 $Y=1.16
c83 20 0 1.54366e-19 $X=3.1 $Y=1.16
r84 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.84
+ $Y=1.16 $X2=1.84 $Y2=1.16
r85 22 23 7.60125 $w=5.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.772 $Y=1.19
+ $X2=1.772 $Y2=1.53
r86 22 28 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=1.772 $Y=1.19
+ $X2=1.772 $Y2=1.16
r87 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=1.16 $X2=3.1 $Y2=1.16
r88 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.1 $Y=1.445
+ $X2=3.1 $Y2=1.16
r89 16 23 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=2.04 $Y=1.53
+ $X2=1.772 $Y2=1.53
r90 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=1.53
+ $X2=3.1 $Y2=1.445
r91 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.935 $Y=1.53
+ $X2=2.04 $Y2=1.53
r92 11 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.325
+ $X2=3.1 $Y2=1.16
r93 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.1 $Y=1.325 $X2=3.1
+ $Y2=1.985
r94 8 20 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=0.995 $X2=3.1
+ $Y2=1.16
r95 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.1 $Y=0.995 $X2=3.1
+ $Y2=0.56
r96 4 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.325
+ $X2=1.84 $Y2=1.16
r97 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.84 $Y=1.325 $X2=1.84
+ $Y2=1.985
r98 1 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=0.995
+ $X2=1.84 $Y2=1.16
r99 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.84 $Y=0.995 $X2=1.84
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%B1 1 3 6 8 10 13 15 22
c43 6 0 1.81811e-19 $X=2.26 $Y=1.985
r44 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.47 $Y=1.16
+ $X2=2.68 $Y2=1.16
r45 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.26 $Y=1.16
+ $X2=2.47 $Y2=1.16
r46 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.16 $X2=2.47 $Y2=1.16
r47 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.16
r48 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.68 $Y=1.325
+ $X2=2.68 $Y2=1.985
r49 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.68 $Y2=1.16
r50 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.68 $Y=0.995
+ $X2=2.68 $Y2=0.56
r51 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.325
+ $X2=2.26 $Y2=1.16
r52 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.26 $Y=1.325 $X2=2.26
+ $Y2=1.985
r53 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=0.995
+ $X2=2.26 $Y2=1.16
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.26 $Y=0.995 $X2=2.26
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A2 1 3 6 8 10 13 17 18 20 21 23 24 25 29 33
c85 29 0 1.50675e-19 $X=4.86 $Y=1.16
c86 18 0 1.80423e-19 $X=3.6 $Y=1.16
c87 8 0 8.35171e-20 $X=4.86 $Y=0.995
r88 30 33 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=4.86 $Y=1.175
+ $X2=5.29 $Y2=1.175
r89 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.86
+ $Y=1.16 $X2=4.86 $Y2=1.16
r90 25 33 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=1.175
+ $X2=5.29 $Y2=1.175
r91 24 30 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=4.82 $Y=1.175 $X2=4.86
+ $Y2=1.175
r92 22 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.735 $Y=1.275
+ $X2=4.82 $Y2=1.175
r93 22 23 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.735 $Y=1.275
+ $X2=4.735 $Y2=1.445
r94 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.65 $Y=1.53
+ $X2=4.735 $Y2=1.445
r95 20 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.65 $Y=1.53
+ $X2=3.765 $Y2=1.53
r96 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=1.16 $X2=3.6 $Y2=1.16
r97 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.6 $Y=1.445
+ $X2=3.765 $Y2=1.53
r98 15 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.6 $Y=1.445
+ $X2=3.6 $Y2=1.16
r99 11 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=1.325
+ $X2=4.86 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.86 $Y=1.325
+ $X2=4.86 $Y2=1.985
r101 8 29 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=0.995
+ $X2=4.86 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.86 $Y=0.995
+ $X2=4.86 $Y2=0.56
r103 4 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.325
+ $X2=3.6 $Y2=1.16
r104 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.6 $Y=1.325 $X2=3.6
+ $Y2=1.985
r105 1 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.995
+ $X2=3.6 $Y2=1.16
r106 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.6 $Y=0.995 $X2=3.6
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A1 1 3 6 8 10 13 15 22
c43 8 0 1.58913e-19 $X=4.44 $Y=0.995
r44 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.23 $Y=1.16
+ $X2=4.44 $Y2=1.16
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.16 $X2=4.23 $Y2=1.16
r46 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.02 $Y=1.16
+ $X2=4.23 $Y2=1.16
r47 15 21 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.23 $Y2=1.175
r48 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=1.325
+ $X2=4.44 $Y2=1.16
r49 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.44 $Y=1.325
+ $X2=4.44 $Y2=1.985
r50 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.44 $Y=0.995
+ $X2=4.44 $Y2=1.16
r51 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.44 $Y=0.995
+ $X2=4.44 $Y2=0.56
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.325
+ $X2=4.02 $Y2=1.16
r53 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.02 $Y=1.325 $X2=4.02
+ $Y2=1.985
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=0.995
+ $X2=4.02 $Y2=1.16
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.02 $Y=0.995 $X2=4.02
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A_27_297# 1 2 3 4 15 17 18 21 24 25 27 29
+ 30 35
c55 35 0 1.24618e-19 $X=2.89 $Y=1.87
c56 30 0 1.24618e-19 $X=2.05 $Y=1.87
c57 25 0 1.50675e-19 $X=1.925 $Y=1.87
r58 35 38 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.89 $Y=1.87 $X2=2.89
+ $Y2=1.96
r59 30 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.05 $Y=1.87 $X2=2.05
+ $Y2=1.96
r60 28 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.175 $Y=1.87
+ $X2=2.05 $Y2=1.87
r61 27 35 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=1.87
+ $X2=2.89 $Y2=1.87
r62 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.765 $Y=1.87
+ $X2=2.175 $Y2=1.87
r63 26 29 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.275 $Y=1.87
+ $X2=1.15 $Y2=1.87
r64 25 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.925 $Y=1.87
+ $X2=2.05 $Y2=1.87
r65 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.925 $Y=1.87
+ $X2=1.275 $Y2=1.87
r66 23 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=1.955
+ $X2=1.15 $Y2=1.87
r67 23 24 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.15 $Y=1.955
+ $X2=1.15 $Y2=2.295
r68 19 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=1.785
+ $X2=1.15 $Y2=1.87
r69 19 21 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.15 $Y=1.785
+ $X2=1.15 $Y2=1.66
r70 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.025 $Y=2.38
+ $X2=1.15 $Y2=2.295
r71 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.025 $Y=2.38
+ $X2=0.435 $Y2=2.38
r72 13 18 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.262 $Y=2.295
+ $X2=0.435 $Y2=2.38
r73 13 15 13.8627 $w=3.43e-07 $l=4.15e-07 $layer=LI1_cond $X=0.262 $Y=2.295
+ $X2=0.262 $Y2=1.88
r74 4 38 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.485 $X2=2.89 $Y2=1.96
r75 3 33 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.485 $X2=2.05 $Y2=1.96
r76 2 21 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.975
+ $Y=1.485 $X2=1.11 $Y2=1.66
r77 1 15 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.27 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%Y 1 2 3 4 19 20 22 23 25 26 27 28 29 38
c72 26 0 1.67842e-19 $X=0.61 $Y=0.765
c73 22 0 8.35171e-20 $X=4.23 $Y=0.73
r74 29 47 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.62
r75 28 47 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.73 $Y=1.53 $X2=0.73
+ $Y2=1.62
r76 27 28 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.73 $Y=1.19
+ $X2=0.73 $Y2=1.53
r77 26 36 3.41797 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0.725
+ $X2=0.69 $Y2=0.725
r78 26 41 3.41797 $w=2.9e-07 $l=2.80936e-07 $layer=LI1_cond $X=0.525 $Y=0.725
+ $X2=0.73 $Y2=0.905
r79 26 27 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.73 $Y=0.92
+ $X2=0.73 $Y2=1.19
r80 26 41 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.73 $Y=0.92
+ $X2=0.73 $Y2=0.905
r81 25 36 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.69 $Y=0.51
+ $X2=0.69 $Y2=0.725
r82 25 38 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.69 $Y=0.51 $X2=0.69
+ $Y2=0.39
r83 22 23 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0.775
+ $X2=4.065 $Y2=0.775
r84 20 23 88.1111 $w=1.78e-07 $l=1.43e-06 $layer=LI1_cond $X=2.635 $Y=0.815
+ $X2=4.065 $Y2=0.815
r85 18 20 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0.775
+ $X2=2.635 $Y2=0.775
r86 18 19 9.3019 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=2.47 $Y=0.775
+ $X2=2.285 $Y2=0.775
r87 14 26 3.10432 $w=1.8e-07 $l=3.7229e-07 $layer=LI1_cond $X=0.855 $Y=0.815
+ $X2=0.525 $Y2=0.725
r88 14 19 88.1111 $w=1.78e-07 $l=1.43e-06 $layer=LI1_cond $X=0.855 $Y=0.815
+ $X2=2.285 $Y2=0.815
r89 4 47 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.485 $X2=0.69 $Y2=1.62
r90 3 22 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.23 $Y2=0.73
r91 2 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.47 $Y2=0.73
r92 1 38 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.69 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A_301_297# 1 2 3 4 5 16 18 20 22 26 28 32
+ 36 39 44 50
c60 28 0 1.50675e-19 $X=4.99 $Y=1.87
c61 22 0 1.50675e-19 $X=4.105 $Y=1.87
c62 20 0 5.9496e-20 $X=3.35 $Y=1.955
r63 44 46 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.47 $Y=2.3 $X2=2.47
+ $Y2=2.38
r64 39 41 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.63 $Y=2.3 $X2=1.63
+ $Y2=2.38
r65 34 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.092 $Y=1.955
+ $X2=5.092 $Y2=1.87
r66 34 36 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=5.092 $Y=1.955
+ $X2=5.092 $Y2=1.96
r67 30 51 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.092 $Y=1.785
+ $X2=5.092 $Y2=1.87
r68 30 32 8.92683 $w=2.03e-07 $l=1.65e-07 $layer=LI1_cond $X=5.092 $Y=1.785
+ $X2=5.092 $Y2=1.62
r69 29 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.355 $Y=1.87
+ $X2=4.23 $Y2=1.87
r70 28 51 2.0246 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.99 $Y=1.87
+ $X2=5.092 $Y2=1.87
r71 28 29 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.99 $Y=1.87
+ $X2=4.355 $Y2=1.87
r72 24 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=1.955
+ $X2=4.23 $Y2=1.87
r73 24 26 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.23 $Y=1.955
+ $X2=4.23 $Y2=1.96
r74 23 49 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=1.87
+ $X2=3.35 $Y2=1.87
r75 22 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.105 $Y=1.87
+ $X2=4.23 $Y2=1.87
r76 22 23 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.105 $Y=1.87
+ $X2=3.475 $Y2=1.87
r77 20 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=1.955
+ $X2=3.35 $Y2=1.87
r78 20 21 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=3.35 $Y=1.955
+ $X2=3.35 $Y2=2.295
r79 19 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.595 $Y=2.38
+ $X2=2.47 $Y2=2.38
r80 18 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.225 $Y=2.38
+ $X2=3.35 $Y2=2.295
r81 18 19 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.225 $Y=2.38
+ $X2=2.595 $Y2=2.38
r82 17 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.755 $Y=2.38
+ $X2=1.63 $Y2=2.38
r83 16 46 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=2.38
+ $X2=2.47 $Y2=2.38
r84 16 17 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.345 $Y=2.38
+ $X2=1.755 $Y2=2.38
r85 5 36 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=4.935
+ $Y=1.485 $X2=5.075 $Y2=1.96
r86 5 32 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=4.935
+ $Y=1.485 $X2=5.075 $Y2=1.62
r87 4 26 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.095
+ $Y=1.485 $X2=4.23 $Y2=1.96
r88 3 49 300 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=2 $X=3.175
+ $Y=1.485 $X2=3.35 $Y2=1.95
r89 2 44 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.485 $X2=2.47 $Y2=2.3
r90 1 39 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.505
+ $Y=1.485 $X2=1.63 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%VPWR 1 2 9 13 16 17 19 20 21 34 35
r70 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r71 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r72 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r73 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r74 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 24 28 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r76 21 29 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r77 21 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 19 31 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.37 $Y2=2.72
r79 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.525 $Y=2.72
+ $X2=4.65 $Y2=2.72
r80 18 34 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.775 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.775 $Y=2.72
+ $X2=4.65 $Y2=2.72
r82 16 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.45 $Y2=2.72
r83 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.81 $Y2=2.72
r84 15 31 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.37 $Y2=2.72
r85 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.81 $Y2=2.72
r86 11 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=2.635
+ $X2=4.65 $Y2=2.72
r87 11 13 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.65 $Y=2.635
+ $X2=4.65 $Y2=2.3
r88 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=2.635
+ $X2=3.81 $Y2=2.72
r89 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.81 $Y=2.635
+ $X2=3.81 $Y2=2.3
r90 2 13 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=1.485 $X2=4.65 $Y2=2.3
r91 1 9 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.485 $X2=3.81 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%VGND 1 2 3 4 13 15 19 23 26 27 29 30 31 52
+ 53 61 67
r71 66 67 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.235
+ $X2=1.715 $Y2=0.235
r72 63 66 0.373774 $w=6.38e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=0.235
+ $X2=1.63 $Y2=0.235
r73 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 60 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r75 59 63 8.59681 $w=6.38e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=0.235
+ $X2=1.61 $Y2=0.235
r76 59 61 9.66931 $w=6.38e-07 $l=1.25e-07 $layer=LI1_cond $X=1.15 $Y=0.235
+ $X2=1.025 $Y2=0.235
r77 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r78 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r79 50 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r80 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r81 47 50 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r82 46 49 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r83 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r84 44 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r85 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r86 41 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r87 41 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r88 40 43 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r89 40 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.715
+ $Y2=0
r90 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r91 37 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r92 36 61 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.025
+ $Y2=0
r93 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r94 34 56 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r95 34 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r96 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r97 31 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r98 29 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.985 $Y=0 $X2=4.83
+ $Y2=0
r99 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0 $X2=5.07
+ $Y2=0
r100 28 52 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.29 $Y2=0
r101 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.07
+ $Y2=0
r102 26 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=2.99
+ $Y2=0
r103 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.355
+ $Y2=0
r104 25 46 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.45
+ $Y2=0
r105 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0 $X2=3.355
+ $Y2=0
r106 21 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.085
+ $X2=5.07 $Y2=0
r107 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.07 $Y=0.085
+ $X2=5.07 $Y2=0.39
r108 17 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0
r109 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0.39
r110 13 56 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.177 $Y2=0
r111 13 15 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.39
r112 4 23 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.935
+ $Y=0.235 $X2=5.07 $Y2=0.39
r113 3 19 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.355 $Y2=0.39
r114 2 66 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.63 $Y2=0.39
r115 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.27 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A_383_47# 1 2 11
r15 8 11 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.05 $Y=0.365
+ $X2=2.89 $Y2=0.365
r16 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.235 $X2=2.89 $Y2=0.39
r17 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.235 $X2=2.05 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A221OI_2%A_735_47# 1 2 7 11 13
c23 13 0 1.58913e-19 $X=4.65 $Y=0.73
r24 11 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=4.69 $Y=0.475
+ $X2=4.69 $Y2=0.365
r25 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.69 $Y=0.475
+ $X2=4.69 $Y2=0.73
r26 7 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.565 $Y=0.365
+ $X2=4.69 $Y2=0.365
r27 7 9 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=4.565 $Y=0.365
+ $X2=3.81 $Y2=0.365
r28 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.235 $X2=4.65 $Y2=0.39
r29 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.235 $X2=4.65 $Y2=0.73
r30 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.235 $X2=3.81 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__dfstp_2.pex.spice
* Created: Tue Sep  1 19:03:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFSTP_2%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.24 $Y=1.235
+ $X2=0.24 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.235 $X2=0.24 $Y2=1.235
r49 15 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.3 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=1.59 $X2=0.3
+ $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.3 $Y=0.88 $X2=0.3
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_27_47# 1 2 9 13 15 17 20 24 28 31 35 36 37
+ 40 42 46 47 50 51 52 54 55 59 61 62 63 64 73 78 85 86 92 93 96
c281 92 0 3.16068e-19 $X=5.155 $Y=1.74
c282 86 0 3.30612e-20 $X=2.765 $Y=1.74
c283 85 0 2.53448e-20 $X=2.765 $Y=1.74
c284 73 0 1.73859e-19 $X=5.29 $Y=1.87
c285 63 0 1.39518e-19 $X=5.145 $Y=1.87
c286 61 0 1.01003e-19 $X=2.385 $Y=1.87
c287 52 0 3.12358e-20 $X=5.05 $Y=0.81
c288 51 0 1.753e-19 $X=5.8 $Y=0.81
c289 47 0 9.52104e-20 $X=2.435 $Y=0.87
c290 46 0 1.76471e-19 $X=2.435 $Y=0.87
c291 40 0 1.78014e-19 $X=0.72 $Y=1.795
c292 24 0 7.39505e-20 $X=5.065 $Y=2.275
r293 93 104 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.155 $Y=1.81
+ $X2=4.965 $Y2=1.81
r294 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.74 $X2=5.155 $Y2=1.74
r295 89 92 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.065 $Y=1.74
+ $X2=5.155 $Y2=1.74
r296 85 88 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.74
+ $X2=2.765 $Y2=1.875
r297 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.74 $X2=2.765 $Y2=1.74
r298 73 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r299 71 86 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.765 $Y2=1.765
r300 71 99 2.12292 $w=3.78e-07 $l=7e-08 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.46 $Y2=1.765
r301 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r302 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.87
+ $X2=0.69 $Y2=1.87
r303 64 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.87
+ $X2=2.53 $Y2=1.87
r304 63 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r305 63 64 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=2.675 $Y2=1.87
r306 62 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.87
+ $X2=0.69 $Y2=1.87
r307 61 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r308 61 62 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=0.835 $Y2=1.87
r309 59 96 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=0.93
+ $X2=5.995 $Y2=0.765
r310 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=0.93 $X2=5.985 $Y2=0.93
r311 55 58 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=5.975 $Y=0.81
+ $X2=5.975 $Y2=0.93
r312 51 55 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.8 $Y=0.81 $X2=5.975
+ $Y2=0.81
r313 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.8 $Y=0.81
+ $X2=5.05 $Y2=0.81
r314 50 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.965 $Y=1.655
+ $X2=4.965 $Y2=1.81
r315 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.965 $Y=0.895
+ $X2=5.05 $Y2=0.81
r316 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.965 $Y=0.895
+ $X2=4.965 $Y2=1.655
r317 47 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.435 $Y=0.87
+ $X2=2.305 $Y2=0.87
r318 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=0.87 $X2=2.435 $Y2=0.87
r319 44 99 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=1.765
r320 44 46 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=0.87
r321 43 78 31.1043 $w=2.7e-07 $l=1.4e-07 $layer=POLY_cond $X=0.75 $Y=1.235
+ $X2=0.89 $Y2=1.235
r322 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.235 $X2=0.75 $Y2=1.235
r323 40 67 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.88
r324 40 42 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.72 $Y=1.795
+ $X2=0.72 $Y2=1.235
r325 39 42 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.72 $Y=0.805
+ $X2=0.72 $Y2=1.235
r326 38 54 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r327 37 67 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.72 $Y2=1.88
r328 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.345 $Y2=1.88
r329 35 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.72 $Y2=0.805
r330 35 36 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.345 $Y2=0.72
r331 29 36 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r332 29 31 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r333 28 96 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.065 $Y=0.445
+ $X2=6.065 $Y2=0.765
r334 22 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=1.74
r335 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=2.275
r336 20 88 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.875
r337 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r338 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r339 11 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r340 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r341 7 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r342 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r343 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r344 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%D 3 7 9 10 14 15
c42 14 0 1.34441e-19 $X=1.855 $Y=1.17
c43 7 0 1.76471e-19 $X=1.83 $Y=2.065
r44 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.335
r45 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.005
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.17 $X2=1.855 $Y2=1.17
r47 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.53
r48 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.17
r49 7 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.335
r50 3 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=0.555
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_193_47# 1 2 9 11 12 15 18 21 23 25 28 31
+ 33 38 40 41 43 44 45 48 52 53 56 57 64
c208 57 0 4.4944e-20 $X=5.31 $Y=1.19
c209 56 0 2.56901e-19 $X=5.31 $Y=1.19
c210 52 0 3.30612e-20 $X=2.99 $Y=0.85
c211 45 0 2.53448e-20 $X=3.135 $Y=1.19
c212 44 0 1.51904e-19 $X=5.165 $Y=1.19
c213 43 0 9.52104e-20 $X=3.027 $Y=1.12
c214 38 0 1.21943e-19 $X=1.1 $Y=1.96
c215 25 0 1.80017e-19 $X=5.605 $Y=2.275
c216 23 0 1.753e-19 $X=5.605 $Y=1.455
c217 9 0 4.43992e-20 $X=2.315 $Y=2.275
r218 64 67 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=1.095
r219 64 66 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=0.765
r220 57 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.26 $X2=5.315 $Y2=1.26
r221 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.31 $Y=1.19
+ $X2=5.31 $Y2=1.19
r222 53 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=0.93 $X2=2.915 $Y2=0.93
r223 52 54 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.965
r224 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.85
r225 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0.85
+ $X2=1.15 $Y2=0.85
r226 44 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.165 $Y=1.19
+ $X2=5.31 $Y2=1.19
r227 44 45 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=5.165 $Y=1.19
+ $X2=3.135 $Y2=1.19
r228 43 45 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.135 $Y2=1.19
r229 43 54 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.027 $Y2=0.965
r230 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=0.85
+ $X2=1.15 $Y2=0.85
r231 40 52 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=2.99 $Y2=0.85
r232 40 41 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=1.295 $Y2=0.85
r233 38 39 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.96
+ $X2=1.12 $Y2=2.045
r234 36 48 54.1147 $w=2.28e-07 $l=1.08e-06 $layer=LI1_cond $X=1.12 $Y=1.93
+ $X2=1.12 $Y2=0.85
r235 36 38 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=1.12 $Y=1.93 $X2=1.12
+ $Y2=1.96
r236 33 48 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.12 $Y=0.68
+ $X2=1.12 $Y2=0.85
r237 33 35 9.01739 $w=2.3e-07 $l=1.7e-07 $layer=LI1_cond $X=1.12 $Y=0.68
+ $X2=1.12 $Y2=0.51
r238 31 39 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=1.125 $Y=2.3
+ $X2=1.125 $Y2=2.045
r239 28 60 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.47 $Y=1.26
+ $X2=5.315 $Y2=1.26
r240 23 28 52.102 $w=1.88e-07 $l=2.09464e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.575 $Y2=1.26
r241 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.605 $Y2=2.275
r242 19 28 36.719 $w=1.88e-07 $l=1.39911e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.575 $Y2=1.26
r243 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.565 $Y2=0.445
r244 18 67 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=1.245
+ $X2=2.855 $Y2=1.095
r245 15 66 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.855 $Y=0.415
+ $X2=2.855 $Y2=0.765
r246 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.855 $Y2=1.245
r247 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.39 $Y2=1.32
r248 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.39 $Y2=1.32
r249 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.315 $Y2=2.275
r250 2 38 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r251 2 31 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=2.3
r252 1 35 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_652_21# 1 2 9 13 15 19 21 25 28 30 31 35
+ 38
c115 38 0 1.30404e-19 $X=4.625 $Y=0.895
c116 35 0 2.11834e-19 $X=4.075 $Y=1.96
c117 28 0 3.15264e-19 $X=4.625 $Y=1.835
c118 21 0 1.75093e-19 $X=4.54 $Y=1.96
r119 36 38 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.435 $Y=0.895
+ $X2=4.625 $Y2=0.895
r120 31 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.905
r121 31 41 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.575
r122 30 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.485 $Y=1.74
+ $X2=3.485 $Y2=1.96
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.74 $X2=3.445 $Y2=1.74
r124 27 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=0.895
r125 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=1.835
r126 23 36 2.53954 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.895
r127 23 25 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.46
r128 22 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.96
+ $X2=4.075 $Y2=1.96
r129 21 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.625 $Y2=1.835
r130 21 22 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.16 $Y2=1.96
r131 17 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=1.96
r132 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=2.21
r133 16 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.485 $Y2=1.96
r134 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=4.075 $Y2=1.96
r135 15 16 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=3.61 $Y2=1.96
r136 13 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.335 $Y=2.275
+ $X2=3.335 $Y2=1.905
r137 9 41 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.335 $Y=0.445
+ $X2=3.335 $Y2=1.575
r138 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.065 $X2=4.075 $Y2=2.21
r139 1 25 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%SET_B 1 3 7 11 14 17 19 23 25 26 28 29 35 36
c135 36 0 1.35144e-19 $X=7.13 $Y=0.85
c136 28 0 2.95874e-19 $X=6.985 $Y=0.85
c137 1 0 9.39349e-20 $X=3.865 $Y=1.145
r138 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r139 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r140 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r141 28 29 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=4.055 $Y2=0.85
r142 26 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=0.98 $X2=3.775 $Y2=0.98
r143 26 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r144 25 36 5.12197 $w=2.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.01 $Y=0.87
+ $X2=7.13 $Y2=0.87
r145 23 43 44.8475 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=0.98
+ $X2=6.845 $Y2=1.145
r146 23 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.845 $Y=0.98
+ $X2=6.845 $Y2=0.815
r147 22 25 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0.9
+ $X2=7.01 $Y2=0.9
r148 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.845
+ $Y=0.98 $X2=6.845 $Y2=0.98
r149 17 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.905 $Y=2.275
+ $X2=6.905 $Y2=1.685
r150 14 19 37.1127 $w=1.7e-07 $l=8.5e-08 $layer=POLY_cond $X=6.895 $Y=1.6
+ $X2=6.895 $Y2=1.685
r151 14 43 192.377 $w=1.7e-07 $l=4.55e-07 $layer=POLY_cond $X=6.895 $Y=1.6
+ $X2=6.895 $Y2=1.145
r152 11 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.785 $Y=0.445
+ $X2=6.785 $Y2=0.815
r153 5 39 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.81 $Y2=0.98
r154 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.905 $Y2=0.445
r155 1 39 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.81 $Y2=0.98
r156 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.865 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_476_47# 1 2 7 9 11 14 16 20 22 24 25 26 30
+ 35 37 38 43 44 53
c157 53 0 1.95729e-19 $X=4.705 $Y=1.4
c158 43 0 4.43992e-20 $X=3.44 $Y=1.3
c159 26 0 1.01003e-19 $X=3.02 $Y=2.335
c160 22 0 3.64688e-20 $X=5.205 $Y=0.735
c161 16 0 1.15925e-19 $X=5.13 $Y=0.825
c162 7 0 3.12358e-20 $X=4.265 $Y=0.735
r163 48 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.705 $Y2=1.4
r164 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.265 $Y2=1.4
r165 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.4 $X2=4.285 $Y2=1.4
r166 44 47 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.245 $Y=1.32
+ $X2=4.245 $Y2=1.4
r167 42 43 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=1.3
+ $X2=3.44 $Y2=1.3
r168 40 42 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.105 $Y=1.3
+ $X2=3.355 $Y2=1.3
r169 38 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=4.245 $Y2=1.32
r170 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=3.44 $Y2=1.32
r171 37 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.195
+ $X2=3.355 $Y2=1.3
r172 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.355 $Y=0.465
+ $X2=3.355 $Y2=1.195
r173 34 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=1.3
r174 34 35 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=2.25
r175 30 36 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=3.355 $Y2=0.465
r176 30 32 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=2.59 $Y2=0.365
r177 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.105 $Y2=2.25
r178 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=2.525 $Y2=2.335
r179 22 24 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=0.735
+ $X2=5.205 $Y2=0.445
r180 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=1.4
r181 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=2.275
r182 17 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=0.825
+ $X2=4.265 $Y2=0.825
r183 16 22 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=5.205 $Y2=0.735
r184 16 17 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=4.34 $Y2=0.825
r185 12 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=1.4
r186 12 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=2.275
r187 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.235
+ $X2=4.265 $Y2=1.4
r188 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=0.825
r189 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=1.235
r190 7 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.825
r191 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.445
r192 2 28 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.065 $X2=2.525 $Y2=2.335
r193 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_1178_261# 1 2 9 13 18 21 25 29 32 34 35 40
c79 34 0 1.80017e-19 $X=7.51 $Y=1.67
c80 18 0 6.36135e-20 $X=6.425 $Y=1.38
r81 38 40 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.615 $Y=0.515
+ $X2=7.785 $Y2=0.515
r82 33 35 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.785 $Y2=1.67
r83 33 34 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.51 $Y2=1.67
r84 32 35 0.716491 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=7.785 $Y=1.575
+ $X2=7.785 $Y2=1.67
r85 31 40 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.785 $Y=0.68
+ $X2=7.785 $Y2=0.515
r86 31 32 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=7.785 $Y=0.68
+ $X2=7.785 $Y2=1.575
r87 27 33 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.67
r88 27 29 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.87
r89 24 34 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=6.075 $Y=1.66
+ $X2=7.51 $Y2=1.66
r90 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.075
+ $Y=1.66 $X2=6.075 $Y2=1.66
r91 20 25 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=6.05 $Y=1.665
+ $X2=6.05 $Y2=1.66
r92 20 21 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=6.05 $Y=1.665
+ $X2=6.05 $Y2=1.825
r93 16 25 36.9668 $w=3.2e-07 $l=2.05e-07 $layer=POLY_cond $X=6.05 $Y=1.455
+ $X2=6.05 $Y2=1.66
r94 16 18 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=6.05 $Y=1.38
+ $X2=6.425 $Y2=1.38
r95 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.425 $Y=1.305
+ $X2=6.425 $Y2=1.38
r96 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.425 $Y=1.305
+ $X2=6.425 $Y2=0.445
r97 9 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.965 $Y=2.275
+ $X2=5.965 $Y2=1.825
r98 2 29 300 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=2 $X=7.455
+ $Y=1.645 $X2=7.595 $Y2=1.87
r99 1 38 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.48
+ $Y=0.235 $X2=7.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_1028_413# 1 2 3 12 16 18 19 22 24 26 27 28
+ 33 34 38 39 40 43 48 50 53 55 57
c159 33 0 7.39505e-20 $X=5.655 $Y=1.915
c160 28 0 1.39518e-19 $X=5.57 $Y=2.29
c161 22 0 1.25086e-19 $X=8.345 $Y=0.56
r162 60 61 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=7.38 $Y=1.26
+ $X2=7.405 $Y2=1.26
r163 56 60 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=7.325 $Y=1.26
+ $X2=7.38 $Y2=1.26
r164 55 57 10.0774 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.325 $Y=1.29
+ $X2=7.14 $Y2=1.29
r165 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.325
+ $Y=1.26 $X2=7.325 $Y2=1.26
r166 46 48 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=2.085
+ $X2=6.66 $Y2=2.21
r167 45 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=6.405 $Y2=1.32
r168 45 57 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=7.14 $Y2=1.32
r169 43 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.235
+ $X2=6.405 $Y2=1.32
r170 42 43 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.405 $Y=0.475
+ $X2=6.405 $Y2=1.235
r171 41 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.74 $Y=2 $X2=5.655
+ $Y2=2
r172 40 46 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.54 $Y=2
+ $X2=6.66 $Y2=2.085
r173 40 41 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.54 $Y=2 $X2=5.74
+ $Y2=2
r174 38 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=6.405 $Y2=1.32
r175 38 39 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=5.74 $Y2=1.32
r176 34 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=6.405 $Y2=0.475
r177 34 36 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=5.805 $Y2=0.39
r178 33 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=1.915
+ $X2=5.655 $Y2=2
r179 32 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.655 $Y=1.405
+ $X2=5.74 $Y2=1.32
r180 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.655 $Y=1.405
+ $X2=5.655 $Y2=1.915
r181 28 50 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.655 $Y=2.29
+ $X2=5.655 $Y2=2
r182 28 30 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.57 $Y=2.29
+ $X2=5.275 $Y2=2.29
r183 24 27 35.9208 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=8.345 $Y=1.41
+ $X2=8.345 $Y2=1.252
r184 24 26 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.345 $Y=1.41
+ $X2=8.345 $Y2=1.985
r185 20 27 35.9208 $w=1.5e-07 $l=1.57e-07 $layer=POLY_cond $X=8.345 $Y=1.095
+ $X2=8.345 $Y2=1.252
r186 20 22 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=8.345 $Y=1.095
+ $X2=8.345 $Y2=0.56
r187 19 61 11.0213 $w=3.28e-07 $l=7.88987e-08 $layer=POLY_cond $X=7.48 $Y=1.252
+ $X2=7.405 $Y2=1.26
r188 18 27 4.4846 $w=3.15e-07 $l=7.5e-08 $layer=POLY_cond $X=8.27 $Y=1.252
+ $X2=8.345 $Y2=1.252
r189 18 19 144.719 $w=3.15e-07 $l=7.9e-07 $layer=POLY_cond $X=8.27 $Y=1.252
+ $X2=7.48 $Y2=1.252
r190 14 61 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.405 $Y=1.095
+ $X2=7.405 $Y2=1.26
r191 14 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.405 $Y=1.095
+ $X2=7.405 $Y2=0.505
r192 10 60 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.38 $Y=1.425
+ $X2=7.38 $Y2=1.26
r193 10 12 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.38 $Y=1.425
+ $X2=7.38 $Y2=2.065
r194 3 48 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.065 $X2=6.695 $Y2=2.21
r195 2 30 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=2.065 $X2=5.275 $Y2=2.33
r196 1 36 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.805 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_1602_47# 1 2 7 9 12 14 16 19 25 30 33 37
+ 39 42
c75 42 0 1.91378e-19 $X=9.185 $Y=1.16
r76 37 38 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.135 $Y=2 $X2=8.135
+ $Y2=1.915
r77 34 42 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=8.765 $Y=1.16
+ $X2=9.185 $Y2=1.16
r78 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.765
+ $Y=1.16 $X2=8.765 $Y2=1.16
r79 31 39 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.3 $Y=1.16
+ $X2=8.175 $Y2=1.16
r80 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.3 $Y=1.16
+ $X2=8.765 $Y2=1.16
r81 30 38 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.175 $Y=1.66
+ $X2=8.175 $Y2=1.915
r82 27 39 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=8.175 $Y=1.325
+ $X2=8.175 $Y2=1.16
r83 27 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.175 $Y=1.325
+ $X2=8.175 $Y2=1.66
r84 23 39 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=8.135 $Y=0.995
+ $X2=8.175 $Y2=1.16
r85 23 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.135 $Y=0.995
+ $X2=8.135 $Y2=0.51
r86 17 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.185 $Y=1.325
+ $X2=9.185 $Y2=1.16
r87 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.185 $Y=1.325
+ $X2=9.185 $Y2=1.985
r88 14 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.185 $Y=0.995
+ $X2=9.185 $Y2=1.16
r89 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.185 $Y=0.995
+ $X2=9.185 $Y2=0.56
r90 10 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.16
r91 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.765 $Y=1.325
+ $X2=8.765 $Y2=1.985
r92 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=1.16
r93 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.765 $Y=0.995
+ $X2=8.765 $Y2=0.56
r94 2 37 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=8.01
+ $Y=1.485 $X2=8.135 $Y2=2
r95 2 30 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.01
+ $Y=1.485 $X2=8.135 $Y2=1.66
r96 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.01
+ $Y=0.235 $X2=8.135 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49 51
+ 53 55 57 63 68 73 81 86 91 97 100 103 110 113 120 123 127
c171 127 0 2.99957e-19 $X=9.43 $Y=2.72
c172 45 0 1.91378e-19 $X=8.555 $Y=1.66
r173 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r174 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r175 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r176 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r177 113 116 10.4269 $w=4.18e-07 $l=3.8e-07 $layer=LI1_cond $X=6.13 $Y=2.34
+ $X2=6.13 $Y2=2.72
r178 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r179 107 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r180 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r181 103 106 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.62 $Y=2.34
+ $X2=3.62 $Y2=2.72
r182 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r183 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 95 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r185 95 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r186 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r187 92 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.64 $Y=2.72
+ $X2=8.555 $Y2=2.72
r188 92 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.64 $Y=2.72
+ $X2=8.97 $Y2=2.72
r189 91 126 4.18617 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.31 $Y=2.72
+ $X2=9.485 $Y2=2.72
r190 91 94 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.31 $Y=2.72
+ $X2=8.97 $Y2=2.72
r191 90 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r192 90 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r193 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r194 87 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.175 $Y2=2.72
r195 87 89 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.59 $Y2=2.72
r196 86 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=2.72
+ $X2=8.555 $Y2=2.72
r197 86 89 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=8.47 $Y=2.72
+ $X2=7.59 $Y2=2.72
r198 85 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r199 85 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r200 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r201 82 116 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.13 $Y2=2.72
r202 82 84 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.67 $Y2=2.72
r203 81 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.175 $Y2=2.72
r204 81 84 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r205 80 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r206 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r207 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r208 77 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r209 76 79 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r210 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r211 74 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.495 $Y2=2.72
r212 74 76 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.83 $Y2=2.72
r213 73 116 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.13 $Y2=2.72
r214 73 79 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.75 $Y2=2.72
r215 72 107 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r216 72 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r217 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r218 69 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r219 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r220 68 106 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=3.62 $Y2=2.72
r221 68 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=2.07 $Y2=2.72
r222 67 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r223 67 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r224 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r225 64 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r226 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r227 63 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r228 63 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r229 57 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r230 55 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r231 53 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r232 53 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r233 49 126 3.06189 $w=2.65e-07 $l=1.04307e-07 $layer=LI1_cond $X=9.442 $Y=2.635
+ $X2=9.485 $Y2=2.72
r234 49 51 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=9.442 $Y=2.635
+ $X2=9.442 $Y2=1.955
r235 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.555 $Y=1.66
+ $X2=8.555 $Y2=2.34
r236 43 123 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=2.635
+ $X2=8.555 $Y2=2.72
r237 43 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.555 $Y=2.635
+ $X2=8.555 $Y2=2.34
r238 39 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.72
r239 39 41 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.21
r240 35 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.72
r241 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.34
r242 34 106 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.62 $Y2=2.72
r243 33 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=4.495 $Y2=2.72
r244 33 34 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.81 $Y2=2.72
r245 29 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r246 29 31 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.22
r247 25 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r248 25 27 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r249 8 51 300 $w=1.7e-07 $l=5.33245e-07 $layer=licon1_PDIFF $count=2 $X=9.26
+ $Y=1.485 $X2=9.395 $Y2=1.955
r250 7 48 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.42
+ $Y=1.485 $X2=8.555 $Y2=2.34
r251 7 45 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.42
+ $Y=1.485 $X2=8.555 $Y2=1.66
r252 6 41 600 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.065 $X2=7.17 $Y2=2.21
r253 5 113 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=2.065 $X2=6.175 $Y2=2.34
r254 4 37 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.065 $X2=4.495 $Y2=2.34
r255 3 103 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.065 $X2=3.595 $Y2=2.34
r256 2 31 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.645 $X2=1.62 $Y2=2.22
r257 1 27 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%A_381_47# 1 2 8 9 10 11 12 15 20
c60 20 0 1.34441e-19 $X=2.04 $Y=1.96
r61 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r62 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.88
r63 11 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.6 $Y2=1.88
r64 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r65 9 10 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.6 $Y2=0.73
r66 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.795
+ $X2=1.6 $Y2=1.88
r67 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.6 $Y2=0.73
r68 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.515 $Y2=1.795
r69 2 20 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.645 $X2=2.04 $Y2=1.96
r70 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%Q 1 2 7 8 9 10 11 12 27 29 37 45
c32 10 0 1.25086e-19 $X=9.345 $Y=0.765
r33 37 45 1.08705 $w=6.34e-07 $l=8.45577e-08 $layer=LI1_cond $X=9.297 $Y=0.895
+ $X2=9.232 $Y2=0.85
r34 27 29 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.975 $Y=1.615
+ $X2=8.975 $Y2=1.66
r35 21 26 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=9.012 $Y=0.765
+ $X2=9.012 $Y2=0.63
r36 12 27 5.02651 $w=7.16e-07 $l=2.55996e-07 $layer=LI1_cond $X=9.192 $Y=1.53
+ $X2=8.975 $Y2=1.615
r37 11 12 4.89445 $w=7.23e-07 $l=2.55e-07 $layer=LI1_cond $X=9.297 $Y=1.19
+ $X2=9.297 $Y2=1.445
r38 10 45 0.384858 $w=6.34e-07 $l=2e-08 $layer=LI1_cond $X=9.232 $Y=0.83
+ $X2=9.232 $Y2=0.85
r39 10 21 6.02774 $w=6.34e-07 $l=2.504e-07 $layer=LI1_cond $X=9.232 $Y=0.83
+ $X2=9.012 $Y2=0.765
r40 10 11 5.92651 $w=5.53e-07 $l=2.75e-07 $layer=LI1_cond $X=9.297 $Y=0.915
+ $X2=9.297 $Y2=1.19
r41 10 37 0.431019 $w=5.53e-07 $l=2e-08 $layer=LI1_cond $X=9.297 $Y=0.915
+ $X2=9.297 $Y2=0.895
r42 9 35 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=8.975 $Y=2.21
+ $X2=8.975 $Y2=2.34
r43 8 9 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.975 $Y=1.87
+ $X2=8.975 $Y2=2.21
r44 8 29 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8.975 $Y=1.87
+ $X2=8.975 $Y2=1.66
r45 7 26 5.64462 $w=2.43e-07 $l=1.2e-07 $layer=LI1_cond $X=9.012 $Y=0.51
+ $X2=9.012 $Y2=0.63
r46 2 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.485 $X2=8.975 $Y2=2.34
r47 2 29 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.84
+ $Y=1.485 $X2=8.975 $Y2=1.66
r48 1 26 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=8.84
+ $Y=0.235 $X2=8.975 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_2%VGND 1 2 3 4 5 6 7 24 28 32 34 38 42 44 46
+ 48 50 52 58 63 71 79 84 90 93 96 99 103 109 113
c156 113 0 2.71124e-20 $X=9.43 $Y=0
c157 79 0 1.35144e-19 $X=8.39 $Y=0
r158 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r159 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r160 103 106 8.97059 $w=6.38e-07 $l=4.8e-07 $layer=LI1_cond $X=7.01 $Y=0
+ $X2=7.01 $Y2=0.48
r161 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r162 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r163 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r164 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r165 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r166 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r167 88 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r168 88 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.51 $Y2=0
r169 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r170 85 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.72 $Y=0
+ $X2=8.555 $Y2=0
r171 85 87 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.72 $Y=0 $X2=8.97
+ $Y2=0
r172 84 112 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=9.482 $Y2=0
r173 84 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=8.97 $Y2=0
r174 83 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r175 83 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.13 $Y2=0
r176 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r177 80 103 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=7.33 $Y=0 $X2=7.01
+ $Y2=0
r178 80 82 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.33 $Y=0 $X2=8.05
+ $Y2=0
r179 79 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.39 $Y=0
+ $X2=8.555 $Y2=0
r180 79 82 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.39 $Y=0 $X2=8.05
+ $Y2=0
r181 78 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r182 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r183 75 78 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r184 75 100 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r185 74 77 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0 $X2=6.67
+ $Y2=0
r186 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r187 72 99 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.92
+ $Y2=0
r188 72 74 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.29
+ $Y2=0
r189 71 103 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=6.69 $Y=0 $X2=7.01
+ $Y2=0
r190 71 77 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.69 $Y=0 $X2=6.67
+ $Y2=0
r191 70 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r192 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r193 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r194 67 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r195 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r196 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r197 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r198 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r199 63 96 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.815
+ $Y2=0
r200 63 69 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.45
+ $Y2=0
r201 62 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r202 62 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r203 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r204 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r205 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r206 58 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r207 58 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r208 52 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r209 50 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r210 48 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r211 48 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r212 44 112 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.482 $Y2=0
r213 44 46 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.44 $Y2=0.38
r214 40 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=0.085
+ $X2=8.555 $Y2=0
r215 40 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.555 $Y=0.085
+ $X2=8.555 $Y2=0.38
r216 36 99 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.92 $Y=0.085
+ $X2=4.92 $Y2=0
r217 36 38 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=4.92 $Y=0.085
+ $X2=4.92 $Y2=0.38
r218 35 96 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=3.815
+ $Y2=0
r219 34 99 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.92
+ $Y2=0
r220 34 35 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.76 $Y=0 $X2=4.02
+ $Y2=0
r221 30 96 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r222 30 32 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.36
r223 26 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r224 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r225 22 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r226 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r227 7 46 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.26
+ $Y=0.235 $X2=9.395 $Y2=0.38
r228 6 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.42
+ $Y=0.235 $X2=8.555 $Y2=0.38
r229 5 106 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.86
+ $Y=0.235 $X2=7.095 $Y2=0.48
r230 4 38 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=4.995 $Y2=0.38
r231 3 32 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.695 $Y2=0.36
r232 2 28 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r233 1 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__ebufn_1.spice
* Created: Tue Sep  1 19:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__ebufn_1.pex.spice"
.subckt sky130_fd_sc_hd__ebufn_1  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.098125 AS=0.1092 PD=1.005 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_193_369#_M1007_d N_TE_B_M1007_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.2583 AS=0.098125 PD=2.07 PS=1.005 NRD=94.284 NRS=51.036 M=1 R=2.8
+ SA=75000.4 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1002 A_531_47# N_A_193_369#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.2275 PD=0.86 PS=2 NRD=9.228 NRS=15.684 M=1 R=4.33333
+ SA=75000.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Z_M1006_d N_A_27_47#_M1006_g A_531_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.286 AS=0.06825 PD=2.18 PS=0.86 NRD=24.912 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_193_369#_M1001_d N_TE_B_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 A_383_297# N_TE_B_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1 AD=0.475
+ AS=0.27 PD=1.95 PS=2.54 NRD=82.7203 NRS=0.9653 M=1 R=6.66667 SA=75000.2
+ SB=75001.3 A=0.15 P=2.3 MULT=1
MM1000 N_Z_M1000_d N_A_27_47#_M1000_g A_383_297# VPB PHIGHVT L=0.15 W=1 AD=0.315
+ AS=0.475 PD=2.63 PS=1.95 NRD=9.8303 NRS=82.7203 M=1 R=6.66667 SA=75001.3
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__ebufn_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nor4bb_4.spice.pex
* Created: Thu Aug 27 14:33:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%C_N 1 3 6 8 14 17
c25 6 0 1.25275e-19 $X=0.49 $Y=1.985
c26 1 0 1.26352e-19 $X=0.49 $Y=0.995
r27 11 14 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.28 $Y=1.16
+ $X2=0.49 $Y2=1.16
r28 8 17 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.22 $X2=0.23
+ $Y2=1.22
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.28
+ $Y=1.16 $X2=0.28 $Y2=1.16
r30 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r31 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r32 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r33 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%D_N 1 3 6 8 13 18
r39 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.16 $X2=1.12 $Y2=1.16
r40 10 13 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.12 $Y2=1.16
r41 8 18 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=1.155 $Y=1.2 $X2=1.12
+ $Y2=1.2
r42 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r43 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325 $X2=0.91
+ $Y2=1.985
r44 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995 $X2=0.91
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A_197_47# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 37 39 43 44 46 48 54 57 64
c124 44 0 1.26352e-19 $X=1.285 $Y=0.82
c125 39 0 1.25275e-19 $X=1.465 $Y=1.62
r126 63 64 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.73 $Y=1.16
+ $X2=3.15 $Y2=1.16
r127 55 63 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.68 $Y=1.16 $X2=2.73
+ $Y2=1.16
r128 55 61 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.68 $Y=1.16
+ $X2=2.31 $Y2=1.16
r129 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.16 $X2=2.68 $Y2=1.16
r130 52 61 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=2 $Y=1.16 $X2=2.31
+ $Y2=1.16
r131 52 58 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2 $Y=1.16 $X2=1.89
+ $Y2=1.16
r132 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2 $Y=1.16 $X2=2.68
+ $Y2=1.16
r133 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2
+ $Y=1.16 $X2=2 $Y2=1.16
r134 49 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=1.16
+ $X2=1.55 $Y2=1.16
r135 49 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.635 $Y=1.16
+ $X2=2 $Y2=1.16
r136 47 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.245
+ $X2=1.55 $Y2=1.16
r137 47 48 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=1.245
+ $X2=1.55 $Y2=1.535
r138 46 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=1.075
+ $X2=1.55 $Y2=1.16
r139 45 46 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.55 $Y=0.905
+ $X2=1.55 $Y2=1.075
r140 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.465 $Y=0.82
+ $X2=1.55 $Y2=0.905
r141 43 44 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.465 $Y=0.82
+ $X2=1.285 $Y2=0.82
r142 39 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.465 $Y=1.62
+ $X2=1.55 $Y2=1.535
r143 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.465 $Y=1.62
+ $X2=1.12 $Y2=1.62
r144 35 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.12 $Y=0.735
+ $X2=1.285 $Y2=0.82
r145 35 37 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.12 $Y=0.735
+ $X2=1.12 $Y2=0.39
r146 31 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.16
r147 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=1.325
+ $X2=3.15 $Y2=1.985
r148 28 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=1.16
r149 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.15 $Y=0.995
+ $X2=3.15 $Y2=0.56
r150 24 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.16
r151 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.985
r152 21 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=0.995
+ $X2=2.73 $Y2=1.16
r153 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.73 $Y=0.995
+ $X2=2.73 $Y2=0.56
r154 17 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.325
+ $X2=2.31 $Y2=1.16
r155 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.31 $Y=1.325
+ $X2=2.31 $Y2=1.985
r156 14 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=0.995
+ $X2=2.31 $Y2=1.16
r157 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.31 $Y=0.995
+ $X2=2.31 $Y2=0.56
r158 10 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=1.16
r159 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.89 $Y=1.325
+ $X2=1.89 $Y2=1.985
r160 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.89 $Y2=1.16
r161 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.89 $Y=0.995
+ $X2=1.89 $Y2=0.56
r162 2 41 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.62
r163 1 37 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A_27_297# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 37 41 44 45 48 49 54 59 66 73
c144 48 0 1.12286e-19 $X=3.44 $Y=1.875
r145 70 71 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.99 $Y=1.16
+ $X2=4.41 $Y2=1.16
r146 65 66 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.79
+ $X2=0.785 $Y2=1.79
r147 64 65 9.85006 $w=5.08e-07 $l=4.2e-07 $layer=LI1_cond $X=0.28 $Y=1.79
+ $X2=0.7 $Y2=1.79
r148 61 64 1.28989 $w=5.08e-07 $l=5.5e-08 $layer=LI1_cond $X=0.225 $Y=1.79
+ $X2=0.28 $Y2=1.79
r149 55 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.74 $Y=1.16 $X2=4.83
+ $Y2=1.16
r150 55 71 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.74 $Y=1.16
+ $X2=4.41 $Y2=1.16
r151 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.74
+ $Y=1.16 $X2=4.74 $Y2=1.16
r152 52 70 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.72 $Y=1.16
+ $X2=3.99 $Y2=1.16
r153 52 67 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.72 $Y=1.16
+ $X2=3.57 $Y2=1.16
r154 51 54 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=3.72 $Y=1.18
+ $X2=4.74 $Y2=1.18
r155 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.72
+ $Y=1.16 $X2=3.72 $Y2=1.16
r156 49 51 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=3.525 $Y=1.18
+ $X2=3.72 $Y2=1.18
r157 47 49 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.44 $Y=1.285
+ $X2=3.525 $Y2=1.18
r158 47 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.44 $Y=1.285
+ $X2=3.44 $Y2=1.875
r159 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.355 $Y=1.96
+ $X2=3.44 $Y2=1.875
r160 45 66 167.668 $w=1.68e-07 $l=2.57e-06 $layer=LI1_cond $X=3.355 $Y=1.96
+ $X2=0.785 $Y2=1.96
r161 44 65 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.7 $Y=1.535
+ $X2=0.7 $Y2=1.79
r162 43 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.895
+ $X2=0.7 $Y2=0.81
r163 43 44 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.7 $Y=0.895 $X2=0.7
+ $Y2=1.535
r164 39 61 4.24724 $w=2.8e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=1.79
r165 39 41 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=2.3
r166 35 59 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.265 $Y=0.81
+ $X2=0.7 $Y2=0.81
r167 35 37 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.265 $Y=0.725
+ $X2=0.265 $Y2=0.39
r168 31 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.83 $Y=1.325
+ $X2=4.83 $Y2=1.16
r169 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.83 $Y=1.325
+ $X2=4.83 $Y2=1.985
r170 28 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.83 $Y=0.995
+ $X2=4.83 $Y2=1.16
r171 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.83 $Y=0.995
+ $X2=4.83 $Y2=0.56
r172 24 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.325
+ $X2=4.41 $Y2=1.16
r173 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.41 $Y=1.325
+ $X2=4.41 $Y2=1.985
r174 21 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=0.995
+ $X2=4.41 $Y2=1.16
r175 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.41 $Y=0.995
+ $X2=4.41 $Y2=0.56
r176 17 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.16
r177 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.99 $Y=1.325
+ $X2=3.99 $Y2=1.985
r178 14 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=1.16
r179 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.99 $Y=0.995
+ $X2=3.99 $Y2=0.56
r180 10 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.16
r181 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.57 $Y=1.325
+ $X2=3.57 $Y2=1.985
r182 7 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=1.16
r183 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.57 $Y=0.995
+ $X2=3.57 $Y2=0.56
r184 2 64 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r185 2 41 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r186 1 37 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%B 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r78 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.94 $Y=1.16 $X2=7.03
+ $Y2=1.16
r79 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.94
+ $Y=1.16 $X2=6.94 $Y2=1.16
r80 37 39 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.61 $Y=1.16
+ $X2=6.94 $Y2=1.16
r81 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.19 $Y=1.16
+ $X2=6.61 $Y2=1.16
r82 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.92 $Y=1.16
+ $X2=6.19 $Y2=1.16
r83 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.92
+ $Y=1.16 $X2=5.92 $Y2=1.16
r84 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.77 $Y=1.16
+ $X2=5.92 $Y2=1.16
r85 29 40 38.8182 $w=2.08e-07 $l=7.35e-07 $layer=LI1_cond $X=6.205 $Y=1.18
+ $X2=6.94 $Y2=1.18
r86 29 35 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=6.205 $Y=1.18
+ $X2=5.92 $Y2=1.18
r87 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.03 $Y=1.325
+ $X2=7.03 $Y2=1.16
r88 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.03 $Y=1.325
+ $X2=7.03 $Y2=1.985
r89 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.03 $Y=0.995
+ $X2=7.03 $Y2=1.16
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.03 $Y=0.995
+ $X2=7.03 $Y2=0.56
r91 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.61 $Y=1.325
+ $X2=6.61 $Y2=1.16
r92 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.61 $Y=1.325
+ $X2=6.61 $Y2=1.985
r93 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.61 $Y=0.995
+ $X2=6.61 $Y2=1.16
r94 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.61 $Y=0.995
+ $X2=6.61 $Y2=0.56
r95 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.19 $Y=1.325
+ $X2=6.19 $Y2=1.16
r96 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.19 $Y=1.325
+ $X2=6.19 $Y2=1.985
r97 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=1.16
r98 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=0.56
r99 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.77 $Y=1.325
+ $X2=5.77 $Y2=1.16
r100 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.77 $Y=1.325
+ $X2=5.77 $Y2=1.985
r101 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=1.16
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 40 41
r71 39 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.62 $Y=1.16 $X2=8.71
+ $Y2=1.16
r72 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.62
+ $Y=1.16 $X2=8.62 $Y2=1.16
r73 37 39 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=8.29 $Y=1.16
+ $X2=8.62 $Y2=1.16
r74 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.87 $Y=1.16
+ $X2=8.29 $Y2=1.16
r75 34 36 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.6 $Y=1.16 $X2=7.87
+ $Y2=1.16
r76 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.6 $Y=1.16
+ $X2=7.6 $Y2=1.16
r77 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.45 $Y=1.16 $X2=7.6
+ $Y2=1.16
r78 29 40 30.368 $w=2.08e-07 $l=5.75e-07 $layer=LI1_cond $X=8.045 $Y=1.18
+ $X2=8.62 $Y2=1.18
r79 29 35 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=8.045 $Y=1.18
+ $X2=7.6 $Y2=1.18
r80 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=1.325
+ $X2=8.71 $Y2=1.16
r81 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.71 $Y=1.325
+ $X2=8.71 $Y2=1.985
r82 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=0.995
+ $X2=8.71 $Y2=1.16
r83 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.71 $Y=0.995
+ $X2=8.71 $Y2=0.56
r84 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.29 $Y=1.325
+ $X2=8.29 $Y2=1.16
r85 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.29 $Y=1.325
+ $X2=8.29 $Y2=1.985
r86 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.29 $Y=0.995
+ $X2=8.29 $Y2=1.16
r87 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.29 $Y=0.995
+ $X2=8.29 $Y2=0.56
r88 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.87 $Y=1.325
+ $X2=7.87 $Y2=1.16
r89 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.87 $Y=1.325
+ $X2=7.87 $Y2=1.985
r90 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.87 $Y=0.995
+ $X2=7.87 $Y2=1.16
r91 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.87 $Y=0.995
+ $X2=7.87 $Y2=0.56
r92 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=1.325
+ $X2=7.45 $Y2=1.16
r93 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.45 $Y=1.325 $X2=7.45
+ $Y2=1.985
r94 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=0.995
+ $X2=7.45 $Y2=1.16
r95 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.45 $Y=0.995 $X2=7.45
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%VPWR 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r106 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r107 48 49 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r108 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r109 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r110 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r111 39 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.625 $Y=2.72
+ $X2=8.5 $Y2=2.72
r112 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.625 $Y=2.72
+ $X2=8.97 $Y2=2.72
r113 38 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r114 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=7.59 $Y2=2.72
r115 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r116 35 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.785 $Y=2.72
+ $X2=7.66 $Y2=2.72
r117 35 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.785 $Y=2.72
+ $X2=8.05 $Y2=2.72
r118 34 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.5 $Y2=2.72
r119 34 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.375 $Y=2.72
+ $X2=8.05 $Y2=2.72
r120 33 49 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 32 33 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r123 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.7 $Y2=2.72
r124 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=1.15 $Y2=2.72
r125 29 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.535 $Y=2.72
+ $X2=7.66 $Y2=2.72
r126 29 32 416.561 $w=1.68e-07 $l=6.385e-06 $layer=LI1_cond $X=7.535 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.7 $Y2=2.72
r128 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r129 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r131 18 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=2.635
+ $X2=8.5 $Y2=2.72
r132 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.5 $Y=2.635
+ $X2=8.5 $Y2=1.96
r133 14 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.66 $Y=2.635
+ $X2=7.66 $Y2=2.72
r134 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.66 $Y=2.635
+ $X2=7.66 $Y2=1.96
r135 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=2.635 $X2=0.7
+ $Y2=2.72
r136 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.7 $Y=2.635
+ $X2=0.7 $Y2=2.3
r137 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.365
+ $Y=1.485 $X2=8.5 $Y2=1.96
r138 2 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.525
+ $Y=1.485 $X2=7.66 $Y2=1.96
r139 1 12 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A_311_297# 1 2 3 4 5 16 24 28 30 34 36 37
r49 32 34 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.055 $Y=2.295
+ $X2=5.055 $Y2=1.96
r50 31 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.325 $Y=2.38
+ $X2=4.2 $Y2=2.38
r51 30 32 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.915 $Y=2.38
+ $X2=5.055 $Y2=2.295
r52 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.915 $Y=2.38
+ $X2=4.325 $Y2=2.38
r53 26 37 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=2.295
+ $X2=4.2 $Y2=2.38
r54 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.2 $Y=2.295
+ $X2=4.2 $Y2=1.96
r55 24 37 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.38
+ $X2=4.2 $Y2=2.38
r56 24 36 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.075 $Y=2.38
+ $X2=3.525 $Y2=2.38
r57 21 23 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=2.52 $Y=2.34
+ $X2=3.36 $Y2=2.34
r58 18 21 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=1.68 $Y=2.34
+ $X2=2.52 $Y2=2.34
r59 16 36 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.4 $Y=2.34
+ $X2=3.525 $Y2=2.34
r60 16 23 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.4 $Y=2.34 $X2=3.36
+ $Y2=2.34
r61 5 34 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.905
+ $Y=1.485 $X2=5.04 $Y2=1.96
r62 4 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.065
+ $Y=1.485 $X2=4.2 $Y2=1.96
r63 3 23 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.485 $X2=3.36 $Y2=2.3
r64 2 21 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.485 $X2=2.52 $Y2=2.3
r65 1 18 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=1.485 $X2=1.68 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 42 43 47
+ 49 53 55 59 61 65 67 71 73 77 79 80 81 82 83 84 85 88 96
r197 90 93 33.3811 $w=2.88e-07 $l=8.4e-07 $layer=LI1_cond $X=2.1 $Y=1.56
+ $X2=2.94 $Y2=1.56
r198 88 96 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=3.015 $Y=1.56
+ $X2=2.985 $Y2=1.56
r199 85 88 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=1.56
+ $X2=3.015 $Y2=1.56
r200 85 96 1.1127 $w=2.88e-07 $l=2.8e-08 $layer=LI1_cond $X=2.957 $Y=1.56
+ $X2=2.985 $Y2=1.56
r201 85 93 0.67557 $w=2.88e-07 $l=1.7e-08 $layer=LI1_cond $X=2.957 $Y=1.56
+ $X2=2.94 $Y2=1.56
r202 75 77 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.5 $Y=0.725
+ $X2=8.5 $Y2=0.39
r203 74 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=0.815
+ $X2=7.66 $Y2=0.815
r204 73 75 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=8.335 $Y=0.815
+ $X2=8.5 $Y2=0.725
r205 73 74 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=8.335 $Y=0.815
+ $X2=7.825 $Y2=0.815
r206 69 84 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.66 $Y=0.725
+ $X2=7.66 $Y2=0.815
r207 69 71 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.66 $Y=0.725
+ $X2=7.66 $Y2=0.39
r208 68 83 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.985 $Y=0.815
+ $X2=6.82 $Y2=0.815
r209 67 84 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=0.815
+ $X2=7.66 $Y2=0.815
r210 67 68 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.495 $Y=0.815
+ $X2=6.985 $Y2=0.815
r211 63 83 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.82 $Y=0.725
+ $X2=6.82 $Y2=0.815
r212 63 65 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.82 $Y=0.725
+ $X2=6.82 $Y2=0.39
r213 62 82 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0.815
+ $X2=5.98 $Y2=0.815
r214 61 83 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.655 $Y=0.815
+ $X2=6.82 $Y2=0.815
r215 61 62 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.655 $Y=0.815
+ $X2=6.145 $Y2=0.815
r216 57 82 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.98 $Y=0.725
+ $X2=5.98 $Y2=0.815
r217 57 59 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.98 $Y=0.725
+ $X2=5.98 $Y2=0.39
r218 56 81 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=0.815
+ $X2=4.62 $Y2=0.815
r219 55 82 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0.815
+ $X2=5.98 $Y2=0.815
r220 55 56 63.4646 $w=1.78e-07 $l=1.03e-06 $layer=LI1_cond $X=5.815 $Y=0.815
+ $X2=4.785 $Y2=0.815
r221 51 81 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.62 $Y=0.725
+ $X2=4.62 $Y2=0.815
r222 51 53 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.62 $Y=0.725
+ $X2=4.62 $Y2=0.39
r223 50 80 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=0.815
+ $X2=3.78 $Y2=0.815
r224 49 81 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0.815
+ $X2=4.62 $Y2=0.815
r225 49 50 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.455 $Y=0.815
+ $X2=3.945 $Y2=0.815
r226 45 80 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.78 $Y=0.725
+ $X2=3.78 $Y2=0.815
r227 45 47 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.78 $Y=0.725
+ $X2=3.78 $Y2=0.39
r228 44 79 4.10651 $w=1.8e-07 $l=2.05e-07 $layer=LI1_cond $X=3.185 $Y=0.815
+ $X2=2.98 $Y2=0.815
r229 43 80 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0.815
+ $X2=3.78 $Y2=0.815
r230 43 44 26.4949 $w=1.78e-07 $l=4.3e-07 $layer=LI1_cond $X=3.615 $Y=0.815
+ $X2=3.185 $Y2=0.815
r231 42 85 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.1 $Y=1.415
+ $X2=3.1 $Y2=1.56
r232 41 79 2.1123 $w=1.7e-07 $l=1.58745e-07 $layer=LI1_cond $X=3.1 $Y=0.905
+ $X2=2.98 $Y2=0.815
r233 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.1 $Y=0.905
+ $X2=3.1 $Y2=1.415
r234 37 79 2.1123 $w=3.3e-07 $l=1.08167e-07 $layer=LI1_cond $X=2.94 $Y=0.725
+ $X2=2.98 $Y2=0.815
r235 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.94 $Y=0.725
+ $X2=2.94 $Y2=0.39
r236 35 79 4.10651 $w=1.8e-07 $l=2.05e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.98 $Y2=0.815
r237 35 36 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.265 $Y2=0.815
r238 31 36 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.1 $Y=0.725
+ $X2=2.265 $Y2=0.815
r239 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.1 $Y=0.725
+ $X2=2.1 $Y2=0.39
r240 10 93 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.485 $X2=2.94 $Y2=1.62
r241 9 90 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.485 $X2=2.1 $Y2=1.62
r242 8 77 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.365
+ $Y=0.235 $X2=8.5 $Y2=0.39
r243 7 71 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.525
+ $Y=0.235 $X2=7.66 $Y2=0.39
r244 6 65 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.685
+ $Y=0.235 $X2=6.82 $Y2=0.39
r245 5 59 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.845
+ $Y=0.235 $X2=5.98 $Y2=0.39
r246 4 53 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.485
+ $Y=0.235 $X2=4.62 $Y2=0.39
r247 3 47 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.645
+ $Y=0.235 $X2=3.78 $Y2=0.39
r248 2 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.805
+ $Y=0.235 $X2=2.94 $Y2=0.39
r249 1 33 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.235 $X2=2.1 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A_729_297# 1 2 3 4 15 19 23 28 30 32 34
r58 24 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.105 $Y=1.54
+ $X2=5.98 $Y2=1.54
r59 23 34 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.695 $Y=1.54
+ $X2=6.82 $Y2=1.54
r60 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.695 $Y=1.54
+ $X2=6.105 $Y2=1.54
r61 20 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.745 $Y=1.54
+ $X2=4.62 $Y2=1.54
r62 19 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.855 $Y=1.54
+ $X2=5.98 $Y2=1.54
r63 19 20 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.855 $Y=1.54
+ $X2=4.745 $Y2=1.54
r64 16 28 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.905 $Y=1.54
+ $X2=3.8 $Y2=1.54
r65 15 30 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=1.54
+ $X2=4.62 $Y2=1.54
r66 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.495 $Y=1.54
+ $X2=3.905 $Y2=1.54
r67 4 34 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.685
+ $Y=1.485 $X2=6.82 $Y2=1.62
r68 3 32 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.845
+ $Y=1.485 $X2=5.98 $Y2=1.62
r69 2 30 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=4.485
+ $Y=1.485 $X2=4.62 $Y2=1.62
r70 1 28 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=3.645
+ $Y=1.485 $X2=3.78 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%A_1087_297# 1 2 3 4 5 18 20 21 24 26 28 29
+ 30 34 36 38 40 42 48
r63 38 50 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.952 $Y=1.625
+ $X2=8.952 $Y2=1.54
r64 38 40 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=8.952 $Y=1.625
+ $X2=8.952 $Y2=2.3
r65 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.205 $Y=1.54
+ $X2=8.08 $Y2=1.54
r66 36 50 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=8.795 $Y=1.54
+ $X2=8.952 $Y2=1.54
r67 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.795 $Y=1.54
+ $X2=8.205 $Y2=1.54
r68 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.08 $Y=1.625
+ $X2=8.08 $Y2=1.54
r69 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=8.08 $Y=1.625
+ $X2=8.08 $Y2=2.3
r70 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.365 $Y=1.54
+ $X2=7.24 $Y2=1.54
r71 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.955 $Y=1.54
+ $X2=8.08 $Y2=1.54
r72 30 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.955 $Y=1.54
+ $X2=7.365 $Y2=1.54
r73 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=2.295
+ $X2=7.24 $Y2=2.38
r74 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=1.625
+ $X2=7.24 $Y2=1.54
r75 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.24 $Y=1.625
+ $X2=7.24 $Y2=2.295
r76 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.525 $Y=2.38
+ $X2=6.4 $Y2=2.38
r77 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.115 $Y=2.38
+ $X2=7.24 $Y2=2.38
r78 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.115 $Y=2.38
+ $X2=6.525 $Y2=2.38
r79 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=2.295
+ $X2=6.4 $Y2=2.38
r80 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.4 $Y=2.295
+ $X2=6.4 $Y2=1.96
r81 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.275 $Y=2.38
+ $X2=6.4 $Y2=2.38
r82 20 21 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.275 $Y=2.38
+ $X2=5.685 $Y2=2.38
r83 16 21 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=5.532 $Y=2.295
+ $X2=5.685 $Y2=2.38
r84 16 18 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=5.532 $Y=2.295
+ $X2=5.532 $Y2=1.96
r85 5 50 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=1.485 $X2=8.92 $Y2=1.62
r86 5 40 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=1.485 $X2=8.92 $Y2=2.3
r87 4 48 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.945
+ $Y=1.485 $X2=8.08 $Y2=1.62
r88 4 34 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.945
+ $Y=1.485 $X2=8.08 $Y2=2.3
r89 3 46 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.105
+ $Y=1.485 $X2=7.24 $Y2=2.3
r90 3 44 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=7.105
+ $Y=1.485 $X2=7.24 $Y2=1.62
r91 2 24 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.265
+ $Y=1.485 $X2=6.4 $Y2=1.96
r92 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=5.435
+ $Y=1.485 $X2=5.56 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__NOR4BB_4%VGND 1 2 3 4 5 6 7 8 9 10 35 37 41 45 49 53
+ 57 61 63 67 69 71 74 75 77 78 80 81 83 84 85 86 87 110 116 119 124 127 129 133
+ 135
r163 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r164 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r165 126 127 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=0.235
+ $X2=5.645 $Y2=0.235
r166 122 126 5.04596 $w=6.38e-07 $l=2.7e-07 $layer=LI1_cond $X=5.29 $Y=0.235
+ $X2=5.56 $Y2=0.235
r167 122 124 13.5939 $w=6.38e-07 $l=3.35e-07 $layer=LI1_cond $X=5.29 $Y=0.235
+ $X2=4.955 $Y2=0.235
r168 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r169 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r170 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r171 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r172 114 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r173 114 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r174 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r175 111 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.08 $Y2=0
r176 111 113 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.165 $Y=0
+ $X2=8.51 $Y2=0
r177 110 132 4.27119 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.835 $Y=0
+ $X2=9.017 $Y2=0
r178 110 113 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.835 $Y=0
+ $X2=8.51 $Y2=0
r179 109 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r180 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r181 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r182 106 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.29 $Y2=0
r183 105 127 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.21 $Y=0
+ $X2=5.645 $Y2=0
r184 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r185 102 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r186 101 124 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.955 $Y2=0
r187 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r188 98 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r189 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r190 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r191 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r192 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r193 92 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r194 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r195 89 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r196 89 91 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.765 $Y=0
+ $X2=2.07 $Y2=0
r197 87 117 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r198 87 135 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r199 85 108 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.155 $Y=0
+ $X2=7.13 $Y2=0
r200 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.155 $Y=0 $X2=7.24
+ $Y2=0
r201 83 105 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.21 $Y2=0
r202 83 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.4
+ $Y2=0
r203 82 108 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.485 $Y=0
+ $X2=7.13 $Y2=0
r204 82 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=0 $X2=6.4
+ $Y2=0
r205 80 97 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=3.91 $Y2=0
r206 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.2
+ $Y2=0
r207 79 101 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.285 $Y=0
+ $X2=4.83 $Y2=0
r208 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.2
+ $Y2=0
r209 77 94 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=2.99 $Y2=0
r210 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.36
+ $Y2=0
r211 76 97 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.91 $Y2=0
r212 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.36
+ $Y2=0
r213 74 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.435 $Y=0
+ $X2=2.07 $Y2=0
r214 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.52
+ $Y2=0
r215 73 94 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=2.99 $Y2=0
r216 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.52
+ $Y2=0
r217 69 132 3.05085 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.972 $Y=0.085
+ $X2=9.017 $Y2=0
r218 69 71 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=8.972 $Y=0.085
+ $X2=8.972 $Y2=0.39
r219 65 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.08 $Y=0.085
+ $X2=8.08 $Y2=0
r220 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.08 $Y=0.085
+ $X2=8.08 $Y2=0.39
r221 64 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=0 $X2=7.24
+ $Y2=0
r222 63 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.08
+ $Y2=0
r223 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.995 $Y=0
+ $X2=7.325 $Y2=0
r224 59 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0
r225 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0.39
r226 55 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=0.085 $X2=6.4
+ $Y2=0
r227 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.4 $Y=0.085
+ $X2=6.4 $Y2=0.39
r228 51 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=0.085 $X2=4.2
+ $Y2=0
r229 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.2 $Y=0.085
+ $X2=4.2 $Y2=0.39
r230 47 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0
r231 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.36 $Y=0.085
+ $X2=3.36 $Y2=0.39
r232 43 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.52 $Y2=0
r233 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.52 $Y=0.085
+ $X2=2.52 $Y2=0.39
r234 39 119 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0
r235 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.68 $Y=0.085
+ $X2=1.68 $Y2=0.39
r236 38 116 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r237 37 119 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.68
+ $Y2=0
r238 37 38 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.595 $Y=0
+ $X2=0.785 $Y2=0
r239 33 116 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0
r240 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.39
r241 10 71 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.785
+ $Y=0.235 $X2=8.92 $Y2=0.39
r242 9 67 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.945
+ $Y=0.235 $X2=8.08 $Y2=0.39
r243 8 61 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.105
+ $Y=0.235 $X2=7.24 $Y2=0.39
r244 7 57 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.265
+ $Y=0.235 $X2=6.4 $Y2=0.39
r245 6 126 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=4.905
+ $Y=0.235 $X2=5.56 $Y2=0.39
r246 5 53 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.235 $X2=4.2 $Y2=0.39
r247 4 49 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.36 $Y2=0.39
r248 3 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.385
+ $Y=0.235 $X2=2.52 $Y2=0.39
r249 2 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.68 $Y2=0.39
r250 1 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.39
.ends


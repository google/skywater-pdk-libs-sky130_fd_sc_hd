* File: sky130_fd_sc_hd__o21bai_4.pxi.spice
* Created: Tue Sep  1 19:22:20 2020
* 
x_PM_SKY130_FD_SC_HD__O21BAI_4%B1_N N_B1_N_M1019_g N_B1_N_M1018_g B1_N
+ N_B1_N_c_108_n N_B1_N_c_109_n N_B1_N_c_110_n PM_SKY130_FD_SC_HD__O21BAI_4%B1_N
x_PM_SKY130_FD_SC_HD__O21BAI_4%A_33_297# N_A_33_297#_M1019_d N_A_33_297#_M1018_s
+ N_A_33_297#_M1002_g N_A_33_297#_M1005_g N_A_33_297#_c_135_n
+ N_A_33_297#_M1003_g N_A_33_297#_M1020_g N_A_33_297#_c_136_n
+ N_A_33_297#_M1009_g N_A_33_297#_M1022_g N_A_33_297#_c_137_n
+ N_A_33_297#_M1024_g N_A_33_297#_c_138_n N_A_33_297#_M1025_g
+ N_A_33_297#_c_148_n N_A_33_297#_c_149_n N_A_33_297#_c_150_n
+ N_A_33_297#_c_139_n N_A_33_297#_c_140_n N_A_33_297#_c_151_n
+ N_A_33_297#_c_190_p N_A_33_297#_c_141_n N_A_33_297#_c_142_n
+ N_A_33_297#_c_143_n PM_SKY130_FD_SC_HD__O21BAI_4%A_33_297#
x_PM_SKY130_FD_SC_HD__O21BAI_4%A2 N_A2_c_230_n N_A2_M1001_g N_A2_M1010_g
+ N_A2_c_231_n N_A2_M1004_g N_A2_M1015_g N_A2_c_232_n N_A2_M1007_g N_A2_M1016_g
+ N_A2_c_233_n N_A2_M1008_g N_A2_M1021_g A2 N_A2_c_234_n N_A2_c_235_n
+ PM_SKY130_FD_SC_HD__O21BAI_4%A2
x_PM_SKY130_FD_SC_HD__O21BAI_4%A1 N_A1_c_315_n N_A1_M1006_g N_A1_M1000_g
+ N_A1_c_316_n N_A1_M1012_g N_A1_M1011_g N_A1_c_317_n N_A1_M1013_g N_A1_M1017_g
+ N_A1_c_318_n N_A1_M1014_g N_A1_M1023_g A1 A1 A1 N_A1_c_320_n
+ PM_SKY130_FD_SC_HD__O21BAI_4%A1
x_PM_SKY130_FD_SC_HD__O21BAI_4%VPWR N_VPWR_M1018_d N_VPWR_M1005_d N_VPWR_M1022_d
+ N_VPWR_M1000_s N_VPWR_M1017_s N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ VPWR N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_394_n
+ N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ PM_SKY130_FD_SC_HD__O21BAI_4%VPWR
x_PM_SKY130_FD_SC_HD__O21BAI_4%Y N_Y_M1003_d N_Y_M1024_d N_Y_M1002_s N_Y_M1020_s
+ N_Y_M1010_d N_Y_M1016_d N_Y_c_494_n N_Y_c_544_n N_Y_c_495_n N_Y_c_510_n
+ N_Y_c_548_n N_Y_c_516_n N_Y_c_496_n N_Y_c_497_n N_Y_c_498_n N_Y_c_499_n
+ N_Y_c_500_n Y N_Y_c_493_n PM_SKY130_FD_SC_HD__O21BAI_4%Y
x_PM_SKY130_FD_SC_HD__O21BAI_4%A_561_297# N_A_561_297#_M1010_s
+ N_A_561_297#_M1015_s N_A_561_297#_M1021_s N_A_561_297#_M1011_d
+ N_A_561_297#_M1023_d N_A_561_297#_c_577_n N_A_561_297#_c_584_n
+ N_A_561_297#_c_578_n N_A_561_297#_c_636_n N_A_561_297#_c_586_n
+ N_A_561_297#_c_579_n N_A_561_297#_c_615_n N_A_561_297#_c_580_n
+ N_A_561_297#_c_619_n N_A_561_297#_c_581_n N_A_561_297#_c_582_n
+ N_A_561_297#_c_599_n N_A_561_297#_c_625_n N_A_561_297#_c_583_n
+ PM_SKY130_FD_SC_HD__O21BAI_4%A_561_297#
x_PM_SKY130_FD_SC_HD__O21BAI_4%VGND N_VGND_M1019_s N_VGND_M1001_d N_VGND_M1007_d
+ N_VGND_M1006_s N_VGND_M1013_s N_VGND_c_642_n N_VGND_c_643_n N_VGND_c_644_n
+ N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n N_VGND_c_648_n N_VGND_c_649_n
+ N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n N_VGND_c_653_n N_VGND_c_654_n
+ N_VGND_c_655_n VGND N_VGND_c_656_n N_VGND_c_657_n
+ PM_SKY130_FD_SC_HD__O21BAI_4%VGND
x_PM_SKY130_FD_SC_HD__O21BAI_4%A_225_47# N_A_225_47#_M1003_s N_A_225_47#_M1009_s
+ N_A_225_47#_M1025_s N_A_225_47#_M1004_s N_A_225_47#_M1008_s
+ N_A_225_47#_M1012_d N_A_225_47#_M1014_d N_A_225_47#_c_740_n
+ N_A_225_47#_c_757_n N_A_225_47#_c_741_n N_A_225_47#_c_742_n
+ N_A_225_47#_c_765_n N_A_225_47#_c_743_n N_A_225_47#_c_773_n
+ N_A_225_47#_c_744_n N_A_225_47#_c_787_n N_A_225_47#_c_745_n
+ N_A_225_47#_c_746_n N_A_225_47#_c_747_n N_A_225_47#_c_748_n
+ N_A_225_47#_c_749_n PM_SKY130_FD_SC_HD__O21BAI_4%A_225_47#
cc_1 VNB N_B1_N_c_108_n 0.0371369f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.16
cc_2 VNB N_B1_N_c_109_n 0.0152198f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.16
cc_3 VNB N_B1_N_c_110_n 0.0249829f $X=-0.19 $Y=-0.24 $X2=0.402 $Y2=0.995
cc_4 VNB N_A_33_297#_c_135_n 0.0199049f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.18
cc_5 VNB N_A_33_297#_c_136_n 0.0160012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_33_297#_c_137_n 0.0159739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_33_297#_c_138_n 0.01577f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_33_297#_c_139_n 0.00568515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_33_297#_c_140_n 0.00292552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_33_297#_c_141_n 0.00392571f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_33_297#_c_142_n 0.00125413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_33_297#_c_143_n 0.100401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_230_n 0.016004f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB N_A2_c_231_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_A2_c_232_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.18
cc_16 VNB N_A2_c_233_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A2_c_234_n 0.00255635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_235_n 0.0621425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_315_n 0.0160112f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_20 VNB N_A1_c_316_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_21 VNB N_A1_c_317_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.18
cc_22 VNB N_A1_c_318_n 0.0214754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB A1 0.0412769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A1_c_320_n 0.0684033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_394_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.00281545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_493_n 0.00104131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_642_n 0.012648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_643_n 0.00616862f $X=-0.19 $Y=-0.24 $X2=0.39 $Y2=1.18
cc_30 VNB N_VGND_c_644_n 0.00411582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_645_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_646_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_647_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_648_n 0.0705945f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_649_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_650_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_651_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_652_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_653_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_654_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_655_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_656_n 0.0283632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_657_n 0.35892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_225_47#_c_740_n 0.00240878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_225_47#_c_741_n 0.003212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_225_47#_c_742_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_225_47#_c_743_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_225_47#_c_744_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_225_47#_c_745_n 0.0126428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_225_47#_c_746_n 0.0184392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_225_47#_c_747_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_225_47#_c_748_n 0.00384439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_225_47#_c_749_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VPB N_B1_N_M1018_g 0.0254799f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_55 VPB N_B1_N_c_108_n 0.00779392f $X=-0.19 $Y=1.305 $X2=0.39 $Y2=1.16
cc_56 VPB N_A_33_297#_M1002_g 0.0178705f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_33_297#_M1005_g 0.0181953f $X=-0.19 $Y=1.305 $X2=0.402 $Y2=0.995
cc_58 VPB N_A_33_297#_M1020_g 0.0182195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_33_297#_M1022_g 0.0220476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_33_297#_c_148_n 0.00915024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_33_297#_c_149_n 0.0308647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_33_297#_c_150_n 0.00174648f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_33_297#_c_151_n 0.00139531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_33_297#_c_143_n 0.0256762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_M1010_g 0.0220691f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_66 VPB N_A2_M1015_g 0.0181358f $X=-0.19 $Y=1.305 $X2=0.402 $Y2=0.995
cc_67 VPB N_A2_M1016_g 0.018138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A2_M1021_g 0.018815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A2_c_235_n 0.0101334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A1_M1000_g 0.0185038f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_71 VPB N_A1_M1011_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.402 $Y2=0.995
cc_72 VPB N_A1_M1017_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A1_M1023_g 0.0226386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB A1 0.060829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A1_c_320_n 0.0104055f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_395_n 0.00428776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_396_n 0.00393015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_397_n 0.00456216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_398_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_399_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_400_n 0.00454762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_401_n 0.056414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_402_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_403_n 0.0167545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_404_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_405_n 0.0265518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_394_n 0.0644246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_407_n 0.0237719f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_408_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_409_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_410_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_494_n 0.00185902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_Y_c_495_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_496_n 0.00273767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_497_n 0.00235124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_498_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_Y_c_499_n 0.00202537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_500_n 0.0023869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB Y 0.0158675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_561_297#_c_577_n 0.00480939f $X=-0.19 $Y=1.305 $X2=0.39 $Y2=1.18
cc_101 VPB N_A_561_297#_c_578_n 0.00179695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_561_297#_c_579_n 0.0036062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_561_297#_c_580_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_561_297#_c_581_n 0.00235082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_561_297#_c_582_n 0.00271811f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_561_297#_c_583_n 0.00204609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 N_B1_N_M1018_g N_A_33_297#_M1002_g 0.0206704f $X=0.52 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_B1_N_M1018_g N_A_33_297#_c_148_n 0.0014856f $X=0.52 $Y=1.985 $X2=0
+ $Y2=0
cc_109 N_B1_N_c_108_n N_A_33_297#_c_148_n 0.00574551f $X=0.39 $Y=1.16 $X2=0
+ $Y2=0
cc_110 N_B1_N_c_109_n N_A_33_297#_c_148_n 0.027113f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_111 N_B1_N_M1018_g N_A_33_297#_c_149_n 0.0101093f $X=0.52 $Y=1.985 $X2=0
+ $Y2=0
cc_112 N_B1_N_M1018_g N_A_33_297#_c_150_n 0.0113567f $X=0.52 $Y=1.985 $X2=0
+ $Y2=0
cc_113 N_B1_N_c_109_n N_A_33_297#_c_150_n 0.0054781f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_N_c_110_n N_A_33_297#_c_139_n 0.00511079f $X=0.402 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_B1_N_c_110_n N_A_33_297#_c_140_n 0.00531722f $X=0.402 $Y=0.995 $X2=0
+ $Y2=0
cc_116 N_B1_N_c_108_n N_A_33_297#_c_151_n 0.00366701f $X=0.39 $Y=1.16 $X2=0
+ $Y2=0
cc_117 N_B1_N_c_110_n N_A_33_297#_c_141_n 0.0027391f $X=0.402 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_B1_N_c_108_n N_A_33_297#_c_142_n 0.0016466f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_N_c_109_n N_A_33_297#_c_142_n 0.0180619f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_N_c_108_n N_A_33_297#_c_143_n 0.0206704f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B1_N_M1018_g N_VPWR_c_395_n 0.00274642f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_N_M1018_g N_VPWR_c_394_n 0.0105294f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_N_M1018_g N_VPWR_c_407_n 0.0054256f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_N_c_108_n N_VGND_c_643_n 0.00429275f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B1_N_c_109_n N_VGND_c_643_n 0.0131644f $X=0.39 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B1_N_c_110_n N_VGND_c_643_n 0.00460417f $X=0.402 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_N_c_110_n N_VGND_c_648_n 0.00542757f $X=0.402 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_N_c_110_n N_VGND_c_657_n 0.0118287f $X=0.402 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_33_297#_c_138_n N_A2_c_230_n 0.014323f $X=2.72 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_33_297#_c_143_n N_A2_c_234_n 2.06878e-19 $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_33_297#_c_143_n N_A2_c_235_n 0.014323f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_33_297#_c_150_n N_VPWR_M1018_d 0.00168387f $X=0.725 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_33_297#_M1002_g N_VPWR_c_395_n 0.00155565f $X=0.94 $Y=1.985 $X2=0
+ $Y2=0
cc_134 N_A_33_297#_c_150_n N_VPWR_c_395_n 0.0133861f $X=0.725 $Y=1.54 $X2=0
+ $Y2=0
cc_135 N_A_33_297#_M1005_g N_VPWR_c_396_n 0.00157837f $X=1.36 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_33_297#_M1020_g N_VPWR_c_396_n 0.00157837f $X=1.78 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_33_297#_M1022_g N_VPWR_c_397_n 0.00338128f $X=2.2 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_33_297#_c_143_n N_VPWR_c_397_n 5.78397e-19 $X=2.72 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_33_297#_M1002_g N_VPWR_c_403_n 0.00585385f $X=0.94 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_33_297#_M1005_g N_VPWR_c_403_n 0.00585385f $X=1.36 $Y=1.985 $X2=0
+ $Y2=0
cc_141 N_A_33_297#_M1020_g N_VPWR_c_404_n 0.00585385f $X=1.78 $Y=1.985 $X2=0
+ $Y2=0
cc_142 N_A_33_297#_M1022_g N_VPWR_c_404_n 0.00585385f $X=2.2 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_33_297#_M1018_s N_VPWR_c_394_n 0.00227274f $X=0.165 $Y=1.485 $X2=0
+ $Y2=0
cc_144 N_A_33_297#_M1002_g N_VPWR_c_394_n 0.010464f $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A_33_297#_M1005_g N_VPWR_c_394_n 0.0104367f $X=1.36 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_33_297#_M1020_g N_VPWR_c_394_n 0.0104367f $X=1.78 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_33_297#_M1022_g N_VPWR_c_394_n 0.0117628f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_33_297#_c_149_n N_VPWR_c_394_n 0.0122408f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_149 N_A_33_297#_c_149_n N_VPWR_c_407_n 0.0176315f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_150 N_A_33_297#_M1002_g N_Y_c_494_n 2.36323e-19 $X=0.94 $Y=1.985 $X2=0 $Y2=0
cc_151 N_A_33_297#_c_150_n N_Y_c_494_n 0.008553f $X=0.725 $Y=1.54 $X2=0 $Y2=0
cc_152 N_A_33_297#_c_190_p N_Y_c_494_n 0.0171818f $X=2.05 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_33_297#_c_143_n N_Y_c_494_n 0.00220041f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A_33_297#_M1005_g N_Y_c_495_n 0.013192f $X=1.36 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_33_297#_M1020_g N_Y_c_495_n 0.0132199f $X=1.78 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_33_297#_c_190_p N_Y_c_495_n 0.0416643f $X=2.05 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_33_297#_c_143_n N_Y_c_495_n 0.0024854f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_33_297#_c_135_n N_Y_c_510_n 0.00778f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_33_297#_c_136_n N_Y_c_510_n 0.00887971f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_33_297#_c_137_n N_Y_c_510_n 0.00969874f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_33_297#_c_139_n N_Y_c_510_n 0.00598948f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_162 N_A_33_297#_c_190_p N_Y_c_510_n 0.037157f $X=2.05 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_33_297#_c_143_n N_Y_c_510_n 0.00487322f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_33_297#_c_138_n N_Y_c_516_n 0.00219452f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_33_297#_c_190_p N_Y_c_498_n 0.0204549f $X=2.05 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_33_297#_c_143_n N_Y_c_498_n 0.00257112f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_33_297#_M1022_g Y 0.0201894f $X=2.2 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A_33_297#_c_190_p Y 0.0280085f $X=2.05 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_33_297#_c_143_n Y 0.0306882f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_33_297#_c_137_n N_Y_c_493_n 0.00414139f $X=2.3 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_33_297#_c_138_n N_Y_c_493_n 0.00342139f $X=2.72 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_33_297#_c_143_n N_Y_c_493_n 0.00839288f $X=2.72 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_33_297#_c_139_n N_VGND_c_643_n 0.0230021f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_174 N_A_33_297#_c_135_n N_VGND_c_648_n 0.00368123f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_33_297#_c_136_n N_VGND_c_648_n 0.00368123f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_33_297#_c_137_n N_VGND_c_648_n 0.00368123f $X=2.3 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_33_297#_c_138_n N_VGND_c_648_n 0.00368123f $X=2.72 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_33_297#_c_139_n N_VGND_c_648_n 0.0171481f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_179 N_A_33_297#_M1019_d N_VGND_c_657_n 0.00211145f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_180 N_A_33_297#_c_135_n N_VGND_c_657_n 0.00657241f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_33_297#_c_136_n N_VGND_c_657_n 0.00524634f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_33_297#_c_137_n N_VGND_c_657_n 0.00524634f $X=2.3 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_33_297#_c_138_n N_VGND_c_657_n 0.00527354f $X=2.72 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_33_297#_c_139_n N_VGND_c_657_n 0.012188f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_185 N_A_33_297#_c_135_n N_A_225_47#_c_740_n 0.00841925f $X=1.46 $Y=0.995
+ $X2=0 $Y2=0
cc_186 N_A_33_297#_c_136_n N_A_225_47#_c_740_n 0.00795669f $X=1.88 $Y=0.995
+ $X2=0 $Y2=0
cc_187 N_A_33_297#_c_137_n N_A_225_47#_c_740_n 0.00795669f $X=2.3 $Y=0.995 $X2=0
+ $Y2=0
cc_188 N_A_33_297#_c_138_n N_A_225_47#_c_740_n 0.00957159f $X=2.72 $Y=0.995
+ $X2=0 $Y2=0
cc_189 N_A_33_297#_c_139_n N_A_225_47#_c_740_n 0.0139972f $X=0.73 $Y=0.39 $X2=0
+ $Y2=0
cc_190 N_A_33_297#_c_190_p N_A_225_47#_c_740_n 0.00817474f $X=2.05 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_33_297#_c_143_n N_A_225_47#_c_740_n 0.00605207f $X=2.72 $Y=1.16 $X2=0
+ $Y2=0
cc_192 N_A2_c_233_n N_A1_c_315_n 0.0150983f $X=4.4 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_193 N_A2_M1021_g N_A1_M1000_g 0.0150983f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A2_c_234_n A1 0.0176526f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A2_c_235_n A1 0.00106988f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A2_c_234_n N_A1_c_320_n 2.06428e-19 $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A2_c_235_n N_A1_c_320_n 0.0150983f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A2_M1010_g N_VPWR_c_397_n 0.00214918f $X=3.14 $Y=1.985 $X2=0 $Y2=0
cc_199 N_A2_M1010_g N_VPWR_c_401_n 0.00357877f $X=3.14 $Y=1.985 $X2=0 $Y2=0
cc_200 N_A2_M1015_g N_VPWR_c_401_n 0.00357877f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A2_M1016_g N_VPWR_c_401_n 0.00357877f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A2_M1021_g N_VPWR_c_401_n 0.00357877f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A2_M1010_g N_VPWR_c_394_n 0.00655123f $X=3.14 $Y=1.985 $X2=0 $Y2=0
cc_204 N_A2_M1015_g N_VPWR_c_394_n 0.00522516f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A2_M1016_g N_VPWR_c_394_n 0.00522516f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_206 N_A2_M1021_g N_VPWR_c_394_n 0.00525237f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_207 N_A2_M1010_g N_Y_c_496_n 0.0124791f $X=3.14 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A2_c_234_n N_Y_c_496_n 0.01103f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A2_M1015_g N_Y_c_497_n 0.0113168f $X=3.56 $Y=1.985 $X2=0 $Y2=0
cc_210 N_A2_M1016_g N_Y_c_497_n 0.0112944f $X=3.98 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A2_c_234_n N_Y_c_497_n 0.0416944f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_235_n N_Y_c_497_n 0.00214321f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A2_c_234_n N_Y_c_499_n 0.0203891f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A2_c_235_n N_Y_c_499_n 0.00222344f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A2_M1021_g N_Y_c_500_n 5.90444e-19 $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A2_c_234_n N_Y_c_500_n 0.0203891f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A2_c_235_n N_Y_c_500_n 0.00222344f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A2_M1010_g Y 8.86727e-19 $X=3.14 $Y=1.985 $X2=0 $Y2=0
cc_219 N_A2_c_234_n Y 0.0170124f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A2_c_235_n Y 0.00671488f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_c_230_n N_Y_c_493_n 9.46264e-19 $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_M1010_g N_A_561_297#_c_584_n 0.00988743f $X=3.14 $Y=1.985 $X2=0
+ $Y2=0
cc_223 N_A2_M1015_g N_A_561_297#_c_584_n 0.00984328f $X=3.56 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A2_M1016_g N_A_561_297#_c_586_n 0.00984328f $X=3.98 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A2_M1021_g N_A_561_297#_c_586_n 0.0121747f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_226 N_A2_M1021_g N_A_561_297#_c_579_n 2.57315e-19 $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A2_c_230_n N_VGND_c_644_n 0.00268723f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_231_n N_VGND_c_644_n 0.00146448f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_232_n N_VGND_c_645_n 0.00146448f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A2_c_233_n N_VGND_c_645_n 0.00146448f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A2_c_230_n N_VGND_c_648_n 0.00423866f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_231_n N_VGND_c_650_n 0.00423334f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_232_n N_VGND_c_650_n 0.00423334f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_233_n N_VGND_c_652_n 0.00423334f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_230_n N_VGND_c_657_n 0.0057566f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A2_c_231_n N_VGND_c_657_n 0.0057163f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_232_n N_VGND_c_657_n 0.0057163f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_233_n N_VGND_c_657_n 0.0057435f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A2_c_230_n N_A_225_47#_c_757_n 0.00209395f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_230_n N_A_225_47#_c_741_n 0.00485693f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_231_n N_A_225_47#_c_741_n 4.58193e-19 $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A2_c_234_n N_A_225_47#_c_741_n 0.00228728f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A2_c_230_n N_A_225_47#_c_742_n 0.00870364f $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A2_c_231_n N_A_225_47#_c_742_n 0.00865686f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A2_c_234_n N_A_225_47#_c_742_n 0.036111f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A2_c_235_n N_A_225_47#_c_742_n 0.00222133f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A2_c_230_n N_A_225_47#_c_765_n 5.22228e-19 $X=3.14 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A2_c_231_n N_A_225_47#_c_765_n 0.00630972f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_232_n N_A_225_47#_c_765_n 0.00630972f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A2_c_233_n N_A_225_47#_c_765_n 5.22228e-19 $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A2_c_232_n N_A_225_47#_c_743_n 0.00870364f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_c_233_n N_A_225_47#_c_743_n 0.00870364f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_234_n N_A_225_47#_c_743_n 0.036111f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A2_c_235_n N_A_225_47#_c_743_n 0.00222133f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A2_c_232_n N_A_225_47#_c_773_n 5.22228e-19 $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A2_c_233_n N_A_225_47#_c_773_n 0.00630972f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A2_c_231_n N_A_225_47#_c_747_n 0.00113286f $X=3.56 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A2_c_232_n N_A_225_47#_c_747_n 0.00113286f $X=3.98 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A2_c_234_n N_A_225_47#_c_747_n 0.0265405f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_260 N_A2_c_235_n N_A_225_47#_c_747_n 0.00230339f $X=4.4 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A2_c_233_n N_A_225_47#_c_748_n 0.00112787f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A2_c_234_n N_A_225_47#_c_748_n 0.00230276f $X=4.25 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A1_M1000_g N_VPWR_c_398_n 0.00302074f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A1_M1011_g N_VPWR_c_398_n 0.00157837f $X=5.24 $Y=1.985 $X2=0 $Y2=0
cc_265 N_A1_M1011_g N_VPWR_c_399_n 0.00585385f $X=5.24 $Y=1.985 $X2=0 $Y2=0
cc_266 N_A1_M1017_g N_VPWR_c_399_n 0.00585385f $X=5.66 $Y=1.985 $X2=0 $Y2=0
cc_267 N_A1_M1017_g N_VPWR_c_400_n 0.00157837f $X=5.66 $Y=1.985 $X2=0 $Y2=0
cc_268 N_A1_M1023_g N_VPWR_c_400_n 0.00302074f $X=6.08 $Y=1.985 $X2=0 $Y2=0
cc_269 N_A1_M1000_g N_VPWR_c_401_n 0.00585385f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A1_M1023_g N_VPWR_c_405_n 0.00585385f $X=6.08 $Y=1.985 $X2=0 $Y2=0
cc_271 A1 N_VPWR_c_405_n 0.015039f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_272 N_A1_M1000_g N_VPWR_c_394_n 0.010464f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A1_M1011_g N_VPWR_c_394_n 0.0104367f $X=5.24 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A1_M1017_g N_VPWR_c_394_n 0.0104367f $X=5.66 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A1_M1023_g N_VPWR_c_394_n 0.0117628f $X=6.08 $Y=1.985 $X2=0 $Y2=0
cc_276 A1 N_VPWR_c_394_n 0.00854752f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_277 A1 N_A_561_297#_c_579_n 0.00771248f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A1_M1000_g N_A_561_297#_c_580_n 0.0132131f $X=4.82 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A1_M1011_g N_A_561_297#_c_580_n 0.0132273f $X=5.24 $Y=1.985 $X2=0 $Y2=0
cc_280 A1 N_A_561_297#_c_580_n 0.041703f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_281 N_A1_c_320_n N_A_561_297#_c_580_n 0.00211509f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A1_M1017_g N_A_561_297#_c_581_n 0.0132273f $X=5.66 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A1_M1023_g N_A_561_297#_c_581_n 0.0134927f $X=6.08 $Y=1.985 $X2=0 $Y2=0
cc_284 A1 N_A_561_297#_c_581_n 0.041703f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_285 N_A1_c_320_n N_A_561_297#_c_581_n 0.00211509f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_286 A1 N_A_561_297#_c_582_n 0.0358133f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_287 A1 N_A_561_297#_c_599_n 0.0645049f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_288 A1 N_A_561_297#_c_583_n 0.0204549f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_289 N_A1_c_320_n N_A_561_297#_c_583_n 0.00220041f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A1_c_315_n N_VGND_c_646_n 0.00146448f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A1_c_316_n N_VGND_c_646_n 0.00146448f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A1_c_317_n N_VGND_c_647_n 0.00146448f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A1_c_318_n N_VGND_c_647_n 0.00268723f $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A1_c_315_n N_VGND_c_652_n 0.00423334f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A1_c_316_n N_VGND_c_654_n 0.00423334f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A1_c_317_n N_VGND_c_654_n 0.00423334f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A1_c_318_n N_VGND_c_656_n 0.00423334f $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A1_c_315_n N_VGND_c_657_n 0.0057435f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A1_c_316_n N_VGND_c_657_n 0.0057163f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A1_c_317_n N_VGND_c_657_n 0.0057163f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_301 N_A1_c_318_n N_VGND_c_657_n 0.00704237f $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A1_c_315_n N_A_225_47#_c_773_n 0.00630972f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A1_c_316_n N_A_225_47#_c_773_n 5.22228e-19 $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A1_c_315_n N_A_225_47#_c_744_n 0.00870364f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A1_c_316_n N_A_225_47#_c_744_n 0.00870364f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_306 A1 N_A_225_47#_c_744_n 0.0362443f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_307 N_A1_c_320_n N_A_225_47#_c_744_n 0.00222133f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A1_c_315_n N_A_225_47#_c_787_n 5.22228e-19 $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A1_c_316_n N_A_225_47#_c_787_n 0.00630972f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A1_c_317_n N_A_225_47#_c_787_n 0.00630972f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A1_c_318_n N_A_225_47#_c_787_n 5.22228e-19 $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A1_c_317_n N_A_225_47#_c_745_n 0.00870364f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A1_c_318_n N_A_225_47#_c_745_n 0.00999903f $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_314 A1 N_A_225_47#_c_745_n 0.0641689f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_315 N_A1_c_320_n N_A_225_47#_c_745_n 0.00222133f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A1_c_317_n N_A_225_47#_c_746_n 5.22228e-19 $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A1_c_318_n N_A_225_47#_c_746_n 0.00630972f $X=6.08 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A1_c_315_n N_A_225_47#_c_748_n 0.00112787f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_319 A1 N_A_225_47#_c_748_n 0.0108485f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_320 N_A1_c_316_n N_A_225_47#_c_749_n 0.00113286f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A1_c_317_n N_A_225_47#_c_749_n 0.00113286f $X=5.66 $Y=0.995 $X2=0 $Y2=0
cc_322 A1 N_A_225_47#_c_749_n 0.0266272f $X=6.585 $Y=1.105 $X2=0 $Y2=0
cc_323 N_A1_c_320_n N_A_225_47#_c_749_n 0.00230339f $X=6.08 $Y=1.16 $X2=0 $Y2=0
cc_324 N_VPWR_c_394_n N_Y_M1002_s 0.00423495f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_325 N_VPWR_c_394_n N_Y_M1020_s 0.00284632f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_326 N_VPWR_c_394_n N_Y_M1010_d 0.00216833f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_394_n N_Y_M1016_d 0.00216833f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_c_403_n N_Y_c_544_n 0.012815f $X=1.445 $Y=2.72 $X2=0 $Y2=0
cc_329 N_VPWR_c_394_n N_Y_c_544_n 0.00801045f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_330 N_VPWR_M1005_d N_Y_c_495_n 0.00165831f $X=1.435 $Y=1.485 $X2=0 $Y2=0
cc_331 N_VPWR_c_396_n N_Y_c_495_n 0.0126919f $X=1.57 $Y=1.96 $X2=0 $Y2=0
cc_332 N_VPWR_c_404_n N_Y_c_548_n 0.0142343f $X=2.285 $Y=2.72 $X2=0 $Y2=0
cc_333 N_VPWR_c_394_n N_Y_c_548_n 0.00955092f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_334 N_VPWR_M1022_d Y 0.00342775f $X=2.275 $Y=1.485 $X2=0 $Y2=0
cc_335 N_VPWR_c_397_n Y 0.0171277f $X=2.41 $Y=1.96 $X2=0 $Y2=0
cc_336 N_VPWR_c_394_n N_A_561_297#_M1010_s 0.0020932f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_337 N_VPWR_c_394_n N_A_561_297#_M1015_s 0.00215203f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_394_n N_A_561_297#_M1021_s 0.00246446f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_394_n N_A_561_297#_M1011_d 0.00284632f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_394_n N_A_561_297#_M1023_d 0.00333334f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_397_n N_A_561_297#_c_577_n 0.0308495f $X=2.41 $Y=1.96 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_401_n N_A_561_297#_c_584_n 0.0330174f $X=4.905 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_394_n N_A_561_297#_c_584_n 0.0204627f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_397_n N_A_561_297#_c_578_n 0.0113145f $X=2.41 $Y=1.96 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_401_n N_A_561_297#_c_578_n 0.0180409f $X=4.905 $Y=2.72 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_394_n N_A_561_297#_c_578_n 0.0107739f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_401_n N_A_561_297#_c_586_n 0.0330174f $X=4.905 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_394_n N_A_561_297#_c_586_n 0.0204627f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_401_n N_A_561_297#_c_615_n 0.0143053f $X=4.905 $Y=2.72 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_394_n N_A_561_297#_c_615_n 0.00962794f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_M1000_s N_A_561_297#_c_580_n 0.00165831f $X=4.895 $Y=1.485 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_398_n N_A_561_297#_c_580_n 0.0126919f $X=5.03 $Y=1.96 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_399_n N_A_561_297#_c_619_n 0.0142343f $X=5.745 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_394_n N_A_561_297#_c_619_n 0.00955092f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_355 N_VPWR_M1017_s N_A_561_297#_c_581_n 0.00165831f $X=5.735 $Y=1.485 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_400_n N_A_561_297#_c_581_n 0.0126919f $X=5.87 $Y=1.96 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_405_n N_A_561_297#_c_599_n 0.0158369f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_394_n N_A_561_297#_c_599_n 0.00955092f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_401_n N_A_561_297#_c_625_n 0.0142933f $X=4.905 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_394_n N_A_561_297#_c_625_n 0.00962421f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_361 N_Y_c_496_n N_A_561_297#_M1010_s 0.00158868f $X=3.225 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_362 Y N_A_561_297#_M1010_s 0.0018459f $X=2.445 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_363 N_Y_c_497_n N_A_561_297#_M1015_s 0.00166124f $X=4.065 $Y=1.535 $X2=0
+ $Y2=0
cc_364 N_Y_c_496_n N_A_561_297#_c_577_n 0.00921788f $X=3.225 $Y=1.535 $X2=0
+ $Y2=0
cc_365 Y N_A_561_297#_c_577_n 0.0105628f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_366 N_Y_M1010_d N_A_561_297#_c_584_n 0.00312348f $X=3.215 $Y=1.485 $X2=0
+ $Y2=0
cc_367 N_Y_c_496_n N_A_561_297#_c_584_n 0.00322336f $X=3.225 $Y=1.535 $X2=0
+ $Y2=0
cc_368 N_Y_c_497_n N_A_561_297#_c_584_n 0.00322336f $X=4.065 $Y=1.535 $X2=0
+ $Y2=0
cc_369 N_Y_c_499_n N_A_561_297#_c_584_n 0.0118865f $X=3.35 $Y=1.62 $X2=0 $Y2=0
cc_370 N_Y_c_497_n N_A_561_297#_c_636_n 0.0127256f $X=4.065 $Y=1.535 $X2=0 $Y2=0
cc_371 N_Y_M1016_d N_A_561_297#_c_586_n 0.00312348f $X=4.055 $Y=1.485 $X2=0
+ $Y2=0
cc_372 N_Y_c_497_n N_A_561_297#_c_586_n 0.00322336f $X=4.065 $Y=1.535 $X2=0
+ $Y2=0
cc_373 N_Y_c_500_n N_A_561_297#_c_586_n 0.0118865f $X=4.19 $Y=1.62 $X2=0 $Y2=0
cc_374 N_Y_c_500_n N_A_561_297#_c_579_n 0.00271526f $X=4.19 $Y=1.62 $X2=0 $Y2=0
cc_375 N_Y_M1003_d N_VGND_c_657_n 0.00220248f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_376 N_Y_M1024_d N_VGND_c_657_n 0.00220248f $X=2.375 $Y=0.235 $X2=0 $Y2=0
cc_377 N_Y_c_510_n N_A_225_47#_M1009_s 0.00334902f $X=2.445 $Y=0.73 $X2=0 $Y2=0
cc_378 N_Y_M1003_d N_A_225_47#_c_740_n 0.00318958f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_379 N_Y_M1024_d N_A_225_47#_c_740_n 0.00317561f $X=2.375 $Y=0.235 $X2=0 $Y2=0
cc_380 N_Y_c_510_n N_A_225_47#_c_740_n 0.0489906f $X=2.445 $Y=0.73 $X2=0 $Y2=0
cc_381 N_Y_c_516_n N_A_225_47#_c_740_n 0.0131314f $X=2.56 $Y=0.815 $X2=0 $Y2=0
cc_382 Y N_A_225_47#_c_740_n 0.00407994f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_383 N_Y_c_496_n N_A_225_47#_c_741_n 0.00638629f $X=3.225 $Y=1.535 $X2=0 $Y2=0
cc_384 Y N_A_225_47#_c_741_n 0.00447631f $X=2.445 $Y=1.445 $X2=0 $Y2=0
cc_385 N_Y_c_493_n N_A_225_47#_c_741_n 0.00406049f $X=2.67 $Y=1.075 $X2=0 $Y2=0
cc_386 N_A_561_297#_c_579_n N_A_225_47#_c_748_n 0.00658191f $X=4.61 $Y=1.625
+ $X2=0 $Y2=0
cc_387 N_VGND_c_657_n N_A_225_47#_M1003_s 0.0021262f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_388 N_VGND_c_657_n N_A_225_47#_M1009_s 0.00218617f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_657_n N_A_225_47#_M1025_s 0.00218529f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_657_n N_A_225_47#_M1004_s 0.00215201f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_657_n N_A_225_47#_M1008_s 0.00215201f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_657_n N_A_225_47#_M1012_d 0.00215201f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_657_n N_A_225_47#_M1014_d 0.00209319f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_648_n N_A_225_47#_c_740_n 0.0745699f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_657_n N_A_225_47#_c_740_n 0.06065f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_648_n N_A_225_47#_c_757_n 0.0114777f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_657_n N_A_225_47#_c_757_n 0.00913984f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_M1001_d N_A_225_47#_c_742_n 0.00162089f $X=3.215 $Y=0.235 $X2=0
+ $Y2=0
cc_399 N_VGND_c_644_n N_A_225_47#_c_742_n 0.0122559f $X=3.35 $Y=0.39 $X2=0 $Y2=0
cc_400 N_VGND_c_648_n N_A_225_47#_c_742_n 0.00198695f $X=3.265 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_650_n N_A_225_47#_c_742_n 0.00198695f $X=4.105 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_657_n N_A_225_47#_c_742_n 0.00835832f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_650_n N_A_225_47#_c_765_n 0.0188551f $X=4.105 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_c_657_n N_A_225_47#_c_765_n 0.0122069f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_M1007_d N_A_225_47#_c_743_n 0.00162089f $X=4.055 $Y=0.235 $X2=0
+ $Y2=0
cc_406 N_VGND_c_645_n N_A_225_47#_c_743_n 0.0122559f $X=4.19 $Y=0.39 $X2=0 $Y2=0
cc_407 N_VGND_c_650_n N_A_225_47#_c_743_n 0.00198695f $X=4.105 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_c_652_n N_A_225_47#_c_743_n 0.00198695f $X=4.945 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_657_n N_A_225_47#_c_743_n 0.00835832f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_652_n N_A_225_47#_c_773_n 0.0188551f $X=4.945 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_657_n N_A_225_47#_c_773_n 0.0122069f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_M1006_s N_A_225_47#_c_744_n 0.00162089f $X=4.895 $Y=0.235 $X2=0
+ $Y2=0
cc_413 N_VGND_c_646_n N_A_225_47#_c_744_n 0.0122559f $X=5.03 $Y=0.39 $X2=0 $Y2=0
cc_414 N_VGND_c_652_n N_A_225_47#_c_744_n 0.00198695f $X=4.945 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_654_n N_A_225_47#_c_744_n 0.00198695f $X=5.785 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_657_n N_A_225_47#_c_744_n 0.00835832f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_c_654_n N_A_225_47#_c_787_n 0.0188551f $X=5.785 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_657_n N_A_225_47#_c_787_n 0.0122069f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_M1013_s N_A_225_47#_c_745_n 0.00162089f $X=5.735 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_VGND_c_647_n N_A_225_47#_c_745_n 0.0122559f $X=5.87 $Y=0.39 $X2=0 $Y2=0
cc_421 N_VGND_c_654_n N_A_225_47#_c_745_n 0.00198695f $X=5.785 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_656_n N_A_225_47#_c_745_n 0.00198695f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_657_n N_A_225_47#_c_745_n 0.00835832f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_656_n N_A_225_47#_c_746_n 0.0209752f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_657_n N_A_225_47#_c_746_n 0.0124119f $X=6.67 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a2bb2o_4.pex.spice
* Created: Tue Sep  1 18:54:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%B1 3 6 8 10 13 15 18 22 23 25 28 29 30
c83 30 0 8.57496e-20 $X=0.41 $Y=0.995
c84 29 0 1.22288e-19 $X=0.41 $Y=1.16
c85 23 0 3.46433e-19 $X=1.73 $Y=1.16
c86 15 0 7.58469e-20 $X=1.515 $Y=1.53
r87 28 31 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r88 28 30 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r89 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r90 25 37 8.29932 $w=4.88e-07 $l=3.4e-07 $layer=LI1_cond $X=0.33 $Y=1.19
+ $X2=0.33 $Y2=1.53
r91 25 29 0.732293 $w=4.88e-07 $l=3e-08 $layer=LI1_cond $X=0.33 $Y=1.19 $X2=0.33
+ $Y2=1.16
r92 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r93 19 22 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.6 $Y=1.16 $X2=1.73
+ $Y2=1.16
r94 17 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=1.245 $X2=1.6
+ $Y2=1.16
r95 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.6 $Y=1.245 $X2=1.6
+ $Y2=1.445
r96 16 37 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.575 $Y=1.53
+ $X2=0.33 $Y2=1.53
r97 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.53
+ $X2=1.6 $Y2=1.445
r98 15 16 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.515 $Y=1.53
+ $X2=0.575 $Y2=1.53
r99 11 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.985
r101 8 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r102 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r103 6 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r104 3 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%B2 1 3 6 8 10 13 15 22
c45 15 0 1.95758e-19 $X=1.155 $Y=1.19
c46 6 0 1.22288e-19 $X=0.89 $Y=1.985
c47 1 0 1.52215e-19 $X=0.89 $Y=0.995
r48 20 22 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.31
+ $Y2=1.16
r49 17 20 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=1.1
+ $Y2=1.16
r50 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r51 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.985
r53 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r54 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r55 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r56 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325 $X2=0.89
+ $Y2=1.985
r57 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995 $X2=0.89
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A_415_21# 1 2 3 10 12 15 17 19 22 24 27 30
+ 32 33 34 35 39 41 45 47 49 50
c139 41 0 7.82236e-20 $X=4.395 $Y=0.815
c140 27 0 1.85277e-19 $X=2.78 $Y=1.16
c141 15 0 7.58469e-20 $X=2.15 $Y=1.985
r142 55 57 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=2.57 $Y2=1.16
r143 50 53 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=1.875
+ $X2=4.14 $Y2=1.96
r144 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=0.725
+ $X2=4.56 $Y2=0.39
r145 42 49 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0.815
+ $X2=3.72 $Y2=0.815
r146 41 43 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=4.56 $Y2=0.725
r147 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.395 $Y=0.815
+ $X2=3.885 $Y2=0.815
r148 37 49 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.72 $Y=0.725
+ $X2=3.72 $Y2=0.815
r149 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.72 $Y=0.725
+ $X2=3.72 $Y2=0.39
r150 36 48 2.30104 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=3.305 $Y=1.875
+ $X2=3.135 $Y2=1.875
r151 35 50 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.015 $Y=1.875
+ $X2=4.14 $Y2=1.875
r152 35 36 43.7475 $w=1.78e-07 $l=7.1e-07 $layer=LI1_cond $X=4.015 $Y=1.875
+ $X2=3.305 $Y2=1.875
r153 33 49 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0.815
+ $X2=3.72 $Y2=0.815
r154 33 34 25.2626 $w=1.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.555 $Y=0.815
+ $X2=3.145 $Y2=0.815
r155 32 48 20.2107 $w=2.35e-07 $l=4.20357e-07 $layer=LI1_cond $X=3.05 $Y=1.495
+ $X2=3.135 $Y2=1.875
r156 31 47 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.245
+ $X2=3.05 $Y2=1.16
r157 31 32 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.05 $Y=1.245
+ $X2=3.05 $Y2=1.495
r158 30 47 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.075
+ $X2=3.05 $Y2=1.16
r159 29 34 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.05 $Y=0.905
+ $X2=3.145 $Y2=0.815
r160 29 30 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.05 $Y=0.905
+ $X2=3.05 $Y2=1.075
r161 27 57 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=1.16
+ $X2=2.57 $Y2=1.16
r162 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.16 $X2=2.78 $Y2=1.16
r163 24 47 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.955 $Y=1.16
+ $X2=3.05 $Y2=1.16
r164 24 26 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.955 $Y=1.16
+ $X2=2.78 $Y2=1.16
r165 20 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.16
r166 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=1.325
+ $X2=2.57 $Y2=1.985
r167 17 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=1.16
r168 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.57 $Y=0.995
+ $X2=2.57 $Y2=0.56
r169 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r170 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r171 10 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=1.16
r172 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.15 $Y=0.995
+ $X2=2.15 $Y2=0.56
r173 3 53 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.96
r174 2 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.39
r175 1 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A1_N 3 6 8 10 13 15 18 19 23 25 28
c90 28 0 5.15455e-19 $X=4.77 $Y=1.16
c91 18 0 1.85277e-19 $X=3.39 $Y=1.105
c92 13 0 1.47656e-19 $X=4.77 $Y=1.985
c93 8 0 7.82236e-20 $X=4.77 $Y=0.995
r94 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=1.325
r95 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.16
+ $X2=3.48 $Y2=0.995
r96 19 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.16 $X2=4.77 $Y2=1.16
r97 18 34 18.5 $w=2.44e-07 $l=3.7e-07 $layer=LI1_cond $X=3.48 $Y=1.16 $X2=3.48
+ $Y2=1.53
r98 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.16 $X2=3.48 $Y2=1.16
r99 17 19 9.12351 $w=3.58e-07 $l=2.85e-07 $layer=LI1_cond $X=4.785 $Y=1.445
+ $X2=4.785 $Y2=1.16
r100 16 34 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=1.53
+ $X2=3.48 $Y2=1.53
r101 15 17 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=4.605 $Y=1.53
+ $X2=4.785 $Y2=1.445
r102 15 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.605 $Y=1.53
+ $X2=3.645 $Y2=1.53
r103 11 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.16
r104 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.77 $Y=1.325
+ $X2=4.77 $Y2=1.985
r105 8 28 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.16
r106 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r107 6 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.51 $Y=1.985
+ $X2=3.51 $Y2=1.325
r108 3 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.56
+ $X2=3.51 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A2_N 1 3 6 8 10 13 15 21 22
r48 20 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.145 $Y=1.16
+ $X2=4.35 $Y2=1.16
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.16 $X2=4.145 $Y2=1.16
r50 17 20 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=4.145 $Y2=1.16
r51 15 21 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=4.145 $Y2=1.175
r52 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.35 $Y=1.325
+ $X2=4.35 $Y2=1.985
r54 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.35 $Y=0.995
+ $X2=4.35 $Y2=0.56
r56 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=1.325
+ $X2=3.93 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.93 $Y=1.325 $X2=3.93
+ $Y2=1.985
r58 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995 $X2=3.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A_193_47# 1 2 3 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 42 45 46 51 55 59 61 62 68 69 77 83
c178 69 0 8.54342e-20 $X=5.315 $Y=1.53
c179 68 0 1.47656e-19 $X=5.315 $Y=1.53
c180 55 0 8.57496e-20 $X=1.1 $Y=0.73
c181 46 0 1.81154e-19 $X=5.46 $Y=1.16
c182 38 0 1.15369e-20 $X=2.195 $Y=0.82
c183 10 0 7.82236e-20 $X=5.19 $Y=0.995
r184 83 85 11.7175 $w=3.54e-07 $l=3.4e-07 $layer=LI1_cond $X=2.427 $Y=1.62
+ $X2=2.427 $Y2=1.96
r185 74 75 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.61 $Y=1.16
+ $X2=6.03 $Y2=1.16
r186 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.315 $Y=1.53
+ $X2=5.315 $Y2=1.53
r187 65 83 3.10169 $w=3.54e-07 $l=9e-08 $layer=LI1_cond $X=2.427 $Y=1.53
+ $X2=2.427 $Y2=1.62
r188 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.53
+ $X2=2.535 $Y2=1.53
r189 62 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.53
+ $X2=2.535 $Y2=1.53
r190 61 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.17 $Y=1.53
+ $X2=5.315 $Y2=1.53
r191 61 62 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=5.17 $Y=1.53
+ $X2=2.68 $Y2=1.53
r192 60 69 10.106 $w=3.23e-07 $l=2.85e-07 $layer=LI1_cond $X=5.297 $Y=1.245
+ $X2=5.297 $Y2=1.53
r193 55 57 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=1.102 $Y=0.73
+ $X2=1.102 $Y2=0.82
r194 52 77 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.21 $Y=1.16
+ $X2=6.45 $Y2=1.16
r195 52 75 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.16
+ $X2=6.03 $Y2=1.16
r196 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=1.16 $X2=6.21 $Y2=1.16
r197 49 74 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.53 $Y=1.16 $X2=5.61
+ $Y2=1.16
r198 49 71 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.53 $Y=1.16
+ $X2=5.19 $Y2=1.16
r199 48 51 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.53 $Y=1.16
+ $X2=6.21 $Y2=1.16
r200 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.16 $X2=5.53 $Y2=1.16
r201 46 60 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=5.46 $Y=1.16
+ $X2=5.297 $Y2=1.245
r202 46 48 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.46 $Y=1.16 $X2=5.53
+ $Y2=1.16
r203 45 65 5.96567 $w=3.54e-07 $l=1.52414e-07 $layer=LI1_cond $X=2.34 $Y=1.415
+ $X2=2.427 $Y2=1.53
r204 44 59 3.46198 $w=2.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.34 $Y=0.905
+ $X2=2.36 $Y2=0.82
r205 44 45 26.9351 $w=2.08e-07 $l=5.1e-07 $layer=LI1_cond $X=2.34 $Y=0.905
+ $X2=2.34 $Y2=1.415
r206 40 59 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.36 $Y2=0.82
r207 40 42 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.36 $Y=0.735
+ $X2=2.36 $Y2=0.39
r208 39 57 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.27 $Y=0.82
+ $X2=1.102 $Y2=0.82
r209 38 59 3.05049 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=2.36 $Y2=0.82
r210 38 39 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=1.27 $Y2=0.82
r211 34 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.16
r212 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.45 $Y=1.325
+ $X2=6.45 $Y2=1.985
r213 31 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=1.16
r214 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.45 $Y=0.995
+ $X2=6.45 $Y2=0.56
r215 27 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.16
r216 27 29 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.03 $Y=1.325
+ $X2=6.03 $Y2=1.985
r217 24 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=1.16
r218 24 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.03 $Y=0.995
+ $X2=6.03 $Y2=0.56
r219 20 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.16
r220 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.61 $Y=1.325
+ $X2=5.61 $Y2=1.985
r221 17 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=1.16
r222 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.61 $Y=0.995
+ $X2=5.61 $Y2=0.56
r223 13 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.16
r224 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.19 $Y=1.325
+ $X2=5.19 $Y2=1.985
r225 10 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=1.16
r226 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.19 $Y=0.995
+ $X2=5.19 $Y2=0.56
r227 3 85 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.96
r228 3 83 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.36 $Y2=1.62
r229 2 42 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.225
+ $Y=0.235 $X2=2.36 $Y2=0.39
r230 1 55 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A_27_297# 1 2 3 4 15 17 18 21 23 31 33 34
+ 35 38
c52 23 0 1.50675e-19 $X=1.815 $Y=1.87
r53 38 40 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.78 $Y=2.3 $X2=2.78
+ $Y2=2.38
r54 33 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.78 $Y2=2.38
r55 33 34 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.655 $Y=2.38
+ $X2=2.065 $Y2=2.38
r56 29 36 3.98977 $w=2.3e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.96 $Y=1.785
+ $X2=1.94 $Y2=1.87
r57 29 31 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=1.785
+ $X2=1.96 $Y2=1.62
r58 26 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=2.065 $Y2=2.38
r59 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.94 $Y=2.295
+ $X2=1.94 $Y2=1.96
r60 25 36 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.955
+ $X2=1.94 $Y2=1.87
r61 25 28 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.94 $Y=1.955
+ $X2=1.94 $Y2=1.96
r62 24 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=1.87
+ $X2=1.1 $Y2=1.87
r63 23 36 2.45049 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=1.87
+ $X2=1.94 $Y2=1.87
r64 23 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.815 $Y=1.87
+ $X2=1.225 $Y2=1.87
r65 19 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.955
+ $X2=1.1 $Y2=1.87
r66 19 21 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.1 $Y=1.955 $X2=1.1
+ $Y2=1.96
r67 17 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=1.87
+ $X2=1.1 $Y2=1.87
r68 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.975 $Y=1.87
+ $X2=0.385 $Y2=1.87
r69 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.385 $Y2=1.87
r70 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.955
+ $X2=0.26 $Y2=1.96
r71 4 38 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.485 $X2=2.78 $Y2=2.3
r72 3 31 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.62
r73 3 28 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=1.96
r74 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.96
r75 1 15 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 43 46 47
+ 48 49 50 52 57 72 79 80 83 86 89 92
c118 33 0 1.23485e-19 $X=4.98 $Y=1.96
r119 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r121 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 80 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=6.67 $Y2=2.72
r124 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 77 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=6.66 $Y2=2.72
r126 77 79 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.785 $Y=2.72
+ $X2=7.13 $Y2=2.72
r127 76 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r128 76 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r129 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r130 73 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=5.82 $Y2=2.72
r131 73 75 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.945 $Y=2.72
+ $X2=6.21 $Y2=2.72
r132 72 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.66 $Y2=2.72
r133 72 75 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.21 $Y2=2.72
r134 71 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r135 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r136 68 71 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 67 70 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r138 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 65 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 65 87 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=1.61 $Y2=2.72
r141 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r142 62 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.52 $Y2=2.72
r143 62 64 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=2.99 $Y2=2.72
r144 61 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r145 61 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r147 58 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=0.68 $Y2=2.72
r148 58 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.805 $Y=2.72
+ $X2=1.15 $Y2=2.72
r149 57 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.52 $Y2=2.72
r150 57 60 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.15 $Y2=2.72
r151 52 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=2.72
+ $X2=0.68 $Y2=2.72
r152 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.555 $Y=2.72
+ $X2=0.23 $Y2=2.72
r153 50 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 50 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 48 70 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.83 $Y2=2.72
r156 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=2.72
+ $X2=4.98 $Y2=2.72
r157 46 64 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.175 $Y=2.72
+ $X2=2.99 $Y2=2.72
r158 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.175 $Y=2.72
+ $X2=3.3 $Y2=2.72
r159 45 67 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.45 $Y2=2.72
r160 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.3 $Y2=2.72
r161 41 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=2.72
r162 41 43 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=6.66 $Y=2.635
+ $X2=6.66 $Y2=1.99
r163 37 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.72
r164 37 39 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.82 $Y2=2.33
r165 36 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.98 $Y2=2.72
r166 35 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.82 $Y2=2.72
r167 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.695 $Y=2.72
+ $X2=5.105 $Y2=2.72
r168 31 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=2.72
r169 31 33 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.98 $Y=2.635
+ $X2=4.98 $Y2=1.96
r170 27 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2.72
r171 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.3 $Y=2.635
+ $X2=3.3 $Y2=2.34
r172 23 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.72
r173 23 25 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.52 $Y=2.635
+ $X2=1.52 $Y2=2.3
r174 19 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r175 19 21 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.3
r176 6 43 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=6.525
+ $Y=1.485 $X2=6.66 $Y2=1.99
r177 5 39 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=2.33
r178 4 33 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=1.96
r179 3 29 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.485 $X2=3.3 $Y2=2.34
r180 2 25 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.3
r181 1 21 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A_717_297# 1 2 7 11 14
c17 11 0 1.25382e-19 $X=4.56 $Y=1.96
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.72 $Y=2.3 $X2=3.72
+ $Y2=2.38
r19 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=2.295
+ $X2=4.56 $Y2=1.96
r20 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=2.38
+ $X2=3.72 $Y2=2.38
r21 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.435 $Y=2.38
+ $X2=4.56 $Y2=2.295
r22 7 8 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.435 $Y=2.38 $X2=3.845
+ $Y2=2.38
r23 2 11 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.96
r24 1 14 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 36
+ 43 44 48
c81 24 0 7.82236e-20 $X=5.565 $Y=0.815
r82 44 48 3.03757 $w=3.1e-07 $l=1.2e-07 $layer=LI1_cond $X=6.765 $Y=1.535
+ $X2=6.765 $Y2=1.415
r83 43 48 8.36451 $w=3.08e-07 $l=2.25e-07 $layer=LI1_cond $X=6.765 $Y=1.19
+ $X2=6.765 $Y2=1.415
r84 42 43 10.595 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=0.905
+ $X2=6.765 $Y2=1.19
r85 40 41 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.24 $Y=1.62
+ $X2=6.24 $Y2=1.87
r86 37 44 7.89872 $w=4.08e-07 $l=2.45e-07 $layer=LI1_cond $X=6.365 $Y=1.535
+ $X2=6.61 $Y2=1.535
r87 36 40 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=1.535
+ $X2=6.24 $Y2=1.62
r88 36 37 0.964185 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=6.24 $Y=1.535
+ $X2=6.365 $Y2=1.535
r89 34 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.405 $Y=0.815
+ $X2=6.24 $Y2=0.815
r90 33 42 7.45983 $w=1.8e-07 $l=1.94872e-07 $layer=LI1_cond $X=6.61 $Y=0.815
+ $X2=6.765 $Y2=0.905
r91 33 34 12.6313 $w=1.78e-07 $l=2.05e-07 $layer=LI1_cond $X=6.61 $Y=0.815
+ $X2=6.405 $Y2=0.815
r92 29 41 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.24 $Y=1.955
+ $X2=6.24 $Y2=1.87
r93 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.24 $Y=1.955
+ $X2=6.24 $Y2=1.96
r94 25 35 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.24 $Y=0.725 $X2=6.24
+ $Y2=0.815
r95 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.24 $Y=0.725
+ $X2=6.24 $Y2=0.39
r96 23 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=6.24 $Y2=0.815
r97 23 24 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.075 $Y=0.815
+ $X2=5.565 $Y2=0.815
r98 21 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.115 $Y=1.87
+ $X2=6.24 $Y2=1.87
r99 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.115 $Y=1.87
+ $X2=5.525 $Y2=1.87
r100 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.4 $Y=1.955
+ $X2=5.525 $Y2=1.87
r101 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.4 $Y=1.955 $X2=5.4
+ $Y2=1.96
r102 13 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.4 $Y=0.725
+ $X2=5.565 $Y2=0.815
r103 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.4 $Y=0.725
+ $X2=5.4 $Y2=0.39
r104 4 40 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.62
r105 4 31 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.485 $X2=6.24 $Y2=1.96
r106 3 19 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.96
r107 2 27 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.105
+ $Y=0.235 $X2=6.24 $Y2=0.39
r108 1 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 38 42 46
+ 49 50 52 53 54 55 57 58 59 84 85 93 96 98
r120 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r121 95 96 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.235
+ $X2=3.385 $Y2=0.235
r122 91 95 5.7935 $w=6.38e-07 $l=3.1e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=3.3 $Y2=0.235
r123 91 93 12.8464 $w=6.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=2.695 $Y2=0.235
r124 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r125 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r126 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r127 82 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r128 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r129 79 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=0 $X2=5.82
+ $Y2=0
r130 79 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.21 $Y2=0
r131 78 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r132 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r133 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r134 75 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r135 74 96 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=3.385 $Y2=0
r136 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r137 71 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r138 70 93 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=2.695 $Y2=0
r139 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r140 67 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r141 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r142 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r143 63 66 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r144 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r145 61 88 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r146 61 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r147 59 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r148 59 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r149 57 81 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.575 $Y=0
+ $X2=6.21 $Y2=0
r150 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.575 $Y=0 $X2=6.66
+ $Y2=0
r151 56 84 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.13 $Y2=0
r152 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0 $X2=6.66
+ $Y2=0
r153 54 77 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.83
+ $Y2=0
r154 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=0 $X2=4.98
+ $Y2=0
r155 52 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=3.91 $Y2=0
r156 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0 $X2=4.14
+ $Y2=0
r157 51 77 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.83 $Y2=0
r158 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.14
+ $Y2=0
r159 49 66 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.61
+ $Y2=0
r160 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.94
+ $Y2=0
r161 48 70 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.53 $Y2=0
r162 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.94
+ $Y2=0
r163 44 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0
r164 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.66 $Y=0.085
+ $X2=6.66 $Y2=0.39
r165 40 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r166 40 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.39
r167 39 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=4.98
+ $Y2=0
r168 38 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.82
+ $Y2=0
r169 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.065 $Y2=0
r170 34 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0
r171 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.98 $Y=0.085
+ $X2=4.98 $Y2=0.39
r172 30 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0
r173 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.14 $Y=0.085
+ $X2=4.14 $Y2=0.39
r174 26 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0
r175 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.94 $Y=0.085
+ $X2=1.94 $Y2=0.39
r176 22 88 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r177 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r178 7 46 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.525
+ $Y=0.235 $X2=6.66 $Y2=0.39
r179 6 42 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.39
r180 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.39
r181 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.39
r182 3 95 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.645
+ $Y=0.235 $X2=3.3 $Y2=0.39
r183 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.39
r184 1 24 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__A2BB2O_4%A_109_47# 1 2 7 9 13
c21 9 0 1.40678e-19 $X=0.68 $Y=0.73
r22 11 16 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.765 $Y=0.365
+ $X2=0.64 $Y2=0.365
r23 11 13 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=0.765 $Y=0.365
+ $X2=1.52 $Y2=0.365
r24 7 16 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.64 $Y=0.475 $X2=0.64
+ $Y2=0.365
r25 7 9 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.64 $Y=0.475
+ $X2=0.64 $Y2=0.73
r26 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
r27 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.39
r28 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.73
.ends


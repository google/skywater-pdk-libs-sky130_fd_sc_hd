* NGSPICE file created from sky130_fd_sc_hd__lpflow_isobufsrc_1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__lpflow_isobufsrc_1 A SLEEP VGND VNB VPB VPWR X
M1000 a_265_297# SLEEP VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=3.146e+11p ps=2.78e+06u
M1001 X SLEEP VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=3.695e+11p ps=3.79e+06u
M1002 X a_74_47# a_265_297# VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1003 VGND A a_74_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1004 VGND a_74_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A a_74_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends


* File: sky130_fd_sc_hd__nor4b_4.spice.SKY130_FD_SC_HD__NOR4B_4.pxi
* Created: Thu Aug 27 14:33:16 2020
* 
x_PM_SKY130_FD_SC_HD__NOR4B_4%A N_A_c_134_n N_A_M1015_g N_A_M1003_g N_A_c_135_n
+ N_A_M1018_g N_A_M1005_g N_A_c_136_n N_A_M1022_g N_A_M1023_g N_A_c_137_n
+ N_A_M1033_g N_A_M1030_g A N_A_c_138_n N_A_c_139_n
+ PM_SKY130_FD_SC_HD__NOR4B_4%A
x_PM_SKY130_FD_SC_HD__NOR4B_4%B N_B_c_210_n N_B_M1019_g N_B_M1000_g N_B_c_211_n
+ N_B_M1024_g N_B_M1006_g N_B_c_212_n N_B_M1028_g N_B_M1026_g N_B_c_213_n
+ N_B_M1029_g N_B_M1031_g B N_B_c_214_n N_B_c_215_n
+ PM_SKY130_FD_SC_HD__NOR4B_4%B
x_PM_SKY130_FD_SC_HD__NOR4B_4%C N_C_c_289_n N_C_M1012_g N_C_M1001_g N_C_c_290_n
+ N_C_M1016_g N_C_M1010_g N_C_c_291_n N_C_M1020_g N_C_M1014_g N_C_c_292_n
+ N_C_M1025_g N_C_M1032_g C N_C_c_293_n N_C_c_294_n
+ PM_SKY130_FD_SC_HD__NOR4B_4%C
x_PM_SKY130_FD_SC_HD__NOR4B_4%A_1191_21# N_A_1191_21#_M1009_s
+ N_A_1191_21#_M1011_s N_A_1191_21#_c_368_n N_A_1191_21#_M1008_g
+ N_A_1191_21#_M1002_g N_A_1191_21#_c_369_n N_A_1191_21#_M1013_g
+ N_A_1191_21#_M1004_g N_A_1191_21#_c_370_n N_A_1191_21#_M1017_g
+ N_A_1191_21#_M1007_g N_A_1191_21#_c_371_n N_A_1191_21#_M1021_g
+ N_A_1191_21#_M1027_g N_A_1191_21#_c_423_p N_A_1191_21#_c_372_n
+ N_A_1191_21#_c_381_n N_A_1191_21#_c_382_n N_A_1191_21#_c_383_n
+ N_A_1191_21#_c_373_n N_A_1191_21#_c_374_n N_A_1191_21#_c_384_n
+ N_A_1191_21#_c_396_p N_A_1191_21#_c_375_n N_A_1191_21#_c_376_n
+ PM_SKY130_FD_SC_HD__NOR4B_4%A_1191_21#
x_PM_SKY130_FD_SC_HD__NOR4B_4%D_N N_D_N_M1009_g N_D_N_M1011_g D_N N_D_N_c_487_n
+ N_D_N_c_488_n D_N PM_SKY130_FD_SC_HD__NOR4B_4%D_N
x_PM_SKY130_FD_SC_HD__NOR4B_4%A_27_297# N_A_27_297#_M1003_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1030_s N_A_27_297#_M1006_s N_A_27_297#_M1031_s
+ N_A_27_297#_c_515_n N_A_27_297#_c_516_n N_A_27_297#_c_517_n
+ N_A_27_297#_c_546_p N_A_27_297#_c_518_n N_A_27_297#_c_519_n
+ N_A_27_297#_c_547_p N_A_27_297#_c_537_n N_A_27_297#_c_566_p
+ N_A_27_297#_c_520_n N_A_27_297#_c_570_p N_A_27_297#_c_521_n
+ N_A_27_297#_c_550_p PM_SKY130_FD_SC_HD__NOR4B_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR4B_4%VPWR N_VPWR_M1003_d N_VPWR_M1023_d N_VPWR_M1011_d
+ N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n VPWR
+ N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n
+ N_VPWR_c_579_n PM_SKY130_FD_SC_HD__NOR4B_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR4B_4%A_445_297# N_A_445_297#_M1000_d
+ N_A_445_297#_M1026_d N_A_445_297#_M1001_d N_A_445_297#_M1014_d
+ N_A_445_297#_c_683_n N_A_445_297#_c_684_n N_A_445_297#_c_685_n
+ N_A_445_297#_c_686_n N_A_445_297#_c_687_n N_A_445_297#_c_688_n
+ N_A_445_297#_c_689_n PM_SKY130_FD_SC_HD__NOR4B_4%A_445_297#
x_PM_SKY130_FD_SC_HD__NOR4B_4%A_803_297# N_A_803_297#_M1001_s
+ N_A_803_297#_M1010_s N_A_803_297#_M1032_s N_A_803_297#_M1004_s
+ N_A_803_297#_M1027_s N_A_803_297#_c_760_n N_A_803_297#_c_744_n
+ N_A_803_297#_c_741_n N_A_803_297#_c_790_n N_A_803_297#_c_746_n
+ N_A_803_297#_c_742_n N_A_803_297#_c_751_n N_A_803_297#_c_800_p
+ N_A_803_297#_c_743_n N_A_803_297#_c_756_n N_A_803_297#_c_777_n
+ N_A_803_297#_c_779_n N_A_803_297#_c_781_n
+ PM_SKY130_FD_SC_HD__NOR4B_4%A_803_297#
x_PM_SKY130_FD_SC_HD__NOR4B_4%Y N_Y_M1015_s N_Y_M1022_s N_Y_M1019_d N_Y_M1028_d
+ N_Y_M1012_d N_Y_M1020_d N_Y_M1008_d N_Y_M1017_d N_Y_M1002_d N_Y_M1007_d
+ N_Y_c_824_n N_Y_c_806_n N_Y_c_807_n N_Y_c_835_n N_Y_c_808_n N_Y_c_840_n
+ N_Y_c_809_n N_Y_c_855_n N_Y_c_810_n N_Y_c_870_n N_Y_c_811_n N_Y_c_877_n
+ N_Y_c_812_n N_Y_c_882_n N_Y_c_813_n N_Y_c_814_n N_Y_c_822_n N_Y_c_917_n
+ N_Y_c_815_n N_Y_c_816_n N_Y_c_817_n N_Y_c_818_n N_Y_c_819_n N_Y_c_820_n
+ N_Y_c_923_n N_Y_c_823_n Y PM_SKY130_FD_SC_HD__NOR4B_4%Y
x_PM_SKY130_FD_SC_HD__NOR4B_4%VGND N_VGND_M1015_d N_VGND_M1018_d N_VGND_M1033_d
+ N_VGND_M1024_s N_VGND_M1029_s N_VGND_M1016_s N_VGND_M1025_s N_VGND_M1013_s
+ N_VGND_M1021_s N_VGND_M1009_d N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n
+ N_VGND_c_1010_n N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n
+ N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n
+ N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n
+ N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n N_VGND_c_1025_n
+ N_VGND_c_1026_n N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n
+ N_VGND_c_1030_n VGND N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n
+ N_VGND_c_1034_n N_VGND_c_1035_n PM_SKY130_FD_SC_HD__NOR4B_4%VGND
cc_1 VNB N_A_c_134_n 0.0216231f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_135_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_c_136_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_c_137_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_c_138_n 0.0100386f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.16
cc_6 VNB N_A_c_139_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_7 VNB N_B_c_210_n 0.0160129f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B_c_211_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_9 VNB N_B_c_212_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_10 VNB N_B_c_213_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_11 VNB N_B_c_214_n 0.00882304f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.16
cc_12 VNB N_B_c_215_n 0.0689331f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_13 VNB N_C_c_289_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_C_c_290_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_15 VNB N_C_c_291_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_16 VNB N_C_c_292_n 0.0159885f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_17 VNB N_C_c_293_n 0.00976873f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.16
cc_18 VNB N_C_c_294_n 0.0689265f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_19 VNB N_A_1191_21#_c_368_n 0.0159859f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_1191_21#_c_369_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_1191_21#_c_370_n 0.0157583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_1191_21#_c_371_n 0.019082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_1191_21#_c_372_n 0.00248213f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_24 VNB N_A_1191_21#_c_373_n 0.0094535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_1191_21#_c_374_n 0.00666161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_1191_21#_c_375_n 0.0302972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_1191_21#_c_376_n 0.0592082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB D_N 0.0226975f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_29 VNB N_D_N_c_487_n 0.0383084f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_30 VNB N_D_N_c_488_n 0.0253599f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_31 VNB N_VPWR_c_579_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_806_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_33 VNB N_Y_c_807_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_34 VNB N_Y_c_808_n 0.00429924f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_35 VNB N_Y_c_809_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.18
cc_36 VNB N_Y_c_810_n 0.00898206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_811_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_812_n 0.0045318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_813_n 8.77122e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_814_n 0.0048242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_815_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_816_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_817_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_818_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_819_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_820_n 4.05044e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_1007_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_48 VNB N_VGND_c_1008_n 0.0072727f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_49 VNB N_VGND_c_1009_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_50 VNB N_VGND_c_1010_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_51 VNB N_VGND_c_1011_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.18
cc_52 VNB N_VGND_c_1012_n 0.00358794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1013_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1014_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1015_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1016_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1017_n 0.0115659f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1018_n 0.00737297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1019_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1020_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1021_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1022_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1023_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1024_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1025_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1026_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1027_n 0.016668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1028_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1029_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1030_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1031_n 0.0199727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1032_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1033_n 0.0197313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1034_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1035_n 0.415684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VPB N_A_M1003_g 0.0252519f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_77 VPB N_A_M1005_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_78 VPB N_A_M1023_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_79 VPB N_A_M1030_g 0.0185045f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_80 VPB N_A_c_139_n 0.0108808f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_81 VPB N_B_M1000_g 0.018818f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_82 VPB N_B_M1006_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_83 VPB N_B_M1026_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_84 VPB N_B_M1031_g 0.0252703f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_85 VPB N_B_c_215_n 0.0108798f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_86 VPB N_C_M1001_g 0.0252703f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_87 VPB N_C_M1010_g 0.0182218f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_88 VPB N_C_M1014_g 0.0182218f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_89 VPB N_C_M1032_g 0.0188099f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_90 VPB N_C_c_294_n 0.0108785f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_91 VPB N_A_1191_21#_M1002_g 0.0187789f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_92 VPB N_A_1191_21#_M1004_g 0.0176643f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_93 VPB N_A_1191_21#_M1007_g 0.0181703f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_94 VPB N_A_1191_21#_M1027_g 0.021923f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_95 VPB N_A_1191_21#_c_381_n 0.0028702f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.18
cc_96 VPB N_A_1191_21#_c_382_n 0.0135429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_1191_21#_c_383_n 8.41749e-19 $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.18
cc_98 VPB N_A_1191_21#_c_384_n 0.00897765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_1191_21#_c_375_n 0.0113164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_1191_21#_c_376_n 0.0102181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_D_N_M1011_g 0.0297081f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_102 VPB N_D_N_c_487_n 0.00983391f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_103 VPB N_A_27_297#_c_515_n 0.0327625f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_104 VPB N_A_27_297#_c_516_n 0.00226814f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_105 VPB N_A_27_297#_c_517_n 0.0152931f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_106 VPB N_A_27_297#_c_518_n 0.00240493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_27_297#_c_519_n 0.00414042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_27_297#_c_520_n 0.0014617f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=1.16
cc_109 VPB N_A_27_297#_c_521_n 0.00204609f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.18
cc_110 VPB N_VPWR_c_580_n 0.00428214f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_111 VPB N_VPWR_c_581_n 0.00454762f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_112 VPB N_VPWR_c_582_n 0.01154f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_113 VPB N_VPWR_c_583_n 0.00789007f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_114 VPB N_VPWR_c_584_n 0.0178658f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_115 VPB N_VPWR_c_585_n 0.0163782f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_116 VPB N_VPWR_c_586_n 0.156607f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_117 VPB N_VPWR_c_587_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_588_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.135 $Y2=1.18
cc_119 VPB N_VPWR_c_579_n 0.0682187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_445_297#_c_683_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.995
cc_121 VPB N_A_445_297#_c_684_n 0.0199604f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_122 VPB N_A_445_297#_c_685_n 0.00235082f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_123 VPB N_A_445_297#_c_686_n 0.00225182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_445_297#_c_687_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_445_297#_c_688_n 0.00202679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_445_297#_c_689_n 0.002258f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_127 VPB N_A_803_297#_c_741_n 0.0014617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_803_297#_c_742_n 0.004421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_803_297#_c_743_n 0.00138574f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=1.16
cc_130 VPB N_Y_c_813_n 0.00127133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_Y_c_822_n 0.00268792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_Y_c_823_n 0.00228462f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 N_A_c_137_n N_B_c_210_n 0.0195974f $X=1.73 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 N_A_M1030_g N_B_M1000_g 0.0195974f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_135 N_A_c_138_n N_B_c_214_n 0.0121231f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_139_n N_B_c_214_n 2.62535e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_138_n N_B_c_215_n 2.62535e-19 $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_c_139_n N_B_c_215_n 0.0195974f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_M1003_g N_A_27_297#_c_515_n 0.0102794f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_M1005_g N_A_27_297#_c_515_n 6.39954e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_A_27_297#_c_516_n 0.0107189f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_M1005_g N_A_27_297#_c_516_n 0.0132714f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A_c_138_n N_A_27_297#_c_516_n 0.0388745f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_c_139_n N_A_27_297#_c_516_n 0.00211509f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_M1003_g N_A_27_297#_c_517_n 0.0014856f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_c_138_n N_A_27_297#_c_517_n 0.002319f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_M1023_g N_A_27_297#_c_518_n 0.0132273f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A_M1030_g N_A_27_297#_c_518_n 0.0132131f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A_c_138_n N_A_27_297#_c_518_n 0.0409754f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_139_n N_A_27_297#_c_518_n 0.00211509f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_c_138_n N_A_27_297#_c_521_n 0.0204549f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_c_139_n N_A_27_297#_c_521_n 0.00220041f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_M1003_g N_VPWR_c_580_n 0.00274642f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_M1005_g N_VPWR_c_580_n 0.00155565f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_M1023_g N_VPWR_c_581_n 0.00157837f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_156 N_A_M1030_g N_VPWR_c_581_n 0.00302074f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_M1003_g N_VPWR_c_584_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_158 N_A_M1005_g N_VPWR_c_585_n 0.00585385f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_M1023_g N_VPWR_c_585_n 0.00585385f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_160 N_A_M1030_g N_VPWR_c_586_n 0.00585385f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_161 N_A_M1003_g N_VPWR_c_579_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_162 N_A_M1005_g N_VPWR_c_579_n 0.0104367f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A_M1023_g N_VPWR_c_579_n 0.0104367f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_M1030_g N_VPWR_c_579_n 0.010464f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A_c_134_n N_Y_c_824_n 0.00539651f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_135_n N_Y_c_824_n 0.00630972f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_136_n N_Y_c_824_n 5.22228e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_135_n N_Y_c_806_n 0.00870364f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_136_n N_Y_c_806_n 0.00870364f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_138_n N_Y_c_806_n 0.0362443f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_139_n N_Y_c_806_n 0.00222133f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_c_134_n N_Y_c_807_n 0.00299247f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_135_n N_Y_c_807_n 0.00113286f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_c_138_n N_Y_c_807_n 0.0266272f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_c_139_n N_Y_c_807_n 0.00230339f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_c_135_n N_Y_c_835_n 5.22228e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_136_n N_Y_c_835_n 0.00630972f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_137_n N_Y_c_835_n 0.00630972f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_137_n N_Y_c_808_n 0.00865686f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_138_n N_Y_c_808_n 0.00826974f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_c_137_n N_Y_c_840_n 5.22228e-19 $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_c_136_n N_Y_c_815_n 0.00113286f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_137_n N_Y_c_815_n 0.00113286f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_138_n N_Y_c_815_n 0.0266272f $X=1.58 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_c_139_n N_Y_c_815_n 0.00230339f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_134_n N_VGND_c_1008_n 0.00338128f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_135_n N_VGND_c_1009_n 0.00146448f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_136_n N_VGND_c_1009_n 0.00146448f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_137_n N_VGND_c_1010_n 0.00146448f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_134_n N_VGND_c_1019_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_135_n N_VGND_c_1019_n 0.00423334f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_136_n N_VGND_c_1021_n 0.00423334f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_137_n N_VGND_c_1021_n 0.00423334f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_134_n N_VGND_c_1035_n 0.0104557f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_135_n N_VGND_c_1035_n 0.0057163f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_136_n N_VGND_c_1035_n 0.0057163f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_137_n N_VGND_c_1035_n 0.0057435f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B_c_214_n N_C_c_293_n 0.0155079f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B_c_215_n N_C_c_293_n 9.30294e-19 $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_214_n N_C_c_294_n 8.91304e-19 $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B_M1000_g N_A_27_297#_c_519_n 2.57315e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_202 N_B_M1000_g N_A_27_297#_c_537_n 0.0121747f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_203 N_B_M1006_g N_A_27_297#_c_537_n 0.00984328f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_204 N_B_M1026_g N_A_27_297#_c_520_n 0.00984328f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_205 N_B_M1031_g N_A_27_297#_c_520_n 0.00988743f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_206 N_B_M1000_g N_VPWR_c_586_n 0.00357877f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_207 N_B_M1006_g N_VPWR_c_586_n 0.00357877f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_208 N_B_M1026_g N_VPWR_c_586_n 0.00357877f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_209 N_B_M1031_g N_VPWR_c_586_n 0.00357877f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B_M1000_g N_VPWR_c_579_n 0.00525237f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B_M1006_g N_VPWR_c_579_n 0.00522516f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B_M1026_g N_VPWR_c_579_n 0.00522516f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B_M1031_g N_VPWR_c_579_n 0.00655123f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B_M1006_g N_A_445_297#_c_683_n 0.0109258f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_215 N_B_M1026_g N_A_445_297#_c_683_n 0.01094f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_216 N_B_c_214_n N_A_445_297#_c_683_n 0.0416643f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B_c_215_n N_A_445_297#_c_683_n 0.00211509f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_218 N_B_M1031_g N_A_445_297#_c_684_n 0.0130871f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_219 N_B_c_214_n N_A_445_297#_c_684_n 0.0313043f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B_M1000_g N_A_445_297#_c_686_n 2.57315e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_221 N_B_c_214_n N_A_445_297#_c_686_n 0.0204292f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_c_215_n N_A_445_297#_c_686_n 0.00219557f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B_c_214_n N_A_445_297#_c_687_n 0.0204292f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B_c_215_n N_A_445_297#_c_687_n 0.00219557f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_225 N_B_c_210_n N_Y_c_835_n 5.22228e-19 $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_210_n N_Y_c_808_n 0.00865686f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B_c_214_n N_Y_c_808_n 0.00826974f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_228 N_B_c_210_n N_Y_c_840_n 0.00630972f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_211_n N_Y_c_840_n 0.00630972f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_212_n N_Y_c_840_n 5.22228e-19 $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B_c_211_n N_Y_c_809_n 0.00870364f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B_c_212_n N_Y_c_809_n 0.00870364f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_214_n N_Y_c_809_n 0.0362443f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_234 N_B_c_215_n N_Y_c_809_n 0.00222133f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B_c_211_n N_Y_c_855_n 5.22228e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_212_n N_Y_c_855_n 0.00630972f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_213_n N_Y_c_855_n 0.0109565f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_213_n N_Y_c_810_n 0.0109318f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B_c_214_n N_Y_c_810_n 0.0286372f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B_c_210_n N_Y_c_816_n 0.00113286f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_211_n N_Y_c_816_n 0.00113286f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B_c_214_n N_Y_c_816_n 0.0266272f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B_c_215_n N_Y_c_816_n 0.00230339f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_244 N_B_c_212_n N_Y_c_817_n 0.00113286f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_245 N_B_c_213_n N_Y_c_817_n 0.00113286f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B_c_214_n N_Y_c_817_n 0.0266272f $X=3.26 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B_c_215_n N_Y_c_817_n 0.00230339f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B_c_210_n N_VGND_c_1010_n 0.00146448f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_211_n N_VGND_c_1011_n 0.00146448f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B_c_212_n N_VGND_c_1011_n 0.00146339f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_c_210_n N_VGND_c_1023_n 0.00423334f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B_c_211_n N_VGND_c_1023_n 0.00423334f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B_c_212_n N_VGND_c_1032_n 0.00423334f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B_c_213_n N_VGND_c_1032_n 0.00423334f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_255 N_B_c_213_n N_VGND_c_1033_n 0.00335921f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_256 N_B_c_210_n N_VGND_c_1035_n 0.0057435f $X=2.15 $Y=0.995 $X2=0 $Y2=0
cc_257 N_B_c_211_n N_VGND_c_1035_n 0.0057163f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B_c_212_n N_VGND_c_1035_n 0.0057163f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_259 N_B_c_213_n N_VGND_c_1035_n 0.0070399f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_260 N_C_c_292_n N_A_1191_21#_c_368_n 0.0190321f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_261 N_C_M1032_g N_A_1191_21#_M1002_g 0.0190321f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_262 N_C_c_293_n N_A_1191_21#_c_376_n 9.94048e-19 $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_263 N_C_c_294_n N_A_1191_21#_c_376_n 0.0190321f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_264 N_C_M1001_g N_VPWR_c_586_n 0.00357877f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_265 N_C_M1010_g N_VPWR_c_586_n 0.00357877f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_266 N_C_M1014_g N_VPWR_c_586_n 0.00357877f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_267 N_C_M1032_g N_VPWR_c_586_n 0.00357877f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_268 N_C_M1001_g N_VPWR_c_579_n 0.00655123f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_269 N_C_M1010_g N_VPWR_c_579_n 0.00522516f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_270 N_C_M1014_g N_VPWR_c_579_n 0.00522516f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_271 N_C_M1032_g N_VPWR_c_579_n 0.00525237f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_272 N_C_M1001_g N_A_445_297#_c_684_n 0.0130871f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_273 N_C_c_293_n N_A_445_297#_c_684_n 0.0332175f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_274 N_C_M1010_g N_A_445_297#_c_685_n 0.01094f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_275 N_C_M1014_g N_A_445_297#_c_685_n 0.0109258f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_276 N_C_c_293_n N_A_445_297#_c_685_n 0.0416643f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_277 N_C_c_294_n N_A_445_297#_c_685_n 0.00211509f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_278 N_C_c_293_n N_A_445_297#_c_688_n 0.0204292f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_279 N_C_c_294_n N_A_445_297#_c_688_n 0.00219557f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_280 N_C_M1032_g N_A_445_297#_c_689_n 2.5798e-19 $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_281 N_C_c_293_n N_A_445_297#_c_689_n 0.0204292f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_282 N_C_c_294_n N_A_445_297#_c_689_n 0.00219557f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_283 N_C_M1001_g N_A_803_297#_c_744_n 0.00988743f $X=4.35 $Y=1.985 $X2=0 $Y2=0
cc_284 N_C_M1010_g N_A_803_297#_c_744_n 0.00984328f $X=4.77 $Y=1.985 $X2=0 $Y2=0
cc_285 N_C_M1014_g N_A_803_297#_c_746_n 0.00988743f $X=5.19 $Y=1.985 $X2=0 $Y2=0
cc_286 N_C_M1032_g N_A_803_297#_c_746_n 0.0121747f $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_287 N_C_M1032_g N_A_803_297#_c_742_n 2.30871e-19 $X=5.61 $Y=1.985 $X2=0 $Y2=0
cc_288 N_C_c_289_n N_Y_c_810_n 0.0109318f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_289 N_C_c_293_n N_Y_c_810_n 0.0305587f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_290 N_C_c_289_n N_Y_c_870_n 0.0109565f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_291 N_C_c_290_n N_Y_c_870_n 0.00630972f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_292 N_C_c_291_n N_Y_c_870_n 5.22228e-19 $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_293 N_C_c_290_n N_Y_c_811_n 0.00870364f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C_c_291_n N_Y_c_811_n 0.00870364f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_c_293_n N_Y_c_811_n 0.0362443f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_296 N_C_c_294_n N_Y_c_811_n 0.00222133f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_297 N_C_c_290_n N_Y_c_877_n 5.22228e-19 $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_c_291_n N_Y_c_877_n 0.00630972f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_299 N_C_c_292_n N_Y_c_877_n 0.00630972f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_292_n N_Y_c_812_n 0.00865686f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_293_n N_Y_c_812_n 0.00826974f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_302 N_C_c_292_n N_Y_c_882_n 5.22228e-19 $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_303 N_C_c_293_n N_Y_c_813_n 0.00785191f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_304 N_C_c_294_n N_Y_c_813_n 8.73873e-19 $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_305 N_C_c_289_n N_Y_c_818_n 0.00113286f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_306 N_C_c_290_n N_Y_c_818_n 0.00113286f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_307 N_C_c_293_n N_Y_c_818_n 0.0266272f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_308 N_C_c_294_n N_Y_c_818_n 0.00230339f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_309 N_C_c_291_n N_Y_c_819_n 0.00113286f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_310 N_C_c_292_n N_Y_c_819_n 0.00113286f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_311 N_C_c_293_n N_Y_c_819_n 0.0266272f $X=5.46 $Y=1.16 $X2=0 $Y2=0
cc_312 N_C_c_294_n N_Y_c_819_n 0.00230339f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_313 N_C_c_290_n N_VGND_c_1012_n 0.00146339f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_314 N_C_c_291_n N_VGND_c_1012_n 0.00146448f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_315 N_C_c_291_n N_VGND_c_1013_n 0.00423334f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_316 N_C_c_292_n N_VGND_c_1013_n 0.00423334f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_317 N_C_c_292_n N_VGND_c_1014_n 0.00146448f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_318 N_C_c_289_n N_VGND_c_1025_n 0.00423334f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_319 N_C_c_290_n N_VGND_c_1025_n 0.00423334f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_320 N_C_c_289_n N_VGND_c_1033_n 0.00335921f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_321 N_C_c_289_n N_VGND_c_1035_n 0.0070399f $X=4.35 $Y=0.995 $X2=0 $Y2=0
cc_322 N_C_c_290_n N_VGND_c_1035_n 0.0057163f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_323 N_C_c_291_n N_VGND_c_1035_n 0.0057163f $X=5.19 $Y=0.995 $X2=0 $Y2=0
cc_324 N_C_c_292_n N_VGND_c_1035_n 0.0057435f $X=5.61 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_1191_21#_c_381_n N_D_N_M1011_g 0.00307757f $X=7.555 $Y=1.455 $X2=0
+ $Y2=0
cc_326 N_A_1191_21#_c_382_n N_D_N_M1011_g 0.0030022f $X=7.85 $Y=1.54 $X2=0 $Y2=0
cc_327 N_A_1191_21#_c_384_n N_D_N_M1011_g 0.00946465f $X=8.02 $Y=1.63 $X2=0
+ $Y2=0
cc_328 N_A_1191_21#_c_382_n D_N 0.0314793f $X=7.85 $Y=1.54 $X2=0 $Y2=0
cc_329 N_A_1191_21#_c_373_n D_N 0.0284697f $X=7.997 $Y=0.735 $X2=0 $Y2=0
cc_330 N_A_1191_21#_c_396_p D_N 0.0185422f $X=7.555 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_1191_21#_c_375_n D_N 0.00244543f $X=7.555 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_1191_21#_c_372_n N_D_N_c_487_n 4.45113e-19 $X=7.555 $Y=1.075 $X2=0
+ $Y2=0
cc_333 N_A_1191_21#_c_381_n N_D_N_c_487_n 2.21427e-19 $X=7.555 $Y=1.455 $X2=0
+ $Y2=0
cc_334 N_A_1191_21#_c_375_n N_D_N_c_487_n 0.00924724f $X=7.555 $Y=1.16 $X2=0
+ $Y2=0
cc_335 N_A_1191_21#_c_372_n N_D_N_c_488_n 0.00213537f $X=7.555 $Y=1.075 $X2=0
+ $Y2=0
cc_336 N_A_1191_21#_c_373_n N_D_N_c_488_n 0.00285661f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_337 N_A_1191_21#_c_374_n N_D_N_c_488_n 0.00560573f $X=8.02 $Y=0.39 $X2=0
+ $Y2=0
cc_338 N_A_1191_21#_c_382_n N_VPWR_c_583_n 0.00836315f $X=7.85 $Y=1.54 $X2=0
+ $Y2=0
cc_339 N_A_1191_21#_M1002_g N_VPWR_c_586_n 0.00357877f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_340 N_A_1191_21#_M1004_g N_VPWR_c_586_n 0.00357877f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_1191_21#_M1007_g N_VPWR_c_586_n 0.00357877f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_1191_21#_M1027_g N_VPWR_c_586_n 0.00357877f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_1191_21#_c_384_n N_VPWR_c_586_n 0.0213966f $X=8.02 $Y=1.63 $X2=0
+ $Y2=0
cc_344 N_A_1191_21#_M1011_s N_VPWR_c_579_n 0.00209319f $X=7.895 $Y=1.485 $X2=0
+ $Y2=0
cc_345 N_A_1191_21#_M1002_g N_VPWR_c_579_n 0.00525237f $X=6.03 $Y=1.985 $X2=0
+ $Y2=0
cc_346 N_A_1191_21#_M1004_g N_VPWR_c_579_n 0.00522516f $X=6.45 $Y=1.985 $X2=0
+ $Y2=0
cc_347 N_A_1191_21#_M1007_g N_VPWR_c_579_n 0.00522516f $X=6.87 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_1191_21#_M1027_g N_VPWR_c_579_n 0.00655123f $X=7.29 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_1191_21#_c_384_n N_VPWR_c_579_n 0.0126193f $X=8.02 $Y=1.63 $X2=0
+ $Y2=0
cc_350 N_A_1191_21#_c_383_n N_A_803_297#_M1027_s 0.0041468f $X=7.64 $Y=1.54
+ $X2=0 $Y2=0
cc_351 N_A_1191_21#_M1002_g N_A_803_297#_c_742_n 2.30871e-19 $X=6.03 $Y=1.985
+ $X2=0 $Y2=0
cc_352 N_A_1191_21#_M1002_g N_A_803_297#_c_751_n 0.0121747f $X=6.03 $Y=1.985
+ $X2=0 $Y2=0
cc_353 N_A_1191_21#_M1004_g N_A_803_297#_c_751_n 0.00985663f $X=6.45 $Y=1.985
+ $X2=0 $Y2=0
cc_354 N_A_1191_21#_M1007_g N_A_803_297#_c_743_n 0.00984328f $X=6.87 $Y=1.985
+ $X2=0 $Y2=0
cc_355 N_A_1191_21#_M1027_g N_A_803_297#_c_743_n 0.0121747f $X=7.29 $Y=1.985
+ $X2=0 $Y2=0
cc_356 N_A_1191_21#_c_384_n N_A_803_297#_c_743_n 0.0120455f $X=8.02 $Y=1.63
+ $X2=0 $Y2=0
cc_357 N_A_1191_21#_c_423_p N_A_803_297#_c_756_n 0.00227909f $X=7.47 $Y=1.18
+ $X2=0 $Y2=0
cc_358 N_A_1191_21#_c_383_n N_A_803_297#_c_756_n 0.0139284f $X=7.64 $Y=1.54
+ $X2=0 $Y2=0
cc_359 N_A_1191_21#_c_384_n N_A_803_297#_c_756_n 0.0327602f $X=8.02 $Y=1.63
+ $X2=0 $Y2=0
cc_360 N_A_1191_21#_c_375_n N_A_803_297#_c_756_n 0.00225697f $X=7.555 $Y=1.16
+ $X2=0 $Y2=0
cc_361 N_A_1191_21#_c_368_n N_Y_c_877_n 5.22228e-19 $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A_1191_21#_c_368_n N_Y_c_812_n 0.0123222f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A_1191_21#_c_368_n N_Y_c_882_n 0.00630972f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_1191_21#_c_369_n N_Y_c_882_n 0.00630972f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A_1191_21#_c_370_n N_Y_c_882_n 5.22228e-19 $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A_1191_21#_c_368_n N_Y_c_813_n 0.00256954f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A_1191_21#_M1002_g N_Y_c_813_n 0.00372438f $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A_1191_21#_c_369_n N_Y_c_813_n 0.0028766f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A_1191_21#_M1004_g N_Y_c_813_n 0.00418415f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A_1191_21#_c_370_n N_Y_c_813_n 4.91375e-19 $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_1191_21#_M1007_g N_Y_c_813_n 7.13641e-19 $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_372 N_A_1191_21#_c_423_p N_Y_c_813_n 0.0166745f $X=7.47 $Y=1.18 $X2=0 $Y2=0
cc_373 N_A_1191_21#_c_376_n N_Y_c_813_n 0.0290684f $X=7.365 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_1191_21#_c_369_n N_Y_c_814_n 0.0060413f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A_1191_21#_c_370_n N_Y_c_814_n 0.00982493f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A_1191_21#_c_371_n N_Y_c_814_n 0.00294361f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A_1191_21#_c_423_p N_Y_c_814_n 0.0465735f $X=7.47 $Y=1.18 $X2=0 $Y2=0
cc_378 N_A_1191_21#_c_373_n N_Y_c_814_n 0.0118927f $X=7.997 $Y=0.735 $X2=0 $Y2=0
cc_379 N_A_1191_21#_c_374_n N_Y_c_814_n 3.40613e-19 $X=8.02 $Y=0.39 $X2=0 $Y2=0
cc_380 N_A_1191_21#_c_376_n N_Y_c_814_n 0.00461638f $X=7.365 $Y=1.16 $X2=0 $Y2=0
cc_381 N_A_1191_21#_M1004_g N_Y_c_822_n 0.00603426f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A_1191_21#_M1007_g N_Y_c_822_n 0.0108817f $X=6.87 $Y=1.985 $X2=0 $Y2=0
cc_383 N_A_1191_21#_c_423_p N_Y_c_822_n 0.0226482f $X=7.47 $Y=1.18 $X2=0 $Y2=0
cc_384 N_A_1191_21#_c_376_n N_Y_c_822_n 0.00219918f $X=7.365 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A_1191_21#_c_369_n N_Y_c_917_n 5.22228e-19 $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A_1191_21#_c_370_n N_Y_c_917_n 0.00630972f $X=6.87 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A_1191_21#_c_371_n N_Y_c_917_n 0.00701638f $X=7.29 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A_1191_21#_c_374_n N_Y_c_917_n 0.00548956f $X=8.02 $Y=0.39 $X2=0 $Y2=0
cc_389 N_A_1191_21#_c_368_n N_Y_c_820_n 0.00221107f $X=6.03 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A_1191_21#_c_369_n N_Y_c_820_n 0.00324953f $X=6.45 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A_1191_21#_M1002_g N_Y_c_923_n 2.5798e-19 $X=6.03 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A_1191_21#_M1004_g N_Y_c_923_n 0.00441257f $X=6.45 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A_1191_21#_M1027_g N_Y_c_823_n 3.17833e-19 $X=7.29 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A_1191_21#_c_423_p N_Y_c_823_n 0.0204292f $X=7.47 $Y=1.18 $X2=0 $Y2=0
cc_395 N_A_1191_21#_c_383_n N_Y_c_823_n 0.00659639f $X=7.64 $Y=1.54 $X2=0 $Y2=0
cc_396 N_A_1191_21#_c_376_n N_Y_c_823_n 0.00219557f $X=7.365 $Y=1.16 $X2=0 $Y2=0
cc_397 N_A_1191_21#_c_373_n N_VGND_M1021_s 0.00408724f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_398 N_A_1191_21#_c_368_n N_VGND_c_1014_n 0.00146448f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_399 N_A_1191_21#_c_369_n N_VGND_c_1015_n 0.00146448f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_400 N_A_1191_21#_c_370_n N_VGND_c_1015_n 0.00146448f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_401 N_A_1191_21#_c_371_n N_VGND_c_1016_n 0.00316354f $X=7.29 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_A_1191_21#_c_423_p N_VGND_c_1016_n 0.00167341f $X=7.47 $Y=1.18 $X2=0
+ $Y2=0
cc_403 N_A_1191_21#_c_373_n N_VGND_c_1016_n 0.00851553f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_404 N_A_1191_21#_c_374_n N_VGND_c_1016_n 0.019325f $X=8.02 $Y=0.39 $X2=0
+ $Y2=0
cc_405 N_A_1191_21#_c_375_n N_VGND_c_1016_n 0.00107514f $X=7.555 $Y=1.16 $X2=0
+ $Y2=0
cc_406 N_A_1191_21#_c_373_n N_VGND_c_1018_n 0.00784313f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_407 N_A_1191_21#_c_368_n N_VGND_c_1027_n 0.00423334f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_408 N_A_1191_21#_c_369_n N_VGND_c_1027_n 0.00423279f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_409 N_A_1191_21#_c_370_n N_VGND_c_1029_n 0.00423334f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_410 N_A_1191_21#_c_371_n N_VGND_c_1029_n 0.00541359f $X=7.29 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_A_1191_21#_c_373_n N_VGND_c_1031_n 0.00335436f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_412 N_A_1191_21#_c_374_n N_VGND_c_1031_n 0.0237059f $X=8.02 $Y=0.39 $X2=0
+ $Y2=0
cc_413 N_A_1191_21#_M1009_s N_VGND_c_1035_n 0.00209319f $X=7.895 $Y=0.235 $X2=0
+ $Y2=0
cc_414 N_A_1191_21#_c_368_n N_VGND_c_1035_n 0.0057435f $X=6.03 $Y=0.995 $X2=0
+ $Y2=0
cc_415 N_A_1191_21#_c_369_n N_VGND_c_1035_n 0.0057153f $X=6.45 $Y=0.995 $X2=0
+ $Y2=0
cc_416 N_A_1191_21#_c_370_n N_VGND_c_1035_n 0.0057163f $X=6.87 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A_1191_21#_c_371_n N_VGND_c_1035_n 0.0108276f $X=7.29 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A_1191_21#_c_373_n N_VGND_c_1035_n 0.00642555f $X=7.997 $Y=0.735 $X2=0
+ $Y2=0
cc_419 N_A_1191_21#_c_374_n N_VGND_c_1035_n 0.0140329f $X=8.02 $Y=0.39 $X2=0
+ $Y2=0
cc_420 N_D_N_M1011_g N_VPWR_c_583_n 0.00513607f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_421 D_N N_VPWR_c_583_n 0.0187446f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_422 N_D_N_c_487_n N_VPWR_c_583_n 0.00498759f $X=8.395 $Y=1.16 $X2=0 $Y2=0
cc_423 N_D_N_M1011_g N_VPWR_c_586_n 0.00541359f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_424 N_D_N_M1011_g N_VPWR_c_579_n 0.0118181f $X=8.23 $Y=1.985 $X2=0 $Y2=0
cc_425 N_D_N_c_488_n N_VGND_c_1016_n 0.00194637f $X=8.357 $Y=0.995 $X2=0 $Y2=0
cc_426 D_N N_VGND_c_1018_n 0.0187437f $X=8.43 $Y=1.105 $X2=0 $Y2=0
cc_427 N_D_N_c_487_n N_VGND_c_1018_n 0.00523789f $X=8.395 $Y=1.16 $X2=0 $Y2=0
cc_428 N_D_N_c_488_n N_VGND_c_1018_n 0.00493171f $X=8.357 $Y=0.995 $X2=0 $Y2=0
cc_429 N_D_N_c_488_n N_VGND_c_1031_n 0.00540385f $X=8.357 $Y=0.995 $X2=0 $Y2=0
cc_430 N_D_N_c_488_n N_VGND_c_1035_n 0.011772f $X=8.357 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A_27_297#_c_516_n N_VPWR_M1003_d 0.00165831f $X=0.975 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_432 N_A_27_297#_c_518_n N_VPWR_M1023_d 0.00165831f $X=1.815 $Y=1.54 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_c_516_n N_VPWR_c_580_n 0.0126919f $X=0.975 $Y=1.54 $X2=0
+ $Y2=0
cc_434 N_A_27_297#_c_518_n N_VPWR_c_581_n 0.0126919f $X=1.815 $Y=1.54 $X2=0
+ $Y2=0
cc_435 N_A_27_297#_c_515_n N_VPWR_c_584_n 0.0210382f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_436 N_A_27_297#_c_546_p N_VPWR_c_585_n 0.0142343f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_437 N_A_27_297#_c_547_p N_VPWR_c_586_n 0.0143053f $X=1.94 $Y=2.295 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_c_537_n N_VPWR_c_586_n 0.0330174f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_c_520_n N_VPWR_c_586_n 0.0489446f $X=3.495 $Y=2.38 $X2=0
+ $Y2=0
cc_440 N_A_27_297#_c_550_p N_VPWR_c_586_n 0.0142933f $X=2.78 $Y=2.38 $X2=0 $Y2=0
cc_441 N_A_27_297#_M1003_s N_VPWR_c_579_n 0.00209319f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_442 N_A_27_297#_M1005_s N_VPWR_c_579_n 0.00284632f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_443 N_A_27_297#_M1030_s N_VPWR_c_579_n 0.00246446f $X=1.805 $Y=1.485 $X2=0
+ $Y2=0
cc_444 N_A_27_297#_M1006_s N_VPWR_c_579_n 0.00215203f $X=2.645 $Y=1.485 $X2=0
+ $Y2=0
cc_445 N_A_27_297#_M1031_s N_VPWR_c_579_n 0.0020932f $X=3.485 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_A_27_297#_c_515_n N_VPWR_c_579_n 0.0124268f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_447 N_A_27_297#_c_546_p N_VPWR_c_579_n 0.00955092f $X=1.1 $Y=2.3 $X2=0 $Y2=0
cc_448 N_A_27_297#_c_547_p N_VPWR_c_579_n 0.00962794f $X=1.94 $Y=2.295 $X2=0
+ $Y2=0
cc_449 N_A_27_297#_c_537_n N_VPWR_c_579_n 0.0204627f $X=2.655 $Y=2.38 $X2=0
+ $Y2=0
cc_450 N_A_27_297#_c_520_n N_VPWR_c_579_n 0.0300869f $X=3.495 $Y=2.38 $X2=0
+ $Y2=0
cc_451 N_A_27_297#_c_550_p N_VPWR_c_579_n 0.00962421f $X=2.78 $Y=2.38 $X2=0
+ $Y2=0
cc_452 N_A_27_297#_c_537_n N_A_445_297#_M1000_d 0.00312348f $X=2.655 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_453 N_A_27_297#_c_520_n N_A_445_297#_M1026_d 0.00312348f $X=3.495 $Y=2.38
+ $X2=0 $Y2=0
cc_454 N_A_27_297#_M1006_s N_A_445_297#_c_683_n 0.00165831f $X=2.645 $Y=1.485
+ $X2=0 $Y2=0
cc_455 N_A_27_297#_c_537_n N_A_445_297#_c_683_n 0.00320918f $X=2.655 $Y=2.38
+ $X2=0 $Y2=0
cc_456 N_A_27_297#_c_566_p N_A_445_297#_c_683_n 0.0126766f $X=2.78 $Y=1.96 $X2=0
+ $Y2=0
cc_457 N_A_27_297#_c_520_n N_A_445_297#_c_683_n 0.00320918f $X=3.495 $Y=2.38
+ $X2=0 $Y2=0
cc_458 N_A_27_297#_M1031_s N_A_445_297#_c_684_n 0.00276279f $X=3.485 $Y=1.485
+ $X2=0 $Y2=0
cc_459 N_A_27_297#_c_520_n N_A_445_297#_c_684_n 0.00320918f $X=3.495 $Y=2.38
+ $X2=0 $Y2=0
cc_460 N_A_27_297#_c_570_p N_A_445_297#_c_684_n 0.0164145f $X=3.62 $Y=1.96 $X2=0
+ $Y2=0
cc_461 N_A_27_297#_c_519_n N_A_445_297#_c_686_n 0.00271526f $X=1.94 $Y=1.625
+ $X2=0 $Y2=0
cc_462 N_A_27_297#_c_537_n N_A_445_297#_c_686_n 0.0118729f $X=2.655 $Y=2.38
+ $X2=0 $Y2=0
cc_463 N_A_27_297#_c_520_n N_A_445_297#_c_687_n 0.0118729f $X=3.495 $Y=2.38
+ $X2=0 $Y2=0
cc_464 N_A_27_297#_c_570_p N_A_803_297#_c_760_n 0.027317f $X=3.62 $Y=1.96 $X2=0
+ $Y2=0
cc_465 N_A_27_297#_c_520_n N_A_803_297#_c_741_n 0.0108671f $X=3.495 $Y=2.38
+ $X2=0 $Y2=0
cc_466 N_A_27_297#_c_518_n N_Y_c_808_n 3.18413e-19 $X=1.815 $Y=1.54 $X2=0 $Y2=0
cc_467 N_A_27_297#_c_519_n N_Y_c_808_n 0.00936521f $X=1.94 $Y=1.625 $X2=0 $Y2=0
cc_468 N_A_27_297#_c_517_n N_VGND_c_1008_n 0.00684525f $X=0.425 $Y=1.54 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_579_n N_A_445_297#_M1000_d 0.00216833f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_470 N_VPWR_c_579_n N_A_445_297#_M1026_d 0.00216833f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_579_n N_A_445_297#_M1001_d 0.00216833f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_579_n N_A_445_297#_M1014_d 0.00216833f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_579_n N_A_803_297#_M1001_s 0.0020932f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_474 N_VPWR_c_579_n N_A_803_297#_M1010_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_579_n N_A_803_297#_M1032_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_579_n N_A_803_297#_M1004_s 0.00215203f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_579_n N_A_803_297#_M1027_s 0.0020932f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_586_n N_A_803_297#_c_744_n 0.0330174f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_579_n N_A_803_297#_c_744_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_586_n N_A_803_297#_c_741_n 0.0159273f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_579_n N_A_803_297#_c_741_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_586_n N_A_803_297#_c_746_n 0.0330174f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_579_n N_A_803_297#_c_746_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_586_n N_A_803_297#_c_751_n 0.0330174f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_579_n N_A_803_297#_c_751_n 0.0204627f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_586_n N_A_803_297#_c_743_n 0.0489446f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_579_n N_A_803_297#_c_743_n 0.0300869f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_586_n N_A_803_297#_c_777_n 0.0142933f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_579_n N_A_803_297#_c_777_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_586_n N_A_803_297#_c_779_n 0.0143053f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_579_n N_A_803_297#_c_779_n 0.00961749f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_586_n N_A_803_297#_c_781_n 0.0142933f $X=8.355 $Y=2.72 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_579_n N_A_803_297#_c_781_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_579_n N_Y_M1002_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_c_579_n N_Y_M1007_d 0.00216833f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_496 N_A_445_297#_c_684_n N_A_803_297#_M1001_s 0.00276279f $X=4.435 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_497 N_A_445_297#_c_685_n N_A_803_297#_M1010_s 0.00165831f $X=5.275 $Y=1.54
+ $X2=0 $Y2=0
cc_498 N_A_445_297#_c_684_n N_A_803_297#_c_760_n 0.0164145f $X=4.435 $Y=1.54
+ $X2=0 $Y2=0
cc_499 N_A_445_297#_M1001_d N_A_803_297#_c_744_n 0.00312348f $X=4.425 $Y=1.485
+ $X2=0 $Y2=0
cc_500 N_A_445_297#_c_684_n N_A_803_297#_c_744_n 0.00320918f $X=4.435 $Y=1.54
+ $X2=0 $Y2=0
cc_501 N_A_445_297#_c_685_n N_A_803_297#_c_744_n 0.00320918f $X=5.275 $Y=1.54
+ $X2=0 $Y2=0
cc_502 N_A_445_297#_c_688_n N_A_803_297#_c_744_n 0.0118729f $X=4.56 $Y=1.62
+ $X2=0 $Y2=0
cc_503 N_A_445_297#_c_685_n N_A_803_297#_c_790_n 0.0126766f $X=5.275 $Y=1.54
+ $X2=0 $Y2=0
cc_504 N_A_445_297#_M1014_d N_A_803_297#_c_746_n 0.00312348f $X=5.265 $Y=1.485
+ $X2=0 $Y2=0
cc_505 N_A_445_297#_c_685_n N_A_803_297#_c_746_n 0.00320918f $X=5.275 $Y=1.54
+ $X2=0 $Y2=0
cc_506 N_A_445_297#_c_689_n N_A_803_297#_c_746_n 0.0118729f $X=5.4 $Y=1.62 $X2=0
+ $Y2=0
cc_507 N_A_445_297#_c_689_n N_A_803_297#_c_742_n 0.00251363f $X=5.4 $Y=1.62
+ $X2=0 $Y2=0
cc_508 N_A_445_297#_c_684_n N_Y_c_810_n 0.00787473f $X=4.435 $Y=1.54 $X2=0 $Y2=0
cc_509 N_A_803_297#_c_751_n N_Y_M1002_d 0.00312348f $X=6.535 $Y=2.38 $X2=0 $Y2=0
cc_510 N_A_803_297#_c_743_n N_Y_M1007_d 0.00312348f $X=7.375 $Y=2.38 $X2=0 $Y2=0
cc_511 N_A_803_297#_c_742_n N_Y_c_812_n 0.00929029f $X=5.82 $Y=1.62 $X2=0 $Y2=0
cc_512 N_A_803_297#_M1004_s N_Y_c_822_n 0.00165831f $X=6.525 $Y=1.485 $X2=0
+ $Y2=0
cc_513 N_A_803_297#_c_751_n N_Y_c_822_n 0.00127075f $X=6.535 $Y=2.38 $X2=0 $Y2=0
cc_514 N_A_803_297#_c_800_p N_Y_c_822_n 0.0126766f $X=6.66 $Y=1.96 $X2=0 $Y2=0
cc_515 N_A_803_297#_c_743_n N_Y_c_822_n 0.00320918f $X=7.375 $Y=2.38 $X2=0 $Y2=0
cc_516 N_A_803_297#_c_742_n N_Y_c_923_n 0.00251363f $X=5.82 $Y=1.62 $X2=0 $Y2=0
cc_517 N_A_803_297#_c_751_n N_Y_c_923_n 0.00214463f $X=6.535 $Y=2.38 $X2=0 $Y2=0
cc_518 N_A_803_297#_c_743_n N_Y_c_823_n 0.0118729f $X=7.375 $Y=2.38 $X2=0 $Y2=0
cc_519 N_A_803_297#_c_751_n Y 0.0118865f $X=6.535 $Y=2.38 $X2=0 $Y2=0
cc_520 N_Y_c_806_n N_VGND_M1018_d 0.00162089f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_521 N_Y_c_808_n N_VGND_M1033_d 0.00162089f $X=2.195 $Y=0.815 $X2=0 $Y2=0
cc_522 N_Y_c_809_n N_VGND_M1024_s 0.00162089f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_523 N_Y_c_810_n N_VGND_M1029_s 0.0108248f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_524 N_Y_c_811_n N_VGND_M1016_s 0.00162089f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_525 N_Y_c_812_n N_VGND_M1025_s 0.00162089f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_526 N_Y_c_814_n N_VGND_M1013_s 0.00162089f $X=6.915 $Y=0.815 $X2=0 $Y2=0
cc_527 N_Y_c_807_n N_VGND_c_1008_n 0.00750114f $X=0.845 $Y=0.815 $X2=0 $Y2=0
cc_528 N_Y_c_806_n N_VGND_c_1009_n 0.0122559f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_529 N_Y_c_808_n N_VGND_c_1010_n 0.0122559f $X=2.195 $Y=0.815 $X2=0 $Y2=0
cc_530 N_Y_c_809_n N_VGND_c_1011_n 0.0122559f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_531 N_Y_c_811_n N_VGND_c_1012_n 0.0122559f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_532 N_Y_c_811_n N_VGND_c_1013_n 0.00198695f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_533 N_Y_c_877_n N_VGND_c_1013_n 0.0188551f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_534 N_Y_c_812_n N_VGND_c_1013_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_535 N_Y_c_812_n N_VGND_c_1014_n 0.0122559f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_536 N_Y_c_814_n N_VGND_c_1015_n 0.0122559f $X=6.915 $Y=0.815 $X2=0 $Y2=0
cc_537 N_Y_c_824_n N_VGND_c_1019_n 0.0188551f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_538 N_Y_c_806_n N_VGND_c_1019_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_539 N_Y_c_806_n N_VGND_c_1021_n 0.00198695f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_540 N_Y_c_835_n N_VGND_c_1021_n 0.0188551f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_541 N_Y_c_808_n N_VGND_c_1021_n 0.00198695f $X=2.195 $Y=0.815 $X2=0 $Y2=0
cc_542 N_Y_c_808_n N_VGND_c_1023_n 0.00198695f $X=2.195 $Y=0.815 $X2=0 $Y2=0
cc_543 N_Y_c_840_n N_VGND_c_1023_n 0.0188551f $X=2.36 $Y=0.39 $X2=0 $Y2=0
cc_544 N_Y_c_809_n N_VGND_c_1023_n 0.00198695f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_545 N_Y_c_810_n N_VGND_c_1025_n 0.00198695f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_546 N_Y_c_870_n N_VGND_c_1025_n 0.0188551f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_547 N_Y_c_811_n N_VGND_c_1025_n 0.00198695f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_548 N_Y_c_812_n N_VGND_c_1027_n 0.00198695f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_549 N_Y_c_882_n N_VGND_c_1027_n 0.0188977f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_550 N_Y_c_814_n N_VGND_c_1027_n 0.00118063f $X=6.915 $Y=0.815 $X2=0 $Y2=0
cc_551 N_Y_c_820_n N_VGND_c_1027_n 8.85324e-19 $X=6.27 $Y=0.815 $X2=0 $Y2=0
cc_552 N_Y_c_814_n N_VGND_c_1029_n 0.00198695f $X=6.915 $Y=0.815 $X2=0 $Y2=0
cc_553 N_Y_c_917_n N_VGND_c_1029_n 0.0188551f $X=7.08 $Y=0.39 $X2=0 $Y2=0
cc_554 N_Y_c_809_n N_VGND_c_1032_n 0.00198695f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_555 N_Y_c_855_n N_VGND_c_1032_n 0.0188551f $X=3.2 $Y=0.39 $X2=0 $Y2=0
cc_556 N_Y_c_810_n N_VGND_c_1032_n 0.00198695f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_557 N_Y_c_810_n N_VGND_c_1033_n 0.0528344f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_558 N_Y_M1015_s N_VGND_c_1035_n 0.00215201f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_559 N_Y_M1022_s N_VGND_c_1035_n 0.00215201f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_560 N_Y_M1019_d N_VGND_c_1035_n 0.00215201f $X=2.225 $Y=0.235 $X2=0 $Y2=0
cc_561 N_Y_M1028_d N_VGND_c_1035_n 0.00215201f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_562 N_Y_M1012_d N_VGND_c_1035_n 0.00215201f $X=4.425 $Y=0.235 $X2=0 $Y2=0
cc_563 N_Y_M1020_d N_VGND_c_1035_n 0.00215201f $X=5.265 $Y=0.235 $X2=0 $Y2=0
cc_564 N_Y_M1008_d N_VGND_c_1035_n 0.00215201f $X=6.105 $Y=0.235 $X2=0 $Y2=0
cc_565 N_Y_M1017_d N_VGND_c_1035_n 0.00215201f $X=6.945 $Y=0.235 $X2=0 $Y2=0
cc_566 N_Y_c_824_n N_VGND_c_1035_n 0.0122069f $X=0.68 $Y=0.39 $X2=0 $Y2=0
cc_567 N_Y_c_806_n N_VGND_c_1035_n 0.00835832f $X=1.355 $Y=0.815 $X2=0 $Y2=0
cc_568 N_Y_c_835_n N_VGND_c_1035_n 0.0122069f $X=1.52 $Y=0.39 $X2=0 $Y2=0
cc_569 N_Y_c_808_n N_VGND_c_1035_n 0.00835832f $X=2.195 $Y=0.815 $X2=0 $Y2=0
cc_570 N_Y_c_840_n N_VGND_c_1035_n 0.0122069f $X=2.36 $Y=0.39 $X2=0 $Y2=0
cc_571 N_Y_c_809_n N_VGND_c_1035_n 0.00835832f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_572 N_Y_c_855_n N_VGND_c_1035_n 0.0122069f $X=3.2 $Y=0.39 $X2=0 $Y2=0
cc_573 N_Y_c_810_n N_VGND_c_1035_n 0.0103256f $X=4.395 $Y=0.815 $X2=0 $Y2=0
cc_574 N_Y_c_870_n N_VGND_c_1035_n 0.0122069f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_575 N_Y_c_811_n N_VGND_c_1035_n 0.00835832f $X=5.235 $Y=0.815 $X2=0 $Y2=0
cc_576 N_Y_c_877_n N_VGND_c_1035_n 0.0122069f $X=5.4 $Y=0.39 $X2=0 $Y2=0
cc_577 N_Y_c_812_n N_VGND_c_1035_n 0.00835832f $X=6.075 $Y=0.815 $X2=0 $Y2=0
cc_578 N_Y_c_882_n N_VGND_c_1035_n 0.01222f $X=6.24 $Y=0.39 $X2=0 $Y2=0
cc_579 N_Y_c_814_n N_VGND_c_1035_n 0.00706837f $X=6.915 $Y=0.815 $X2=0 $Y2=0
cc_580 N_Y_c_917_n N_VGND_c_1035_n 0.0122069f $X=7.08 $Y=0.39 $X2=0 $Y2=0
cc_581 N_Y_c_820_n N_VGND_c_1035_n 0.00138075f $X=6.27 $Y=0.815 $X2=0 $Y2=0

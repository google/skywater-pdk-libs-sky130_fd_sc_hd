* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 Y a_105_352# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.05e+11p pd=2.61e+06u as=6.365e+11p ps=5.36e+06u
M1001 a_388_297# A2 Y VPB phighvt w=1e+06u l=150000u
+  ad=2.55e+11p pd=2.51e+06u as=0p ps=0u
M1002 a_297_47# a_105_352# Y VNB nshort w=650000u l=150000u
+  ad=3.705e+11p pd=3.74e+06u as=1.69e+11p ps=1.82e+06u
M1003 VPWR A1 a_388_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_297_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.847e+11p ps=3.2e+06u
M1005 VPWR B1_N a_105_352# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1006 VGND A2 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_105_352# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__inv_16.spice.pex
* Created: Thu Aug 27 14:22:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_16%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34 36
+ 38 41 43 45 48 50 52 55 57 59 62 64 66 69 71 73 76 78 80 83 85 87 90 92 94 97
+ 99 101 104 106 108 111 113 114 115 116 117 118 143 147
r313 146 147 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.415 $Y=1.16
+ $X2=6.835 $Y2=1.16
r314 145 146 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.995 $Y=1.16
+ $X2=6.415 $Y2=1.16
r315 144 145 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.575 $Y=1.16
+ $X2=5.995 $Y2=1.16
r316 142 144 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.36 $Y=1.16
+ $X2=5.575 $Y2=1.16
r317 142 143 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=5.36
+ $Y=1.16 $X2=5.36 $Y2=1.16
r318 140 142 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.155 $Y=1.16
+ $X2=5.36 $Y2=1.16
r319 139 140 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.735 $Y=1.16
+ $X2=5.155 $Y2=1.16
r320 138 139 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.315 $Y=1.16
+ $X2=4.735 $Y2=1.16
r321 137 138 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.895 $Y=1.16
+ $X2=4.315 $Y2=1.16
r322 136 137 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.475 $Y=1.16
+ $X2=3.895 $Y2=1.16
r323 135 136 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.055 $Y=1.16
+ $X2=3.475 $Y2=1.16
r324 134 135 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.635 $Y=1.16
+ $X2=3.055 $Y2=1.16
r325 133 134 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.215 $Y=1.16
+ $X2=2.635 $Y2=1.16
r326 132 133 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.795 $Y=1.16
+ $X2=2.215 $Y2=1.16
r327 131 132 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.375 $Y=1.16
+ $X2=1.795 $Y2=1.16
r328 130 131 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.955 $Y=1.16
+ $X2=1.375 $Y2=1.16
r329 129 130 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.535 $Y=1.16
+ $X2=0.955 $Y2=1.16
r330 126 129 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.295 $Y=1.16
+ $X2=0.535 $Y2=1.16
r331 118 143 47.5383 $w=2.38e-07 $l=9.9e-07 $layer=LI1_cond $X=4.37 $Y=1.195
+ $X2=5.36 $Y2=1.195
r332 117 118 22.0885 $w=2.38e-07 $l=4.6e-07 $layer=LI1_cond $X=3.91 $Y=1.195
+ $X2=4.37 $Y2=1.195
r333 116 117 44.177 $w=2.38e-07 $l=9.2e-07 $layer=LI1_cond $X=2.99 $Y=1.195
+ $X2=3.91 $Y2=1.195
r334 115 116 44.177 $w=2.38e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=1.195
+ $X2=2.99 $Y2=1.195
r335 114 115 44.177 $w=2.38e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=1.195
+ $X2=2.07 $Y2=1.195
r336 113 114 44.177 $w=2.38e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=1.195
+ $X2=1.15 $Y2=1.195
r337 113 126 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=0.295
+ $Y=1.16 $X2=0.295 $Y2=1.16
r338 109 147 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=1.325
+ $X2=6.835 $Y2=1.16
r339 109 111 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.835 $Y=1.325
+ $X2=6.835 $Y2=1.985
r340 106 147 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.835 $Y=0.995
+ $X2=6.835 $Y2=1.16
r341 106 108 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.835 $Y=0.995
+ $X2=6.835 $Y2=0.56
r342 102 146 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.325
+ $X2=6.415 $Y2=1.16
r343 102 104 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.415 $Y=1.325
+ $X2=6.415 $Y2=1.985
r344 99 146 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=0.995
+ $X2=6.415 $Y2=1.16
r345 99 101 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.415 $Y=0.995
+ $X2=6.415 $Y2=0.56
r346 95 145 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.16
r347 95 97 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.995 $Y=1.325
+ $X2=5.995 $Y2=1.985
r348 92 145 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=1.16
r349 92 94 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.995 $Y=0.995
+ $X2=5.995 $Y2=0.56
r350 88 144 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.325
+ $X2=5.575 $Y2=1.16
r351 88 90 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.575 $Y=1.325
+ $X2=5.575 $Y2=1.985
r352 85 144 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=0.995
+ $X2=5.575 $Y2=1.16
r353 85 87 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.575 $Y=0.995
+ $X2=5.575 $Y2=0.56
r354 81 140 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.325
+ $X2=5.155 $Y2=1.16
r355 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.155 $Y=1.325
+ $X2=5.155 $Y2=1.985
r356 78 140 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=0.995
+ $X2=5.155 $Y2=1.16
r357 78 80 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.155 $Y=0.995
+ $X2=5.155 $Y2=0.56
r358 74 139 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.325
+ $X2=4.735 $Y2=1.16
r359 74 76 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.735 $Y=1.325
+ $X2=4.735 $Y2=1.985
r360 71 139 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=0.995
+ $X2=4.735 $Y2=1.16
r361 71 73 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.735 $Y=0.995
+ $X2=4.735 $Y2=0.56
r362 67 138 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.325
+ $X2=4.315 $Y2=1.16
r363 67 69 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.315 $Y=1.325
+ $X2=4.315 $Y2=1.985
r364 64 138 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=1.16
r365 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.315 $Y=0.995
+ $X2=4.315 $Y2=0.56
r366 60 137 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.325
+ $X2=3.895 $Y2=1.16
r367 60 62 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.895 $Y=1.325
+ $X2=3.895 $Y2=1.985
r368 57 137 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=0.995
+ $X2=3.895 $Y2=1.16
r369 57 59 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.895 $Y=0.995
+ $X2=3.895 $Y2=0.56
r370 53 136 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.475 $Y=1.325
+ $X2=3.475 $Y2=1.16
r371 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.475 $Y=1.325
+ $X2=3.475 $Y2=1.985
r372 50 136 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.475 $Y=0.995
+ $X2=3.475 $Y2=1.16
r373 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.475 $Y=0.995
+ $X2=3.475 $Y2=0.56
r374 46 135 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.16
r375 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.325
+ $X2=3.055 $Y2=1.985
r376 43 135 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=0.995
+ $X2=3.055 $Y2=1.16
r377 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.055 $Y=0.995
+ $X2=3.055 $Y2=0.56
r378 39 134 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=1.16
r379 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=1.985
r380 36 134 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=0.995
+ $X2=2.635 $Y2=1.16
r381 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.635 $Y=0.995
+ $X2=2.635 $Y2=0.56
r382 32 133 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.325
+ $X2=2.215 $Y2=1.16
r383 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=1.325
+ $X2=2.215 $Y2=1.985
r384 29 133 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.215 $Y2=1.16
r385 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.215 $Y=0.995
+ $X2=2.215 $Y2=0.56
r386 25 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=1.16
r387 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.795 $Y=1.325
+ $X2=1.795 $Y2=1.985
r388 22 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=0.995
+ $X2=1.795 $Y2=1.16
r389 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.795 $Y=0.995
+ $X2=1.795 $Y2=0.56
r390 18 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.16
r391 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.985
r392 15 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=1.16
r393 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=0.56
r394 11 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r395 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r396 8 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.16
r397 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r398 4 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.325
+ $X2=0.535 $Y2=1.16
r399 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.535 $Y=1.325
+ $X2=0.535 $Y2=1.985
r400 1 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=1.16
r401 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.535 $Y=0.995
+ $X2=0.535 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_16%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 56 60 64 66 68 71 72 74 75 77 78 79 80 82 83 84 103 111 114 118
r116 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r117 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r119 106 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 103 117 3.63957 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=7.16 $Y2=2.72
r122 103 105 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=6.67 $Y2=2.72
r123 102 106 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r124 102 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r125 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r126 99 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=2.72
+ $X2=5.365 $Y2=2.72
r127 99 101 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.45 $Y=2.72
+ $X2=5.75 $Y2=2.72
r128 98 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r130 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r132 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r135 89 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r136 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 86 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.165 $Y2=2.72
r138 86 88 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=2.72
+ $X2=1.61 $Y2=2.72
r139 84 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 84 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r141 82 101 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.12 $Y=2.72
+ $X2=5.75 $Y2=2.72
r142 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=2.72
+ $X2=6.205 $Y2=2.72
r143 81 105 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.29 $Y=2.72
+ $X2=6.67 $Y2=2.72
r144 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.29 $Y=2.72
+ $X2=6.205 $Y2=2.72
r145 79 97 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.44 $Y=2.72 $X2=4.37
+ $Y2=2.72
r146 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=2.72
+ $X2=4.525 $Y2=2.72
r147 77 94 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=2.72 $X2=3.45
+ $Y2=2.72
r148 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.72
+ $X2=3.685 $Y2=2.72
r149 76 97 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.77 $Y=2.72 $X2=4.37
+ $Y2=2.72
r150 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.72
+ $X2=3.685 $Y2=2.72
r151 74 91 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.76 $Y=2.72
+ $X2=2.53 $Y2=2.72
r152 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=2.72
+ $X2=2.845 $Y2=2.72
r153 73 94 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=3.45 $Y2=2.72
r154 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=2.845 $Y2=2.72
r155 71 88 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=1.61 $Y2=2.72
r156 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.72
+ $X2=2.005 $Y2=2.72
r157 70 91 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=2.72
+ $X2=2.53 $Y2=2.72
r158 70 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=2.72
+ $X2=2.005 $Y2=2.72
r159 66 117 3.27562 $w=2.1e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.16 $Y2=2.72
r160 66 68 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=7.065 $Y=2.635
+ $X2=7.065 $Y2=2
r161 62 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=2.635
+ $X2=6.205 $Y2=2.72
r162 62 64 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.205 $Y=2.635
+ $X2=6.205 $Y2=2
r163 58 114 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=2.635
+ $X2=5.365 $Y2=2.72
r164 58 60 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.365 $Y=2.635
+ $X2=5.365 $Y2=2
r165 57 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=2.72
+ $X2=4.525 $Y2=2.72
r166 56 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=2.72
+ $X2=5.365 $Y2=2.72
r167 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.28 $Y=2.72
+ $X2=4.61 $Y2=2.72
r168 52 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=2.635
+ $X2=4.525 $Y2=2.72
r169 52 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.525 $Y=2.635
+ $X2=4.525 $Y2=2
r170 48 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.635
+ $X2=3.685 $Y2=2.72
r171 48 50 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.685 $Y=2.635
+ $X2=3.685 $Y2=2
r172 44 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=2.635
+ $X2=2.845 $Y2=2.72
r173 44 46 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.845 $Y=2.635
+ $X2=2.845 $Y2=2
r174 40 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=2.635
+ $X2=2.005 $Y2=2.72
r175 40 42 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.005 $Y=2.635
+ $X2=2.005 $Y2=2
r176 36 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.635
+ $X2=1.165 $Y2=2.72
r177 36 38 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.165 $Y=2.635
+ $X2=1.165 $Y2=2
r178 35 108 3.63491 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=0.205 $Y2=2.72
r179 34 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2.72
+ $X2=1.165 $Y2=2.72
r180 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.08 $Y=2.72
+ $X2=0.41 $Y2=2.72
r181 30 33 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=0.305 $Y=1.65
+ $X2=0.305 $Y2=2.34
r182 28 108 3.28028 $w=2.1e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.205 $Y2=2.72
r183 28 33 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.305 $Y2=2.34
r184 9 68 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.91
+ $Y=1.485 $X2=7.045 $Y2=2
r185 8 64 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=6.07
+ $Y=1.485 $X2=6.205 $Y2=2
r186 7 60 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=5.23
+ $Y=1.485 $X2=5.365 $Y2=2
r187 6 54 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.39
+ $Y=1.485 $X2=4.525 $Y2=2
r188 5 50 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.55
+ $Y=1.485 $X2=3.685 $Y2=2
r189 4 46 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.71
+ $Y=1.485 $X2=2.845 $Y2=2
r190 3 42 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.87
+ $Y=1.485 $X2=2.005 $Y2=2
r191 2 38 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=2
r192 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.485 $X2=0.325 $Y2=2.34
r193 1 30 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.485 $X2=0.325 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__INV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 53 55 57 58 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 105 107 111 115 117
+ 119 123 127 129 131 135 139 143 145 146 148 149 151 152 154 155 157 158 160
+ 163 164 165
r288 164 169 3.19459 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=6.625 $Y=0.81
+ $X2=6.625 $Y2=0.905
r289 164 165 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.625 $Y=0.92
+ $X2=6.625 $Y2=1.19
r290 164 169 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=6.625 $Y=0.92
+ $X2=6.625 $Y2=0.905
r291 161 165 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.625 $Y=1.495
+ $X2=6.625 $Y2=1.19
r292 161 163 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.625 $Y=1.495
+ $X2=6.625 $Y2=1.58
r293 137 163 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.625 $Y=1.665
+ $X2=6.625 $Y2=1.58
r294 137 139 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.625 $Y=1.665
+ $X2=6.625 $Y2=2.34
r295 133 164 3.19459 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=6.625 $Y=0.715
+ $X2=6.625 $Y2=0.81
r296 133 135 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.625 $Y=0.715
+ $X2=6.625 $Y2=0.38
r297 132 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=1.58
+ $X2=5.785 $Y2=1.58
r298 131 163 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=1.58
+ $X2=6.625 $Y2=1.58
r299 131 132 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.46 $Y=1.58
+ $X2=5.95 $Y2=1.58
r300 130 158 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=0.81
+ $X2=5.785 $Y2=0.81
r301 129 164 3.38787 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=0.81
+ $X2=6.625 $Y2=0.81
r302 129 130 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=6.46 $Y=0.81
+ $X2=5.95 $Y2=0.81
r303 125 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=1.665
+ $X2=5.785 $Y2=1.58
r304 125 127 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.785 $Y=1.665
+ $X2=5.785 $Y2=2.34
r305 121 158 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.785 $Y=0.715
+ $X2=5.785 $Y2=0.81
r306 121 123 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.785 $Y=0.715
+ $X2=5.785 $Y2=0.38
r307 120 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=1.58
+ $X2=4.945 $Y2=1.58
r308 119 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=1.58
+ $X2=5.785 $Y2=1.58
r309 119 120 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.62 $Y=1.58
+ $X2=5.11 $Y2=1.58
r310 118 155 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.11 $Y=0.81
+ $X2=4.945 $Y2=0.81
r311 117 158 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0.81
+ $X2=5.785 $Y2=0.81
r312 117 118 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=5.62 $Y=0.81
+ $X2=5.11 $Y2=0.81
r313 113 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=1.665
+ $X2=4.945 $Y2=1.58
r314 113 115 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.945 $Y=1.665
+ $X2=4.945 $Y2=2.34
r315 109 155 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.945 $Y=0.715
+ $X2=4.945 $Y2=0.81
r316 109 111 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.945 $Y=0.715
+ $X2=4.945 $Y2=0.38
r317 108 154 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=1.58
+ $X2=4.105 $Y2=1.58
r318 107 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=1.58
+ $X2=4.945 $Y2=1.58
r319 107 108 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.78 $Y=1.58
+ $X2=4.27 $Y2=1.58
r320 106 152 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0.81
+ $X2=4.105 $Y2=0.81
r321 105 155 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.78 $Y=0.81
+ $X2=4.945 $Y2=0.81
r322 105 106 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=4.78 $Y=0.81
+ $X2=4.27 $Y2=0.81
r323 101 154 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=1.665
+ $X2=4.105 $Y2=1.58
r324 101 103 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.105 $Y=1.665
+ $X2=4.105 $Y2=2.34
r325 97 152 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.105 $Y=0.715
+ $X2=4.105 $Y2=0.81
r326 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=0.715
+ $X2=4.105 $Y2=0.38
r327 96 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=1.58
+ $X2=3.265 $Y2=1.58
r328 95 154 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.94 $Y=1.58
+ $X2=4.105 $Y2=1.58
r329 95 96 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.94 $Y=1.58
+ $X2=3.43 $Y2=1.58
r330 94 149 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=0.81
+ $X2=3.265 $Y2=0.81
r331 93 152 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.94 $Y=0.81
+ $X2=4.105 $Y2=0.81
r332 93 94 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.94 $Y=0.81
+ $X2=3.43 $Y2=0.81
r333 89 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=1.665
+ $X2=3.265 $Y2=1.58
r334 89 91 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.265 $Y=1.665
+ $X2=3.265 $Y2=2.34
r335 85 149 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.265 $Y=0.715
+ $X2=3.265 $Y2=0.81
r336 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=0.715
+ $X2=3.265 $Y2=0.38
r337 84 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=1.58
+ $X2=2.425 $Y2=1.58
r338 83 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=1.58
+ $X2=3.265 $Y2=1.58
r339 83 84 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.1 $Y=1.58
+ $X2=2.59 $Y2=1.58
r340 82 146 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0.81
+ $X2=2.425 $Y2=0.81
r341 81 149 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=0.81
+ $X2=3.265 $Y2=0.81
r342 81 82 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=3.1 $Y=0.81
+ $X2=2.59 $Y2=0.81
r343 77 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=1.665
+ $X2=2.425 $Y2=1.58
r344 77 79 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.425 $Y=1.665
+ $X2=2.425 $Y2=2.34
r345 73 146 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.425 $Y=0.715
+ $X2=2.425 $Y2=0.81
r346 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.425 $Y=0.715
+ $X2=2.425 $Y2=0.38
r347 72 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=1.58
+ $X2=1.585 $Y2=1.58
r348 71 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=1.58
+ $X2=2.425 $Y2=1.58
r349 71 72 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.26 $Y=1.58
+ $X2=1.75 $Y2=1.58
r350 70 143 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=0.81
+ $X2=1.585 $Y2=0.81
r351 69 146 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0.81
+ $X2=2.425 $Y2=0.81
r352 69 70 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.26 $Y=0.81
+ $X2=1.75 $Y2=0.81
r353 65 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.665
+ $X2=1.585 $Y2=1.58
r354 65 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.585 $Y=1.665
+ $X2=1.585 $Y2=2.34
r355 61 143 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.585 $Y=0.715
+ $X2=1.585 $Y2=0.81
r356 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.585 $Y=0.715
+ $X2=1.585 $Y2=0.38
r357 60 142 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=1.58
+ $X2=0.745 $Y2=1.58
r358 59 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=1.58
+ $X2=1.585 $Y2=1.58
r359 59 60 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.42 $Y=1.58
+ $X2=0.91 $Y2=1.58
r360 57 143 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=0.81
+ $X2=1.585 $Y2=0.81
r361 57 58 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=1.42 $Y=0.81
+ $X2=0.91 $Y2=0.81
r362 53 142 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=1.58
r363 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=2.34
r364 49 58 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.745 $Y=0.715
+ $X2=0.91 $Y2=0.81
r365 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.745 $Y=0.715
+ $X2=0.745 $Y2=0.38
r366 16 163 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.485 $X2=6.625 $Y2=1.65
r367 16 139 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.49
+ $Y=1.485 $X2=6.625 $Y2=2.34
r368 15 160 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=5.65
+ $Y=1.485 $X2=5.785 $Y2=1.65
r369 15 127 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.65
+ $Y=1.485 $X2=5.785 $Y2=2.34
r370 14 157 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.485 $X2=4.945 $Y2=1.65
r371 14 115 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.485 $X2=4.945 $Y2=2.34
r372 13 154 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.485 $X2=4.105 $Y2=1.65
r373 13 103 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.485 $X2=4.105 $Y2=2.34
r374 12 151 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.485 $X2=3.265 $Y2=1.65
r375 12 91 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.485 $X2=3.265 $Y2=2.34
r376 11 148 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.425 $Y2=1.65
r377 11 79 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.485 $X2=2.425 $Y2=2.34
r378 10 145 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.585 $Y2=1.65
r379 10 67 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.585 $Y2=2.34
r380 9 142 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.485 $X2=0.745 $Y2=1.65
r381 9 55 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.485 $X2=0.745 $Y2=2.34
r382 8 135 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.49
+ $Y=0.235 $X2=6.625 $Y2=0.38
r383 7 123 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.65
+ $Y=0.235 $X2=5.785 $Y2=0.38
r384 6 111 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.235 $X2=4.945 $Y2=0.38
r385 5 99 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.97
+ $Y=0.235 $X2=4.105 $Y2=0.38
r386 4 87 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.235 $X2=3.265 $Y2=0.38
r387 3 75 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.235 $X2=2.425 $Y2=0.38
r388 2 63 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.45
+ $Y=0.235 $X2=1.585 $Y2=0.38
r389 1 51 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.235 $X2=0.745 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__INV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 32 36 40 44 48
+ 52 54 58 62 64 66 69 70 72 73 75 76 77 78 80 81 82 101 109 112 116
r136 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r137 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r138 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r139 104 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r140 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r141 101 115 3.63957 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.16
+ $Y2=0
r142 101 103 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=6.67 $Y2=0
r143 100 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r144 100 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r145 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r146 97 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=0 $X2=5.365
+ $Y2=0
r147 97 99 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.45 $Y=0 $X2=5.75
+ $Y2=0
r148 96 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r149 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r150 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r151 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r152 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r153 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r154 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r155 87 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r156 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r157 84 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.165
+ $Y2=0
r158 84 86 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.61
+ $Y2=0
r159 82 110 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r160 82 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r161 80 99 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.12 $Y=0 $X2=5.75
+ $Y2=0
r162 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=0 $X2=6.205
+ $Y2=0
r163 79 103 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.29 $Y=0 $X2=6.67
+ $Y2=0
r164 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.29 $Y=0 $X2=6.205
+ $Y2=0
r165 77 95 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.37
+ $Y2=0
r166 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.525
+ $Y2=0
r167 75 92 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.45
+ $Y2=0
r168 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0 $X2=3.685
+ $Y2=0
r169 74 95 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.77 $Y=0 $X2=4.37
+ $Y2=0
r170 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=0 $X2=3.685
+ $Y2=0
r171 72 89 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.53
+ $Y2=0
r172 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.845
+ $Y2=0
r173 71 92 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=3.45
+ $Y2=0
r174 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0 $X2=2.845
+ $Y2=0
r175 69 86 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.61
+ $Y2=0
r176 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.005
+ $Y2=0
r177 68 89 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.53
+ $Y2=0
r178 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.005
+ $Y2=0
r179 64 115 3.27562 $w=2.1e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.065 $Y=0.085
+ $X2=7.16 $Y2=0
r180 64 66 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=7.065 $Y=0.085
+ $X2=7.065 $Y2=0.38
r181 60 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=0.085
+ $X2=6.205 $Y2=0
r182 60 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.205 $Y=0.085
+ $X2=6.205 $Y2=0.38
r183 56 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0
r184 56 58 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0.38
r185 55 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=0 $X2=4.525
+ $Y2=0
r186 54 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=0 $X2=5.365
+ $Y2=0
r187 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.28 $Y=0 $X2=4.61
+ $Y2=0
r188 50 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0
r189 50 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0.38
r190 46 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r191 46 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.38
r192 42 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0
r193 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.845 $Y=0.085
+ $X2=2.845 $Y2=0.38
r194 38 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0
r195 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.005 $Y=0.085
+ $X2=2.005 $Y2=0.38
r196 34 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0
r197 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.165 $Y=0.085
+ $X2=1.165 $Y2=0.38
r198 33 106 3.78596 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=0
+ $X2=0.205 $Y2=0
r199 32 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=0 $X2=1.165
+ $Y2=0
r200 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.41
+ $Y2=0
r201 28 106 3.23192 $w=2.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.205 $Y2=0
r202 28 30 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.38
r203 9 66 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.91
+ $Y=0.235 $X2=7.045 $Y2=0.38
r204 8 62 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.235 $X2=6.205 $Y2=0.38
r205 7 58 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.23
+ $Y=0.235 $X2=5.365 $Y2=0.38
r206 6 52 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.235 $X2=4.525 $Y2=0.38
r207 5 48 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.235 $X2=3.685 $Y2=0.38
r208 4 44 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.845 $Y2=0.38
r209 3 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.235 $X2=2.005 $Y2=0.38
r210 2 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.38
r211 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.2
+ $Y=0.235 $X2=0.325 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o41ai_4.pex.spice
* Created: Tue Sep  1 19:26:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O41AI_4%B1 3 7 11 15 19 23 25 27 31 33 34 35 36
r76 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r77 42 44 34.1782 $w=2.75e-07 $l=1.95e-07 $layer=POLY_cond $X=0.275 $Y=1.16
+ $X2=0.47 $Y2=1.16
r78 36 49 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.52 $Y2=1.175
r79 35 49 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.52 $Y2=1.175
r80 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r81 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r82 33 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r83 25 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.52 $Y2=1.16
r84 25 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.985
r85 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.73 $Y=1.025
+ $X2=1.73 $Y2=0.56
r86 17 48 36.8073 $w=2.75e-07 $l=2.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.52 $Y2=1.16
r87 17 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.31 $Y=1.295
+ $X2=1.31 $Y2=1.985
r88 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.31 $Y=1.025
+ $X2=1.31 $Y2=0.56
r89 9 17 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=1.31 $Y2=1.16
r90 9 44 73.6145 $w=2.75e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.16
+ $X2=0.47 $Y2=1.16
r91 9 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.89 $Y=1.295
+ $X2=0.89 $Y2=1.985
r92 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.89 $Y=1.025
+ $X2=0.89 $Y2=0.56
r93 5 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.305
+ $X2=0.47 $Y2=1.16
r94 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.47 $Y=1.305 $X2=0.47
+ $Y2=1.985
r95 1 44 16.9318 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=1.16
r96 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A4 1 3 6 10 14 18 22 24 26 30 32 33 34 35
r96 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.72
+ $Y=1.16 $X2=3.72 $Y2=1.16
r97 41 43 26.3063 $w=2.84e-07 $l=1.55e-07 $layer=POLY_cond $X=2.515 $Y=1.16
+ $X2=2.67 $Y2=1.16
r98 35 48 11.9227 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=3.935 $Y=1.175
+ $X2=3.72 $Y2=1.175
r99 34 48 13.5864 $w=1.98e-07 $l=2.45e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.72 $Y2=1.175
r100 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.475 $Y2=1.175
r101 32 33 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=2.515 $Y=1.175
+ $X2=3.015 $Y2=1.175
r102 32 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.515
+ $Y=1.16 $X2=2.515 $Y2=1.16
r103 24 47 35.6408 $w=2.84e-07 $l=2.1e-07 $layer=POLY_cond $X=3.93 $Y=1.16
+ $X2=3.72 $Y2=1.16
r104 24 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.985
r105 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.93 $Y=1.025
+ $X2=3.93 $Y2=0.56
r106 16 47 35.6408 $w=2.84e-07 $l=2.1e-07 $layer=POLY_cond $X=3.51 $Y=1.16
+ $X2=3.72 $Y2=1.16
r107 16 22 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.51 $Y=1.295
+ $X2=3.51 $Y2=1.985
r108 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=1.025
+ $X2=3.51 $Y2=0.56
r109 8 16 71.2817 $w=2.84e-07 $l=4.2e-07 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=3.51 $Y2=1.16
r110 8 43 71.2817 $w=2.84e-07 $l=4.2e-07 $layer=POLY_cond $X=3.09 $Y=1.16
+ $X2=2.67 $Y2=1.16
r111 8 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.09 $Y=1.295
+ $X2=3.09 $Y2=1.985
r112 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.09 $Y=1.025
+ $X2=3.09 $Y2=0.56
r113 4 43 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.16
r114 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.325
+ $X2=2.67 $Y2=1.985
r115 1 43 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r116 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 41 43
c93 36 0 1.75804e-19 $X=5.775 $Y=1.19
c94 7 0 6.60366e-20 $X=4.35 $Y=1.985
r95 52 53 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=5.19 $Y=1.16 $X2=5.61
+ $Y2=1.16
r96 51 52 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.16 $X2=5.19
+ $Y2=1.16
r97 49 51 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.77 $Y2=1.16
r98 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.56
+ $Y=1.16 $X2=4.56 $Y2=1.16
r99 46 49 46.6565 $w=2.7e-07 $l=2.1e-07 $layer=POLY_cond $X=4.35 $Y=1.16
+ $X2=4.56 $Y2=1.16
r100 41 53 16.663 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.685 $Y=1.16
+ $X2=5.61 $Y2=1.16
r101 41 43 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=5.685 $Y=1.16
+ $X2=5.815 $Y2=1.16
r102 36 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.815
+ $Y=1.16 $X2=5.815 $Y2=1.16
r103 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=5.315 $Y=1.175
+ $X2=5.775 $Y2=1.175
r104 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=5.315 $Y2=1.175
r105 34 50 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=1.175
+ $X2=4.56 $Y2=1.175
r106 33 50 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.175
+ $X2=4.56 $Y2=1.175
r107 29 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.16
r108 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.295
+ $X2=5.61 $Y2=1.985
r109 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=1.16
r110 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.61 $Y=1.025
+ $X2=5.61 $Y2=0.56
r111 21 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.16
r112 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.19 $Y=1.295
+ $X2=5.19 $Y2=1.985
r113 17 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=1.16
r114 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.19 $Y=1.025
+ $X2=5.19 $Y2=0.56
r115 13 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.16
r116 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=1.295
+ $X2=4.77 $Y2=1.985
r117 9 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=1.16
r118 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.77 $Y=1.025
+ $X2=4.77 $Y2=0.56
r119 5 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.16
r120 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.985
r121 1 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=1.16
r122 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.35 $Y=1.025
+ $X2=4.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 50 51
c100 51 0 1.75804e-19 $X=7.81 $Y=1.16
r101 49 51 7.77608 $w=2.7e-07 $l=3.5e-08 $layer=POLY_cond $X=7.775 $Y=1.16
+ $X2=7.81 $Y2=1.16
r102 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.775
+ $Y=1.16 $X2=7.775 $Y2=1.16
r103 47 49 85.5369 $w=2.7e-07 $l=3.85e-07 $layer=POLY_cond $X=7.39 $Y=1.16
+ $X2=7.775 $Y2=1.16
r104 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.97 $Y=1.16
+ $X2=7.39 $Y2=1.16
r105 45 46 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.55 $Y=1.16
+ $X2=6.97 $Y2=1.16
r106 42 45 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=6.53 $Y=1.16 $X2=6.55
+ $Y2=1.16
r107 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.16 $X2=6.53 $Y2=1.16
r108 36 50 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=7.635 $Y=1.175
+ $X2=7.775 $Y2=1.175
r109 35 36 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=7.175 $Y=1.175
+ $X2=7.635 $Y2=1.175
r110 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.715 $Y=1.175
+ $X2=7.175 $Y2=1.175
r111 34 43 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=6.715 $Y=1.175
+ $X2=6.53 $Y2=1.175
r112 33 43 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=6.255 $Y=1.175
+ $X2=6.53 $Y2=1.175
r113 29 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.16
r114 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.81 $Y=1.295
+ $X2=7.81 $Y2=1.985
r115 25 51 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.81 $Y=1.025
+ $X2=7.81 $Y2=1.16
r116 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.81 $Y=1.025
+ $X2=7.81 $Y2=0.56
r117 21 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.39 $Y=1.295
+ $X2=7.39 $Y2=1.16
r118 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.39 $Y=1.295
+ $X2=7.39 $Y2=1.985
r119 17 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.39 $Y=1.025
+ $X2=7.39 $Y2=1.16
r120 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.39 $Y=1.025
+ $X2=7.39 $Y2=0.56
r121 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.16
r122 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.97 $Y=1.295
+ $X2=6.97 $Y2=1.985
r123 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.97 $Y=1.025
+ $X2=6.97 $Y2=1.16
r124 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.97 $Y=1.025
+ $X2=6.97 $Y2=0.56
r125 5 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.16
r126 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.55 $Y=1.295
+ $X2=6.55 $Y2=1.985
r127 1 45 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=1.16
r128 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.55 $Y=1.025
+ $X2=6.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 50 62
r88 48 50 9.99782 $w=2.7e-07 $l=4.5e-08 $layer=POLY_cond $X=9.49 $Y=1.16
+ $X2=9.535 $Y2=1.16
r89 47 48 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.07 $Y=1.16 $X2=9.49
+ $Y2=1.16
r90 46 47 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=8.65 $Y=1.16 $X2=9.07
+ $Y2=1.16
r91 44 46 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=8.32 $Y=1.16
+ $X2=8.65 $Y2=1.16
r92 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.32
+ $Y=1.16 $X2=8.32 $Y2=1.16
r93 41 44 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=8.23 $Y=1.16 $X2=8.32
+ $Y2=1.16
r94 36 62 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=9.935 $Y=1.175
+ $X2=9.93 $Y2=1.175
r95 35 62 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=9.475 $Y=1.175
+ $X2=9.93 $Y2=1.175
r96 35 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.535
+ $Y=1.16 $X2=9.535 $Y2=1.16
r97 34 35 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=9.015 $Y=1.175
+ $X2=9.475 $Y2=1.175
r98 33 34 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=8.555 $Y=1.175
+ $X2=9.015 $Y2=1.175
r99 33 45 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=8.555 $Y=1.175
+ $X2=8.32 $Y2=1.175
r100 29 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.49 $Y=1.295
+ $X2=9.49 $Y2=1.16
r101 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.49 $Y=1.295
+ $X2=9.49 $Y2=1.985
r102 25 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.49 $Y=1.025
+ $X2=9.49 $Y2=1.16
r103 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.49 $Y=1.025
+ $X2=9.49 $Y2=0.56
r104 21 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.07 $Y=1.295
+ $X2=9.07 $Y2=1.16
r105 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.07 $Y=1.295
+ $X2=9.07 $Y2=1.985
r106 17 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.07 $Y=1.025
+ $X2=9.07 $Y2=1.16
r107 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.07 $Y=1.025
+ $X2=9.07 $Y2=0.56
r108 13 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.65 $Y=1.295
+ $X2=8.65 $Y2=1.16
r109 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.65 $Y=1.295
+ $X2=8.65 $Y2=1.985
r110 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.65 $Y=1.025
+ $X2=8.65 $Y2=1.16
r111 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.65 $Y=1.025
+ $X2=8.65 $Y2=0.56
r112 5 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.23 $Y=1.295
+ $X2=8.23 $Y2=1.16
r113 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.23 $Y=1.295
+ $X2=8.23 $Y2=1.985
r114 1 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.23 $Y=1.025
+ $X2=8.23 $Y2=1.16
r115 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.23 $Y=1.025
+ $X2=8.23 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%VPWR 1 2 3 4 5 16 18 24 28 32 36 39 40 42 43
+ 45 46 47 53 65 66 72
c129 3 0 8.32868e-20 $X=1.805 $Y=1.485
r130 72 73 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r131 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r132 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r133 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r134 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r135 60 73 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 59 60 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r137 57 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=1.98 $Y2=2.72
r138 57 59 387.856 $w=1.68e-07 $l=5.945e-06 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=8.05 $Y2=2.72
r139 56 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r140 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r141 53 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.98 $Y2=2.72
r142 53 55 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r143 52 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r144 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r145 49 69 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r146 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 47 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 47 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r149 45 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.195 $Y=2.72
+ $X2=8.97 $Y2=2.72
r150 45 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.195 $Y=2.72
+ $X2=9.28 $Y2=2.72
r151 44 65 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.365 $Y=2.72
+ $X2=9.89 $Y2=2.72
r152 44 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=2.72
+ $X2=9.28 $Y2=2.72
r153 42 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.05 $Y2=2.72
r154 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=2.72
+ $X2=8.44 $Y2=2.72
r155 41 62 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.525 $Y=2.72
+ $X2=8.97 $Y2=2.72
r156 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=2.72
+ $X2=8.44 $Y2=2.72
r157 39 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r158 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=1.1 $Y2=2.72
r159 38 55 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.61 $Y2=2.72
r160 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=2.72
+ $X2=1.1 $Y2=2.72
r161 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.28 $Y2=2.72
r162 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.28 $Y2=2
r163 30 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=2.635
+ $X2=8.44 $Y2=2.72
r164 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.44 $Y=2.635
+ $X2=8.44 $Y2=2
r165 26 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2.72
r166 26 28 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.98 $Y=2.635
+ $X2=1.98 $Y2=2
r167 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r168 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r169 18 21 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r170 16 69 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r171 16 21 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r172 5 36 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=2
r173 4 32 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=2
r174 3 28 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.485 $X2=1.94 $Y2=2
r175 2 24 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r176 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r177 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%Y 1 2 3 4 5 6 19 27 29 33 35 36 37 38 39 40
+ 41 42 55 59 62 70 77
c98 59 0 8.32868e-20 $X=1.87 $Y=1.53
c99 29 0 6.60366e-20 $X=3.555 $Y=1.53
c100 19 0 7.2785e-20 $X=1.87 $Y=0.77
r101 77 80 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.52 $Y=1.66
+ $X2=1.52 $Y2=2.34
r102 70 73 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.68 $Y=1.66
+ $X2=0.68 $Y2=2.34
r103 42 59 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.015 $Y=1.53
+ $X2=1.87 $Y2=1.53
r104 41 42 8.2563 $w=4.58e-07 $l=2.55e-07 $layer=LI1_cond $X=2.015 $Y=1.19
+ $X2=2.015 $Y2=1.445
r105 40 62 3.29198 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=2.015 $Y=0.77
+ $X2=2.015 $Y2=0.905
r106 40 41 10.7296 $w=2.88e-07 $l=2.7e-07 $layer=LI1_cond $X=2.015 $Y=0.92
+ $X2=2.015 $Y2=1.19
r107 40 62 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.015 $Y=0.92
+ $X2=2.015 $Y2=0.905
r108 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.53
+ $X2=1.355 $Y2=1.53
r109 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.53
+ $X2=1.685 $Y2=1.53
r110 39 77 2.33884 $w=4.83e-07 $l=4.5e-08 $layer=LI1_cond $X=1.52 $Y=1.615
+ $X2=1.52 $Y2=1.66
r111 39 59 11.6128 $w=1.68e-07 $l=1.78e-07 $layer=LI1_cond $X=1.692 $Y=1.53
+ $X2=1.87 $Y2=1.53
r112 39 60 0.456684 $w=1.68e-07 $l=7e-09 $layer=LI1_cond $X=1.692 $Y=1.53
+ $X2=1.685 $Y2=1.53
r113 38 55 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.155 $Y=1.53
+ $X2=1.355 $Y2=1.53
r114 38 56 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.155 $Y=1.53
+ $X2=0.845 $Y2=1.53
r115 37 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.53
+ $X2=0.845 $Y2=1.53
r116 37 70 2.46016 $w=4.98e-07 $l=4.5e-08 $layer=LI1_cond $X=0.68 $Y=1.615
+ $X2=0.68 $Y2=1.66
r117 35 42 20.2515 $w=3.38e-07 $l=5.55e-07 $layer=LI1_cond $X=2.715 $Y=1.53
+ $X2=2.16 $Y2=1.53
r118 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.715 $Y=1.53
+ $X2=2.88 $Y2=1.53
r119 31 33 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.72 $Y=1.615
+ $X2=3.72 $Y2=1.66
r120 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=1.53
+ $X2=2.88 $Y2=1.53
r121 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.72 $Y2=1.615
r122 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.555 $Y=1.53
+ $X2=3.045 $Y2=1.53
r123 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=2.88 $Y2=1.53
r124 25 27 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.88 $Y=1.615
+ $X2=2.88 $Y2=1.66
r125 21 24 35.8538 $w=2.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.68 $Y=0.77
+ $X2=1.52 $Y2=0.77
r126 19 40 3.53583 $w=2.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.87 $Y=0.77
+ $X2=2.015 $Y2=0.77
r127 19 24 14.9391 $w=2.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.87 $Y=0.77
+ $X2=1.52 $Y2=0.77
r128 6 33 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.485 $X2=3.72 $Y2=1.66
r129 5 27 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.485 $X2=2.88 $Y2=1.66
r130 4 80 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=2.34
r131 4 77 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.66
r132 3 73 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=2.34
r133 3 70 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.66
r134 2 24 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.72
r135 1 21 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A_467_297# 1 2 3 4 5 18 20 21 24 26 28 32 36
+ 38 42 44 47
c71 32 0 1.18248e-19 $X=4.815 $Y=1.53
r72 40 42 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.82 $Y=1.615
+ $X2=5.82 $Y2=1.66
r73 39 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=1.53
+ $X2=4.98 $Y2=1.53
r74 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.655 $Y=1.53
+ $X2=5.82 $Y2=1.615
r75 38 39 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.655 $Y=1.53
+ $X2=5.145 $Y2=1.53
r76 34 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.615
+ $X2=4.98 $Y2=1.53
r77 34 36 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.98 $Y=1.615
+ $X2=4.98 $Y2=1.66
r78 33 46 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=1.53
+ $X2=4.14 $Y2=1.53
r79 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=1.53
+ $X2=4.98 $Y2=1.53
r80 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.815 $Y=1.53
+ $X2=4.225 $Y2=1.53
r81 29 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.14 $Y=2.295
+ $X2=4.14 $Y2=2.29
r82 28 46 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=1.615
+ $X2=4.14 $Y2=1.53
r83 28 31 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.14 $Y=1.615
+ $X2=4.14 $Y2=2.29
r84 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2.38 $X2=3.3
+ $Y2=2.38
r85 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=2.38
+ $X2=4.14 $Y2=2.295
r86 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.055 $Y=2.38
+ $X2=3.385 $Y2=2.38
r87 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.295 $X2=3.3
+ $Y2=2.38
r88 22 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.3 $Y=2.295 $X2=3.3
+ $Y2=1.95
r89 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.38 $X2=3.3
+ $Y2=2.38
r90 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.215 $Y=2.38
+ $X2=2.545 $Y2=2.38
r91 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.42 $Y=2.295
+ $X2=2.545 $Y2=2.38
r92 16 18 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.42 $Y=2.295
+ $X2=2.42 $Y2=1.95
r93 5 42 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.485 $X2=5.82 $Y2=1.66
r94 4 36 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.485 $X2=4.98 $Y2=1.66
r95 3 46 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=1.61
r96 3 31 400 $w=1.7e-07 $l=8.69885e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.14 $Y2=2.29
r97 2 24 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.485 $X2=3.3 $Y2=1.95
r98 1 18 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.485 $X2=2.46 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A_885_297# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r41 31 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.6 $Y=2.295 $X2=7.6
+ $Y2=1.95
r42 30 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=2.38
+ $X2=6.76 $Y2=2.38
r43 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.515 $Y=2.38
+ $X2=7.6 $Y2=2.295
r44 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.515 $Y=2.38
+ $X2=6.845 $Y2=2.38
r45 25 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=2.295
+ $X2=6.76 $Y2=2.38
r46 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.76 $Y=2.295
+ $X2=6.76 $Y2=1.95
r47 24 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=2.38 $X2=5.4
+ $Y2=2.38
r48 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=2.38
+ $X2=6.76 $Y2=2.38
r49 23 24 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=6.675 $Y=2.38
+ $X2=5.485 $Y2=2.38
r50 19 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=2.295 $X2=5.4
+ $Y2=2.38
r51 19 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.4 $Y=2.295 $X2=5.4
+ $Y2=1.95
r52 17 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=2.38 $X2=5.4
+ $Y2=2.38
r53 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.315 $Y=2.38
+ $X2=4.645 $Y2=2.38
r54 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.52 $Y=2.295
+ $X2=4.645 $Y2=2.38
r55 13 15 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.52 $Y=2.295
+ $X2=4.52 $Y2=1.95
r56 4 33 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=1.95
r57 3 27 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=1.95
r58 2 21 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.265
+ $Y=1.485 $X2=5.4 $Y2=1.95
r59 1 15 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.425
+ $Y=1.485 $X2=4.56 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A_1243_297# 1 2 3 4 5 18 20 21 24 26 30 34
+ 38 42 46 50 51 52
r85 46 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.7 $Y=1.66 $X2=9.7
+ $Y2=2.34
r86 44 46 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.7 $Y=1.615 $X2=9.7
+ $Y2=1.66
r87 43 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=1.53
+ $X2=8.86 $Y2=1.53
r88 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.535 $Y=1.53
+ $X2=9.7 $Y2=1.615
r89 42 43 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.535 $Y=1.53
+ $X2=9.025 $Y2=1.53
r90 38 40 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.86 $Y=1.66
+ $X2=8.86 $Y2=2.34
r91 36 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=1.615
+ $X2=8.86 $Y2=1.53
r92 36 38 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.86 $Y=1.615
+ $X2=8.86 $Y2=1.66
r93 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=1.53
+ $X2=8.02 $Y2=1.53
r94 34 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=1.53
+ $X2=8.86 $Y2=1.53
r95 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.695 $Y=1.53
+ $X2=8.185 $Y2=1.53
r96 30 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.02 $Y=1.66
+ $X2=8.02 $Y2=2.34
r97 28 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=1.615
+ $X2=8.02 $Y2=1.53
r98 28 30 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.02 $Y=1.615
+ $X2=8.02 $Y2=1.66
r99 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=1.53
+ $X2=7.18 $Y2=1.53
r100 26 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.855 $Y=1.53
+ $X2=8.02 $Y2=1.53
r101 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.855 $Y=1.53
+ $X2=7.345 $Y2=1.53
r102 22 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=1.615
+ $X2=7.18 $Y2=1.53
r103 22 24 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.18 $Y=1.615
+ $X2=7.18 $Y2=1.66
r104 20 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=1.53
+ $X2=7.18 $Y2=1.53
r105 20 21 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.015 $Y=1.53
+ $X2=6.505 $Y2=1.53
r106 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.34 $Y=1.615
+ $X2=6.505 $Y2=1.53
r107 16 18 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.34 $Y=1.615
+ $X2=6.34 $Y2=1.66
r108 5 48 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.565
+ $Y=1.485 $X2=9.7 $Y2=2.34
r109 5 46 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=9.565
+ $Y=1.485 $X2=9.7 $Y2=1.66
r110 4 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=2.34
r111 4 38 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=1.66
r112 3 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=2.34
r113 3 30 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=1.66
r114 2 24 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=1.66
r115 1 18 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=6.215
+ $Y=1.485 $X2=6.34 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 44 50 53 54 55 58 60 64 66 70 72 76 78 82 84 88 90 94 96 100 102 106 112 113
+ 114 115 116 117 118 119
c227 66 0 1.18248e-19 $X=4.815 $Y=0.82
c228 3 0 7.2785e-20 $X=1.805 $Y=0.235
r229 104 106 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=9.7 $Y=0.735
+ $X2=9.7 $Y2=0.38
r230 103 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=0.82
+ $X2=8.86 $Y2=0.82
r231 102 104 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.535 $Y=0.82
+ $X2=9.7 $Y2=0.735
r232 102 103 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.535 $Y=0.82
+ $X2=9.025 $Y2=0.82
r233 98 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=0.735
+ $X2=8.86 $Y2=0.82
r234 98 100 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.86 $Y=0.735
+ $X2=8.86 $Y2=0.38
r235 97 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=0.82
+ $X2=8.02 $Y2=0.82
r236 96 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=0.82
+ $X2=8.86 $Y2=0.82
r237 96 97 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.695 $Y=0.82
+ $X2=8.185 $Y2=0.82
r238 92 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=0.735
+ $X2=8.02 $Y2=0.82
r239 92 94 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.02 $Y=0.735
+ $X2=8.02 $Y2=0.38
r240 91 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.345 $Y=0.82
+ $X2=7.18 $Y2=0.82
r241 90 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.855 $Y=0.82
+ $X2=8.02 $Y2=0.82
r242 90 91 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.855 $Y=0.82
+ $X2=7.345 $Y2=0.82
r243 86 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0.735
+ $X2=7.18 $Y2=0.82
r244 86 88 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=7.18 $Y=0.735
+ $X2=7.18 $Y2=0.38
r245 85 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=0.82
+ $X2=6.34 $Y2=0.82
r246 84 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=0.82
+ $X2=7.18 $Y2=0.82
r247 84 85 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.015 $Y=0.82
+ $X2=6.505 $Y2=0.82
r248 80 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=0.735
+ $X2=6.34 $Y2=0.82
r249 80 82 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.34 $Y=0.735
+ $X2=6.34 $Y2=0.38
r250 79 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=0.82
+ $X2=5.82 $Y2=0.82
r251 78 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=0.82
+ $X2=6.34 $Y2=0.82
r252 78 79 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.175 $Y=0.82
+ $X2=5.985 $Y2=0.82
r253 74 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.735
+ $X2=5.82 $Y2=0.82
r254 74 76 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.82 $Y=0.735
+ $X2=5.82 $Y2=0.38
r255 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=0.82
+ $X2=4.98 $Y2=0.82
r256 72 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=0.82
+ $X2=5.82 $Y2=0.82
r257 72 73 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.655 $Y=0.82
+ $X2=5.145 $Y2=0.82
r258 68 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=0.735
+ $X2=4.98 $Y2=0.82
r259 68 70 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.98 $Y=0.735
+ $X2=4.98 $Y2=0.38
r260 67 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0.82
+ $X2=4.14 $Y2=0.82
r261 66 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0.82
+ $X2=4.98 $Y2=0.82
r262 66 67 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.815 $Y=0.82
+ $X2=4.305 $Y2=0.82
r263 62 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.735
+ $X2=4.14 $Y2=0.82
r264 62 64 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.14 $Y=0.735
+ $X2=4.14 $Y2=0.38
r265 61 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0.82
+ $X2=3.3 $Y2=0.82
r266 60 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0.82
+ $X2=4.14 $Y2=0.82
r267 60 61 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=0.82
+ $X2=3.465 $Y2=0.82
r268 56 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.735
+ $X2=3.3 $Y2=0.82
r269 56 58 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.3 $Y=0.735
+ $X2=3.3 $Y2=0.38
r270 54 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0.82
+ $X2=3.3 $Y2=0.82
r271 54 55 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.135 $Y=0.82
+ $X2=2.625 $Y2=0.82
r272 51 55 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=2.487 $Y=0.735
+ $X2=2.625 $Y2=0.82
r273 51 53 0.628605 $w=2.73e-07 $l=1.5e-08 $layer=LI1_cond $X=2.487 $Y=0.735
+ $X2=2.487 $Y2=0.72
r274 50 111 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=2.487 $Y=0.465
+ $X2=2.487 $Y2=0.36
r275 50 53 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=2.487 $Y=0.465
+ $X2=2.487 $Y2=0.72
r276 47 49 44.3636 $w=2.08e-07 $l=8.4e-07 $layer=LI1_cond $X=1.1 $Y=0.36
+ $X2=1.94 $Y2=0.36
r277 45 109 3.8266 $w=2.1e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=0.215 $Y2=0.36
r278 45 47 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=1.1 $Y2=0.36
r279 44 111 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=2.35 $Y=0.36
+ $X2=2.487 $Y2=0.36
r280 44 49 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.35 $Y=0.36
+ $X2=1.94 $Y2=0.36
r281 40 109 3.09071 $w=2.6e-07 $l=1.05e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.36
r282 40 42 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.72
r283 13 106 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=9.565
+ $Y=0.235 $X2=9.7 $Y2=0.38
r284 12 100 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.725
+ $Y=0.235 $X2=8.86 $Y2=0.38
r285 11 94 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.38
r286 10 88 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.045
+ $Y=0.235 $X2=7.18 $Y2=0.38
r287 9 82 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.215
+ $Y=0.235 $X2=6.34 $Y2=0.38
r288 8 76 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.685
+ $Y=0.235 $X2=5.82 $Y2=0.38
r289 7 70 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.845
+ $Y=0.235 $X2=4.98 $Y2=0.38
r290 6 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.005
+ $Y=0.235 $X2=4.14 $Y2=0.38
r291 5 58 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.165
+ $Y=0.235 $X2=3.3 $Y2=0.38
r292 4 111 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.38
r293 4 53 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.72
r294 3 49 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r295 2 47 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.38
r296 1 109 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r297 1 42 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__O41AI_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 45 49 53
+ 57 60 61 63 64 66 67 69 70 71 72 74 75 77 78 79 111 112 115
r163 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r164 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r165 109 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r166 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r167 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r168 106 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r169 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r170 103 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=0 $X2=7.6
+ $Y2=0
r171 103 105 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.685 $Y=0
+ $X2=8.05 $Y2=0
r172 102 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r173 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r174 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r175 98 101 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r176 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r177 96 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r178 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r179 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r180 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r181 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r182 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r183 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r184 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r185 82 86 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r186 79 87 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r187 79 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r188 77 108 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=8.97 $Y2=0
r189 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.195 $Y=0 $X2=9.28
+ $Y2=0
r190 76 111 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=9.89 $Y2=0
r191 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.28
+ $Y2=0
r192 74 105 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.355 $Y=0
+ $X2=8.05 $Y2=0
r193 74 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0 $X2=8.44
+ $Y2=0
r194 73 108 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.525 $Y=0
+ $X2=8.97 $Y2=0
r195 73 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.44
+ $Y2=0
r196 71 101 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.67
+ $Y2=0
r197 71 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.76
+ $Y2=0
r198 69 95 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.29
+ $Y2=0
r199 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.4
+ $Y2=0
r200 68 98 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.485 $Y=0
+ $X2=5.75 $Y2=0
r201 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.4
+ $Y2=0
r202 66 92 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.475 $Y=0
+ $X2=4.37 $Y2=0
r203 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.56
+ $Y2=0
r204 65 95 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=5.29 $Y2=0
r205 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=0 $X2=4.56
+ $Y2=0
r206 63 89 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.635 $Y=0
+ $X2=3.45 $Y2=0
r207 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.72
+ $Y2=0
r208 62 92 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=4.37
+ $Y2=0
r209 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.72
+ $Y2=0
r210 60 86 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.53 $Y2=0
r211 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.88
+ $Y2=0
r212 59 89 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.965 $Y=0
+ $X2=3.45 $Y2=0
r213 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.88
+ $Y2=0
r214 55 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0
r215 55 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0.38
r216 51 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0
r217 51 53 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0.38
r218 47 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0
r219 47 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.6 $Y=0.085
+ $X2=7.6 $Y2=0.38
r220 46 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=0 $X2=6.76
+ $Y2=0
r221 45 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=0 $X2=7.6
+ $Y2=0
r222 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.515 $Y=0
+ $X2=6.845 $Y2=0
r223 41 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=0.085
+ $X2=6.76 $Y2=0
r224 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.76 $Y=0.085
+ $X2=6.76 $Y2=0.38
r225 37 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.4 $Y=0.085 $X2=5.4
+ $Y2=0
r226 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.4 $Y=0.085
+ $X2=5.4 $Y2=0.38
r227 33 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0
r228 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.56 $Y=0.085
+ $X2=4.56 $Y2=0.38
r229 29 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r230 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.38
r231 25 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0
r232 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.88 $Y=0.085
+ $X2=2.88 $Y2=0.38
r233 8 57 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.145
+ $Y=0.235 $X2=9.28 $Y2=0.38
r234 7 53 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.38
r235 6 49 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.465
+ $Y=0.235 $X2=7.6 $Y2=0.38
r236 5 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.38
r237 4 39 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.235 $X2=5.4 $Y2=0.38
r238 3 35 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.38
r239 2 31 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
r240 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.38
.ends


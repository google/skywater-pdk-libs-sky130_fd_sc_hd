* File: sky130_fd_sc_hd__a211oi_2.spice.SKY130_FD_SC_HD__A211OI_2.pxi
* Created: Thu Aug 27 13:59:49 2020
* 
x_PM_SKY130_FD_SC_HD__A211OI_2%C1 N_C1_c_74_n N_C1_M1002_g N_C1_M1009_g
+ N_C1_c_75_n N_C1_M1007_g N_C1_M1015_g C1 C1 N_C1_c_76_n N_C1_c_77_n
+ PM_SKY130_FD_SC_HD__A211OI_2%C1
x_PM_SKY130_FD_SC_HD__A211OI_2%B1 N_B1_c_116_n N_B1_M1005_g N_B1_M1003_g
+ N_B1_c_117_n N_B1_M1012_g N_B1_M1010_g B1 B1 B1 N_B1_c_120_n N_B1_c_121_n
+ PM_SKY130_FD_SC_HD__A211OI_2%B1
x_PM_SKY130_FD_SC_HD__A211OI_2%A1 N_A1_c_169_n N_A1_M1008_g N_A1_M1004_g
+ N_A1_c_170_n N_A1_M1013_g N_A1_M1011_g A1 A1 N_A1_c_172_n
+ PM_SKY130_FD_SC_HD__A211OI_2%A1
x_PM_SKY130_FD_SC_HD__A211OI_2%A2 N_A2_c_210_n N_A2_M1000_g N_A2_M1001_g
+ N_A2_c_211_n N_A2_M1006_g N_A2_M1014_g A2 A2 A2 N_A2_c_213_n N_A2_c_223_n
+ N_A2_c_214_n PM_SKY130_FD_SC_HD__A211OI_2%A2
x_PM_SKY130_FD_SC_HD__A211OI_2%A_37_297# N_A_37_297#_M1009_s N_A_37_297#_M1015_s
+ N_A_37_297#_M1010_d N_A_37_297#_c_250_n N_A_37_297#_c_257_n
+ N_A_37_297#_c_251_n N_A_37_297#_c_260_n N_A_37_297#_c_261_n
+ N_A_37_297#_c_252_n N_A_37_297#_c_253_n N_A_37_297#_c_276_p
+ PM_SKY130_FD_SC_HD__A211OI_2%A_37_297#
x_PM_SKY130_FD_SC_HD__A211OI_2%Y N_Y_M1002_d N_Y_M1005_s N_Y_M1008_d N_Y_M1009_d
+ N_Y_c_288_n N_Y_c_285_n N_Y_c_303_n Y Y Y Y Y Y N_Y_c_297_n
+ PM_SKY130_FD_SC_HD__A211OI_2%Y
x_PM_SKY130_FD_SC_HD__A211OI_2%A_292_297# N_A_292_297#_M1003_s
+ N_A_292_297#_M1004_s N_A_292_297#_M1001_s N_A_292_297#_c_338_n
+ N_A_292_297#_c_373_p N_A_292_297#_c_339_n N_A_292_297#_c_340_n
+ N_A_292_297#_c_374_p N_A_292_297#_c_341_n N_A_292_297#_c_342_n
+ PM_SKY130_FD_SC_HD__A211OI_2%A_292_297#
x_PM_SKY130_FD_SC_HD__A211OI_2%VPWR N_VPWR_M1004_d N_VPWR_M1011_d N_VPWR_M1014_d
+ N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n
+ N_VPWR_c_388_n VPWR N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n
+ N_VPWR_c_382_n VPWR PM_SKY130_FD_SC_HD__A211OI_2%VPWR
x_PM_SKY130_FD_SC_HD__A211OI_2%VGND N_VGND_M1002_s N_VGND_M1007_s N_VGND_M1012_d
+ N_VGND_M1000_d N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n
+ N_VGND_c_448_n VGND N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ VGND PM_SKY130_FD_SC_HD__A211OI_2%VGND
x_PM_SKY130_FD_SC_HD__A211OI_2%A_485_47# N_A_485_47#_M1008_s N_A_485_47#_M1013_s
+ N_A_485_47#_M1006_s N_A_485_47#_c_517_n N_A_485_47#_c_518_n
+ N_A_485_47#_c_531_n N_A_485_47#_c_519_n PM_SKY130_FD_SC_HD__A211OI_2%A_485_47#
cc_1 VNB N_C1_c_74_n 0.0216096f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_2 VNB N_C1_c_75_n 0.0161657f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_C1_c_76_n 0.0160237f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_4 VNB N_C1_c_77_n 0.0545373f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.16
cc_5 VNB N_B1_c_116_n 0.0161947f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_6 VNB N_B1_c_117_n 0.0212151f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_7 VNB B1 3.55996e-19 $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.445
cc_8 VNB B1 0.00228294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_120_n 0.0347254f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.16
cc_10 VNB N_B1_c_121_n 0.00445813f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.19
cc_11 VNB N_A1_c_169_n 0.0220814f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_12 VNB N_A1_c_170_n 0.0164438f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_13 VNB A1 0.00382387f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.445
cc_14 VNB N_A1_c_172_n 0.049908f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.16
cc_15 VNB N_A2_c_210_n 0.0162447f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.995
cc_16 VNB N_A2_c_211_n 0.0218823f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_17 VNB A2 7.0678e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_213_n 0.0528524f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.19
cc_19 VNB N_A2_c_214_n 0.0130932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_285_n 0.00909221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB Y 0.0010466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_382_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_444_n 0.011635f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.985
cc_24 VNB N_VGND_c_445_n 0.0265578f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.105
cc_25 VNB N_VGND_c_446_n 3.22457e-19 $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_26 VNB N_VGND_c_447_n 0.00545368f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_27 VNB N_VGND_c_448_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_449_n 0.0150118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_450_n 0.0115717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_451_n 0.0341603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_452_n 0.0169345f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_453_n 0.245166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_454_n 0.00436214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_455_n 0.00510188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_456_n 0.00436092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_485_47#_c_517_n 0.00253853f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.56
cc_37 VNB N_A_485_47#_c_518_n 0.00964039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_485_47#_c_519_n 0.0141126f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_39 VPB N_C1_M1009_g 0.0213135f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.985
cc_40 VPB N_C1_M1015_g 0.0189631f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_41 VPB N_C1_c_76_n 0.0148894f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_42 VPB N_C1_c_77_n 0.014379f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.16
cc_43 VPB N_B1_M1003_g 0.0188751f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.985
cc_44 VPB N_B1_M1010_g 0.0253813f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_45 VPB B1 0.00335108f $X=-0.19 $Y=1.305 $X2=0.125 $Y2=1.445
cc_46 VPB N_B1_c_120_n 0.004558f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.16
cc_47 VPB N_A1_M1004_g 0.0253911f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.985
cc_48 VPB N_A1_M1011_g 0.0187394f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_49 VPB N_A1_c_172_n 0.0115351f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.16
cc_50 VPB N_A2_M1001_g 0.0187334f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.985
cc_51 VPB N_A2_M1014_g 0.0219845f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_52 VPB A2 0.0192321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A2_c_213_n 0.0134886f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.19
cc_54 VPB N_A_37_297#_c_250_n 0.0191356f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_55 VPB N_A_37_297#_c_251_n 0.00746418f $X=-0.19 $Y=1.305 $X2=0.125 $Y2=1.105
cc_56 VPB N_A_37_297#_c_252_n 0.00245421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_37_297#_c_253_n 0.0047302f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.16
cc_58 VPB Y 9.40669e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_292_297#_c_338_n 0.0197398f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_60 VPB N_A_292_297#_c_339_n 0.00551179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_292_297#_c_340_n 0.00269649f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_62 VPB N_A_292_297#_c_341_n 0.00229067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_292_297#_c_342_n 0.00244502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_383_n 0.00449918f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.985
cc_65 VPB N_VPWR_c_384_n 0.00391697f $X=-0.19 $Y=1.305 $X2=0.125 $Y2=1.445
cc_66 VPB N_VPWR_c_385_n 0.0134573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_386_n 0.00449918f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_68 VPB N_VPWR_c_387_n 0.017463f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_69 VPB N_VPWR_c_388_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.16
cc_70 VPB N_VPWR_c_389_n 0.0605569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_390_n 0.017463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_391_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_382_n 0.0595597f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_C1_c_75_n N_B1_c_116_n 0.0207423f $X=0.955 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_75 N_C1_M1015_g N_B1_M1003_g 0.0207423f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_76 N_C1_c_77_n B1 0.00230308f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C1_c_77_n N_B1_c_120_n 0.0207423f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C1_c_77_n N_B1_c_121_n 0.00280717f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C1_c_76_n N_A_37_297#_M1009_s 0.00356172f $X=0.315 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_80 N_C1_c_76_n N_A_37_297#_c_250_n 0.0222304f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_81 N_C1_c_77_n N_A_37_297#_c_250_n 9.19108e-19 $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C1_M1009_g N_A_37_297#_c_257_n 0.0115808f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_83 N_C1_M1015_g N_A_37_297#_c_257_n 0.0115808f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_84 N_C1_c_75_n N_Y_c_288_n 0.0150488f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_85 N_C1_c_74_n Y 0.0105578f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_86 N_C1_M1009_g Y 0.0118058f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_87 N_C1_c_75_n Y 0.0029727f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_88 N_C1_M1015_g Y 0.00126907f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_89 N_C1_c_76_n Y 0.0414198f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_90 N_C1_c_77_n Y 0.0215468f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_91 N_C1_M1009_g Y 0.00374759f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_92 N_C1_M1015_g Y 0.00465665f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_93 N_C1_c_74_n N_Y_c_297_n 0.00455058f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_94 N_C1_M1015_g N_A_292_297#_c_341_n 4.06986e-19 $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_95 N_C1_M1009_g N_VPWR_c_389_n 0.00359964f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_96 N_C1_M1015_g N_VPWR_c_389_n 0.00359964f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_97 N_C1_M1009_g N_VPWR_c_382_n 0.00625772f $X=0.525 $Y=1.985 $X2=0 $Y2=0
cc_98 N_C1_M1015_g N_VPWR_c_382_n 0.00530646f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_99 N_C1_c_74_n N_VGND_c_445_n 0.00673673f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_100 N_C1_c_76_n N_VGND_c_445_n 0.02077f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_101 N_C1_c_77_n N_VGND_c_445_n 0.00167802f $X=0.955 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C1_c_74_n N_VGND_c_446_n 4.76231e-19 $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_103 N_C1_c_75_n N_VGND_c_446_n 0.00671303f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_104 N_C1_c_74_n N_VGND_c_449_n 0.0054895f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C1_c_75_n N_VGND_c_449_n 0.00355956f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_106 N_C1_c_74_n N_VGND_c_453_n 0.0108426f $X=0.525 $Y=0.995 $X2=0 $Y2=0
cc_107 N_C1_c_75_n N_VGND_c_453_n 0.00415355f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_108 B1 A1 0.00867894f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B1_c_120_n A1 0.00241506f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_110 B1 N_A1_c_172_n 2.31323e-19 $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B1_c_120_n N_A1_c_172_n 0.00766527f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_112 B1 N_A_37_297#_M1015_s 0.00302257f $X=1.045 $Y=1.445 $X2=0 $Y2=0
cc_113 B1 N_A_37_297#_c_260_n 0.0147759f $X=1.045 $Y=1.445 $X2=0 $Y2=0
cc_114 N_B1_M1003_g N_A_37_297#_c_261_n 0.0124676f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_115 N_B1_M1010_g N_A_37_297#_c_261_n 0.0102357f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_116 N_B1_c_116_n N_Y_c_288_n 0.0115344f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_117 B1 N_Y_c_288_n 0.0137473f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B1_c_121_n N_Y_c_288_n 0.0155699f $X=1.145 $Y=1.285 $X2=0 $Y2=0
cc_119 N_B1_c_117_n N_Y_c_285_n 0.0153909f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_120 B1 N_Y_c_285_n 0.00458497f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_121 B1 N_Y_c_303_n 0.0135093f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B1_c_120_n N_Y_c_303_n 0.00241526f $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_123 B1 Y 0.0150355f $X=1.045 $Y=1.445 $X2=0 $Y2=0
cc_124 N_B1_c_120_n Y 3.83894e-19 $X=1.815 $Y=1.16 $X2=0 $Y2=0
cc_125 N_B1_c_121_n Y 0.0199672f $X=1.145 $Y=1.285 $X2=0 $Y2=0
cc_126 N_B1_M1010_g N_A_292_297#_c_338_n 0.0136412f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_127 B1 N_A_292_297#_c_338_n 0.0013794f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_M1003_g N_A_292_297#_c_341_n 0.00871063f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_129 N_B1_M1010_g N_A_292_297#_c_341_n 0.0118005f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_130 B1 N_A_292_297#_c_341_n 0.00753021f $X=1.045 $Y=1.445 $X2=0 $Y2=0
cc_131 B1 N_A_292_297#_c_341_n 0.0268811f $X=1.505 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B1_c_120_n N_A_292_297#_c_341_n 0.00243382f $X=1.815 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_B1_M1010_g N_VPWR_c_383_n 0.00220691f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_134 N_B1_M1003_g N_VPWR_c_389_n 0.00359964f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B1_M1010_g N_VPWR_c_389_n 0.00359964f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B1_M1003_g N_VPWR_c_382_n 0.00530646f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B1_M1010_g N_VPWR_c_382_n 0.00658082f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B1_c_116_n N_VGND_c_446_n 0.00675326f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_117_n N_VGND_c_446_n 6.26587e-19 $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_116_n N_VGND_c_447_n 6.26587e-19 $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_117_n N_VGND_c_447_n 0.00785251f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B1_c_116_n N_VGND_c_450_n 0.00355956f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B1_c_117_n N_VGND_c_450_n 0.00355956f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B1_c_116_n N_VGND_c_453_n 0.00419786f $X=1.385 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B1_c_117_n N_VGND_c_453_n 0.00419786f $X=1.815 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_c_170_n N_A2_c_210_n 0.0232066f $X=3.195 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A1_M1011_g N_A2_M1001_g 0.0232066f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_148 A1 N_A2_c_213_n 8.79505e-19 $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A1_c_172_n N_A2_c_213_n 0.0232066f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_150 A1 N_A2_c_223_n 0.00673927f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A1_c_172_n N_A2_c_223_n 8.79437e-19 $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A1_c_169_n N_Y_c_285_n 0.0117564f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_170_n N_Y_c_285_n 0.00304782f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_154 A1 N_Y_c_285_n 0.0449091f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A1_c_172_n N_Y_c_285_n 0.00852911f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_M1004_g N_A_292_297#_c_338_n 0.0166683f $X=2.765 $Y=1.985 $X2=0
+ $Y2=0
cc_157 A1 N_A_292_297#_c_338_n 0.0349893f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A1_c_172_n N_A_292_297#_c_338_n 0.00636978f $X=3.195 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A1_M1011_g N_A_292_297#_c_339_n 0.018462f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_160 A1 N_A_292_297#_c_342_n 0.0194515f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_172_n N_A_292_297#_c_342_n 0.0024449f $X=3.195 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A1_M1004_g N_VPWR_c_383_n 0.0033198f $X=2.765 $Y=1.985 $X2=0 $Y2=0
cc_163 N_A1_M1011_g N_VPWR_c_384_n 0.00157243f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A1_M1004_g N_VPWR_c_387_n 0.00585385f $X=2.765 $Y=1.985 $X2=0 $Y2=0
cc_165 N_A1_M1011_g N_VPWR_c_387_n 0.00585385f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A1_M1004_g N_VPWR_c_382_n 0.0118268f $X=2.765 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_M1011_g N_VPWR_c_382_n 0.0105525f $X=3.195 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_c_169_n N_VGND_c_447_n 0.00248811f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_170_n N_VGND_c_448_n 0.00125518f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_169_n N_VGND_c_451_n 0.00359964f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_170_n N_VGND_c_451_n 0.00359964f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A1_c_169_n N_VGND_c_453_n 0.00658082f $X=2.765 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_170_n N_VGND_c_453_n 0.00534735f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_169_n N_A_485_47#_c_517_n 0.00881608f $X=2.765 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A1_c_170_n N_A_485_47#_c_517_n 0.0134173f $X=3.195 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_A_292_297#_c_339_n 0.0162109f $X=3.625 $Y=1.985 $X2=0
+ $Y2=0
cc_177 N_A2_M1014_g N_A_292_297#_c_340_n 2.85064e-19 $X=4.055 $Y=1.985 $X2=0
+ $Y2=0
cc_178 A2 N_A_292_297#_c_340_n 0.00228239f $X=4.285 $Y=1.445 $X2=0 $Y2=0
cc_179 N_A2_c_213_n N_A_292_297#_c_340_n 0.0024449f $X=4.265 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A2_c_223_n N_A_292_297#_c_340_n 0.0194515f $X=4.175 $Y=1.16 $X2=0 $Y2=0
cc_181 A2 N_VPWR_M1014_d 0.00444487f $X=4.285 $Y=1.445 $X2=0 $Y2=0
cc_182 N_A2_M1001_g N_VPWR_c_384_n 0.00157243f $X=3.625 $Y=1.985 $X2=0 $Y2=0
cc_183 N_A2_M1014_g N_VPWR_c_386_n 0.0033198f $X=4.055 $Y=1.985 $X2=0 $Y2=0
cc_184 A2 N_VPWR_c_386_n 0.0168982f $X=4.285 $Y=1.445 $X2=0 $Y2=0
cc_185 N_A2_c_213_n N_VPWR_c_386_n 8.03343e-19 $X=4.265 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_VPWR_c_390_n 0.00585385f $X=3.625 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A2_M1014_g N_VPWR_c_390_n 0.00585385f $X=4.055 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A2_M1001_g N_VPWR_c_382_n 0.0105525f $X=3.625 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A2_M1014_g N_VPWR_c_382_n 0.0115195f $X=4.055 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A2_c_210_n N_VGND_c_448_n 0.00763332f $X=3.625 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_211_n N_VGND_c_448_n 0.00838216f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_210_n N_VGND_c_451_n 0.00353537f $X=3.625 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_211_n N_VGND_c_452_n 0.00353537f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_210_n N_VGND_c_453_n 0.00418339f $X=3.625 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_211_n N_VGND_c_453_n 0.00518765f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_210_n N_A_485_47#_c_518_n 0.0141171f $X=3.625 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_211_n N_A_485_47#_c_518_n 0.0131275f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_213_n N_A_485_47#_c_518_n 0.00753832f $X=4.265 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A2_c_223_n N_A_485_47#_c_518_n 0.0259645f $X=4.175 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_214_n N_A_485_47#_c_518_n 0.0206749f $X=4.337 $Y=1.285 $X2=0 $Y2=0
cc_201 N_A_37_297#_c_257_n N_Y_M1009_d 0.00340138f $X=1.075 $Y=2.37 $X2=0 $Y2=0
cc_202 N_A_37_297#_c_257_n Y 0.0151669f $X=1.075 $Y=2.37 $X2=0 $Y2=0
cc_203 N_A_37_297#_c_261_n N_A_292_297#_M1003_s 0.00341854f $X=1.935 $Y=2.355
+ $X2=-0.19 $Y2=1.305
cc_204 N_A_37_297#_M1010_d N_A_292_297#_c_338_n 0.0030713f $X=1.89 $Y=1.485
+ $X2=0 $Y2=0
cc_205 N_A_37_297#_c_261_n N_A_292_297#_c_338_n 0.00303673f $X=1.935 $Y=2.355
+ $X2=0 $Y2=0
cc_206 N_A_37_297#_c_253_n N_A_292_297#_c_338_n 0.0210743f $X=2.03 $Y=2 $X2=0
+ $Y2=0
cc_207 N_A_37_297#_c_261_n N_A_292_297#_c_341_n 0.0154266f $X=1.935 $Y=2.355
+ $X2=0 $Y2=0
cc_208 N_A_37_297#_c_252_n N_VPWR_c_383_n 0.0140847f $X=2.075 $Y=2.255 $X2=0
+ $Y2=0
cc_209 N_A_37_297#_c_253_n N_VPWR_c_383_n 0.0273982f $X=2.03 $Y=2 $X2=0 $Y2=0
cc_210 N_A_37_297#_c_257_n N_VPWR_c_389_n 0.0339793f $X=1.075 $Y=2.37 $X2=0
+ $Y2=0
cc_211 N_A_37_297#_c_251_n N_VPWR_c_389_n 0.0168262f $X=0.405 $Y=2.37 $X2=0
+ $Y2=0
cc_212 N_A_37_297#_c_261_n N_VPWR_c_389_n 0.0342716f $X=1.935 $Y=2.355 $X2=0
+ $Y2=0
cc_213 N_A_37_297#_c_252_n N_VPWR_c_389_n 0.018073f $X=2.075 $Y=2.255 $X2=0
+ $Y2=0
cc_214 N_A_37_297#_c_276_p N_VPWR_c_389_n 0.0117613f $X=1.17 $Y=2.355 $X2=0
+ $Y2=0
cc_215 N_A_37_297#_M1009_s N_VPWR_c_382_n 0.00213754f $X=0.185 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_A_37_297#_M1015_s N_VPWR_c_382_n 0.00223591f $X=1.03 $Y=1.485 $X2=0
+ $Y2=0
cc_217 N_A_37_297#_M1010_d N_VPWR_c_382_n 0.00213754f $X=1.89 $Y=1.485 $X2=0
+ $Y2=0
cc_218 N_A_37_297#_c_257_n N_VPWR_c_382_n 0.0232862f $X=1.075 $Y=2.37 $X2=0
+ $Y2=0
cc_219 N_A_37_297#_c_251_n N_VPWR_c_382_n 0.00995632f $X=0.405 $Y=2.37 $X2=0
+ $Y2=0
cc_220 N_A_37_297#_c_261_n N_VPWR_c_382_n 0.0233735f $X=1.935 $Y=2.355 $X2=0
+ $Y2=0
cc_221 N_A_37_297#_c_252_n N_VPWR_c_382_n 0.0107056f $X=2.075 $Y=2.255 $X2=0
+ $Y2=0
cc_222 N_A_37_297#_c_276_p N_VPWR_c_382_n 0.00727972f $X=1.17 $Y=2.355 $X2=0
+ $Y2=0
cc_223 N_Y_c_285_n N_A_292_297#_c_338_n 0.016748f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_224 N_Y_c_285_n N_A_292_297#_c_339_n 6.64236e-19 $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_225 N_Y_M1009_d N_VPWR_c_382_n 0.0022523f $X=0.6 $Y=1.485 $X2=0 $Y2=0
cc_226 N_Y_c_288_n N_VGND_M1007_s 0.00356881f $X=1.505 $Y=0.755 $X2=0 $Y2=0
cc_227 N_Y_c_285_n N_VGND_M1012_d 0.00729184f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_228 N_Y_c_288_n N_VGND_c_446_n 0.0154687f $X=1.505 $Y=0.755 $X2=0 $Y2=0
cc_229 N_Y_c_285_n N_VGND_c_447_n 0.0199465f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_230 N_Y_c_288_n N_VGND_c_449_n 0.00218985f $X=1.505 $Y=0.755 $X2=0 $Y2=0
cc_231 N_Y_c_297_n N_VGND_c_449_n 0.0156896f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_232 N_Y_c_288_n N_VGND_c_450_n 0.00237557f $X=1.505 $Y=0.755 $X2=0 $Y2=0
cc_233 N_Y_c_285_n N_VGND_c_450_n 0.00237557f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_234 Y N_VGND_c_450_n 0.0103239f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_235 N_Y_c_285_n N_VGND_c_451_n 0.00335954f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_236 N_Y_M1002_d N_VGND_c_453_n 0.00239726f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_237 N_Y_M1005_s N_VGND_c_453_n 0.00259724f $X=1.46 $Y=0.235 $X2=0 $Y2=0
cc_238 N_Y_M1008_d N_VGND_c_453_n 0.0022523f $X=2.84 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_288_n N_VGND_c_453_n 0.00916746f $X=1.505 $Y=0.755 $X2=0 $Y2=0
cc_240 N_Y_c_285_n N_VGND_c_453_n 0.0124734f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_241 Y N_VGND_c_453_n 5.9298e-19 $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_242 Y N_VGND_c_453_n 0.00709824f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_243 N_Y_c_297_n N_VGND_c_453_n 0.00975383f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_244 N_Y_c_285_n N_A_485_47#_M1008_s 0.0049028f $X=2.98 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_245 N_Y_M1008_d N_A_485_47#_c_517_n 0.00331038f $X=2.84 $Y=0.235 $X2=0 $Y2=0
cc_246 N_Y_c_285_n N_A_485_47#_c_517_n 0.0390804f $X=2.98 $Y=0.755 $X2=0 $Y2=0
cc_247 N_A_292_297#_c_338_n N_VPWR_M1004_d 0.00337897f $X=2.845 $Y=1.555
+ $X2=-0.19 $Y2=1.305
cc_248 N_A_292_297#_c_339_n N_VPWR_M1011_d 0.00181657f $X=3.705 $Y=1.555 $X2=0
+ $Y2=0
cc_249 N_A_292_297#_c_338_n N_VPWR_c_383_n 0.0155267f $X=2.845 $Y=1.555 $X2=0
+ $Y2=0
cc_250 N_A_292_297#_c_339_n N_VPWR_c_384_n 0.0130834f $X=3.705 $Y=1.555 $X2=0
+ $Y2=0
cc_251 N_A_292_297#_c_373_p N_VPWR_c_387_n 0.0152923f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_252 N_A_292_297#_c_374_p N_VPWR_c_390_n 0.0152923f $X=3.84 $Y=2.3 $X2=0 $Y2=0
cc_253 N_A_292_297#_M1003_s N_VPWR_c_382_n 0.0022523f $X=1.46 $Y=1.485 $X2=0
+ $Y2=0
cc_254 N_A_292_297#_M1004_s N_VPWR_c_382_n 0.00257947f $X=2.84 $Y=1.485 $X2=0
+ $Y2=0
cc_255 N_A_292_297#_M1001_s N_VPWR_c_382_n 0.00257947f $X=3.7 $Y=1.485 $X2=0
+ $Y2=0
cc_256 N_A_292_297#_c_373_p N_VPWR_c_382_n 0.0103212f $X=2.98 $Y=2.3 $X2=0 $Y2=0
cc_257 N_A_292_297#_c_374_p N_VPWR_c_382_n 0.0103212f $X=3.84 $Y=2.3 $X2=0 $Y2=0
cc_258 N_A_292_297#_c_339_n N_A_485_47#_c_518_n 0.00464805f $X=3.705 $Y=1.555
+ $X2=0 $Y2=0
cc_259 N_A_292_297#_c_339_n N_A_485_47#_c_531_n 0.00556674f $X=3.705 $Y=1.555
+ $X2=0 $Y2=0
cc_260 N_VGND_c_453_n N_A_485_47#_M1008_s 0.00213789f $X=4.37 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_261 N_VGND_c_453_n N_A_485_47#_M1013_s 0.00245191f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_453_n N_A_485_47#_M1006_s 0.00233744f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_447_n N_A_485_47#_c_517_n 0.017007f $X=2.03 $Y=0.38 $X2=0 $Y2=0
cc_264 N_VGND_c_451_n N_A_485_47#_c_517_n 0.0611481f $X=3.675 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_453_n N_A_485_47#_c_517_n 0.039988f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_M1000_d N_A_485_47#_c_518_n 0.00333086f $X=3.7 $Y=0.235 $X2=0
+ $Y2=0
cc_267 N_VGND_c_448_n N_A_485_47#_c_518_n 0.0154649f $X=3.84 $Y=0.36 $X2=0 $Y2=0
cc_268 N_VGND_c_451_n N_A_485_47#_c_518_n 0.00260024f $X=3.675 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_452_n N_A_485_47#_c_518_n 0.00260024f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_453_n N_A_485_47#_c_518_n 0.0105918f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_271 N_VGND_c_452_n N_A_485_47#_c_519_n 0.0162389f $X=4.37 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_453_n N_A_485_47#_c_519_n 0.0094641f $X=4.37 $Y=0 $X2=0 $Y2=0

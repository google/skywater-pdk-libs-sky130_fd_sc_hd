* File: sky130_fd_sc_hd__einvp_8.spice.SKY130_FD_SC_HD__EINVP_8.pxi
* Created: Thu Aug 27 14:20:57 2020
* 
x_PM_SKY130_FD_SC_HD__EINVP_8%TE N_TE_c_133_n N_TE_M1030_g N_TE_M1023_g
+ N_TE_c_134_n N_TE_c_135_n N_TE_c_136_n N_TE_M1010_g N_TE_c_137_n N_TE_c_138_n
+ N_TE_M1012_g N_TE_c_139_n N_TE_c_140_n N_TE_M1014_g N_TE_c_141_n N_TE_c_142_n
+ N_TE_M1015_g N_TE_c_143_n N_TE_c_144_n N_TE_M1016_g N_TE_c_145_n N_TE_c_146_n
+ N_TE_M1019_g N_TE_c_147_n N_TE_c_148_n N_TE_M1020_g N_TE_c_149_n N_TE_c_150_n
+ N_TE_M1021_g N_TE_c_151_n N_TE_c_152_n N_TE_c_153_n N_TE_c_154_n N_TE_c_155_n
+ N_TE_c_156_n N_TE_c_157_n TE TE PM_SKY130_FD_SC_HD__EINVP_8%TE
x_PM_SKY130_FD_SC_HD__EINVP_8%A_27_47# N_A_27_47#_M1030_s N_A_27_47#_M1023_s
+ N_A_27_47#_c_274_n N_A_27_47#_M1000_g N_A_27_47#_c_275_n N_A_27_47#_c_276_n
+ N_A_27_47#_c_277_n N_A_27_47#_M1001_g N_A_27_47#_c_278_n N_A_27_47#_c_279_n
+ N_A_27_47#_M1005_g N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_M1008_g
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_M1009_g N_A_27_47#_c_284_n
+ N_A_27_47#_c_285_n N_A_27_47#_M1013_g N_A_27_47#_c_286_n N_A_27_47#_c_287_n
+ N_A_27_47#_M1024_g N_A_27_47#_c_288_n N_A_27_47#_M1027_g N_A_27_47#_c_289_n
+ N_A_27_47#_c_290_n N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n
+ N_A_27_47#_c_294_n N_A_27_47#_c_269_n N_A_27_47#_c_295_n N_A_27_47#_c_270_n
+ N_A_27_47#_c_271_n N_A_27_47#_c_296_n N_A_27_47#_c_272_n N_A_27_47#_c_273_n
+ N_A_27_47#_c_340_n PM_SKY130_FD_SC_HD__EINVP_8%A_27_47#
x_PM_SKY130_FD_SC_HD__EINVP_8%A N_A_c_432_n N_A_M1003_g N_A_M1002_g N_A_c_433_n
+ N_A_M1004_g N_A_M1007_g N_A_M1006_g N_A_M1017_g N_A_M1011_g N_A_M1018_g
+ N_A_c_438_n N_A_M1028_g N_A_M1022_g N_A_c_439_n N_A_M1031_g N_A_M1025_g
+ N_A_M1032_g N_A_M1026_g N_A_c_442_n N_A_M1033_g N_A_M1029_g A A A A A A
+ PM_SKY130_FD_SC_HD__EINVP_8%A
x_PM_SKY130_FD_SC_HD__EINVP_8%VPWR N_VPWR_M1023_d N_VPWR_M1000_s N_VPWR_M1005_s
+ N_VPWR_M1009_s N_VPWR_M1024_s N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n
+ N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n
+ N_VPWR_c_574_n VPWR N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n
+ N_VPWR_c_578_n N_VPWR_c_565_n N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n
+ PM_SKY130_FD_SC_HD__EINVP_8%VPWR
x_PM_SKY130_FD_SC_HD__EINVP_8%A_215_309# N_A_215_309#_M1000_d
+ N_A_215_309#_M1001_d N_A_215_309#_M1008_d N_A_215_309#_M1013_d
+ N_A_215_309#_M1027_d N_A_215_309#_M1007_s N_A_215_309#_M1018_s
+ N_A_215_309#_M1025_s N_A_215_309#_M1029_s N_A_215_309#_c_689_n
+ N_A_215_309#_c_696_n N_A_215_309#_c_686_n N_A_215_309#_c_745_n
+ N_A_215_309#_c_702_n N_A_215_309#_c_749_n N_A_215_309#_c_706_n
+ N_A_215_309#_c_753_n N_A_215_309#_c_710_n N_A_215_309#_c_720_n
+ N_A_215_309#_c_759_n N_A_215_309#_c_782_p N_A_215_309#_c_722_n
+ N_A_215_309#_c_784_p N_A_215_309#_c_724_n N_A_215_309#_c_786_p
+ N_A_215_309#_c_687_n N_A_215_309#_c_688_n N_A_215_309#_c_692_n
+ N_A_215_309#_c_693_n N_A_215_309#_c_694_n N_A_215_309#_c_767_n
+ N_A_215_309#_c_769_n N_A_215_309#_c_771_n
+ PM_SKY130_FD_SC_HD__EINVP_8%A_215_309#
x_PM_SKY130_FD_SC_HD__EINVP_8%Z N_Z_M1003_s N_Z_M1006_s N_Z_M1028_s N_Z_M1032_s
+ N_Z_M1002_d N_Z_M1017_d N_Z_M1022_d N_Z_M1026_d N_Z_c_788_n N_Z_c_807_n Z Z Z
+ Z Z Z Z Z N_Z_c_792_n Z N_Z_c_793_n N_Z_c_794_n N_Z_c_848_n
+ PM_SKY130_FD_SC_HD__EINVP_8%Z
x_PM_SKY130_FD_SC_HD__EINVP_8%VGND N_VGND_M1030_d N_VGND_M1012_d N_VGND_M1015_d
+ N_VGND_M1019_d N_VGND_M1021_d N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n
+ N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n
+ N_VGND_c_893_n N_VGND_c_894_n VGND N_VGND_c_895_n N_VGND_c_896_n
+ N_VGND_c_897_n N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n N_VGND_c_901_n
+ PM_SKY130_FD_SC_HD__EINVP_8%VGND
x_PM_SKY130_FD_SC_HD__EINVP_8%A_193_47# N_A_193_47#_M1010_s N_A_193_47#_M1014_s
+ N_A_193_47#_M1016_s N_A_193_47#_M1020_s N_A_193_47#_M1003_d
+ N_A_193_47#_M1004_d N_A_193_47#_M1011_d N_A_193_47#_M1031_d
+ N_A_193_47#_M1033_d N_A_193_47#_c_1016_n N_A_193_47#_c_1017_n
+ N_A_193_47#_c_1020_n N_A_193_47#_c_1080_n N_A_193_47#_c_1022_n
+ N_A_193_47#_c_1087_n N_A_193_47#_c_1025_n N_A_193_47#_c_1094_n
+ N_A_193_47#_c_1012_n N_A_193_47#_c_1013_n N_A_193_47#_c_1014_n
+ N_A_193_47#_c_1015_n N_A_193_47#_c_1030_n N_A_193_47#_c_1031_n
+ N_A_193_47#_c_1032_n PM_SKY130_FD_SC_HD__EINVP_8%A_193_47#
cc_1 VNB N_TE_c_133_n 0.0186243f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_2 VNB N_TE_c_134_n 0.0144728f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=1.035
cc_3 VNB N_TE_c_135_n 0.0390839f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.035
cc_4 VNB N_TE_c_136_n 0.0141775f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.96
cc_5 VNB N_TE_c_137_n 0.0152216f $X=-0.19 $Y=-0.24 $X2=1.255 $Y2=1.035
cc_6 VNB N_TE_c_138_n 0.0141947f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.96
cc_7 VNB N_TE_c_139_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.035
cc_8 VNB N_TE_c_140_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.96
cc_9 VNB N_TE_c_141_n 0.00896022f $X=-0.19 $Y=-0.24 $X2=2.095 $Y2=1.035
cc_10 VNB N_TE_c_142_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.96
cc_11 VNB N_TE_c_143_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=1.035
cc_12 VNB N_TE_c_144_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.96
cc_13 VNB N_TE_c_145_n 0.00896022f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=1.035
cc_14 VNB N_TE_c_146_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=0.96
cc_15 VNB N_TE_c_147_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=1.035
cc_16 VNB N_TE_c_148_n 0.0140273f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.96
cc_17 VNB N_TE_c_149_n 0.016072f $X=-0.19 $Y=-0.24 $X2=3.775 $Y2=1.035
cc_18 VNB N_TE_c_150_n 0.018285f $X=-0.19 $Y=-0.24 $X2=3.85 $Y2=0.96
cc_19 VNB N_TE_c_151_n 0.00661167f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.035
cc_20 VNB N_TE_c_152_n 0.0053816f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.035
cc_21 VNB N_TE_c_153_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.035
cc_22 VNB N_TE_c_154_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.035
cc_23 VNB N_TE_c_155_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=1.035
cc_24 VNB N_TE_c_156_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.035
cc_25 VNB N_TE_c_157_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=1.035
cc_26 VNB TE 0.0134173f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_A_27_47#_c_269_n 0.0156779f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_28 VNB N_A_27_47#_c_270_n 0.00754597f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_29 VNB N_A_27_47#_c_271_n 7.10498e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.142
cc_30 VNB N_A_27_47#_c_272_n 0.00764942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_273_n 0.0274243f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_c_432_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_33 VNB N_A_c_433_n 0.0155271f $X=-0.19 $Y=-0.24 $X2=0.815 $Y2=1.035
cc_34 VNB N_A_M1006_g 0.0173901f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.56
cc_35 VNB N_A_M1017_g 4.49313e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_36 VNB N_A_M1011_g 0.0174037f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.96
cc_37 VNB N_A_M1018_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=1.035
cc_38 VNB N_A_c_438_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.56
cc_39 VNB N_A_c_439_n 0.0160053f $X=-0.19 $Y=-0.24 $X2=3.355 $Y2=1.035
cc_40 VNB N_A_M1032_g 0.0174037f $X=-0.19 $Y=-0.24 $X2=3.85 $Y2=0.56
cc_41 VNB N_A_M1026_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=1.035
cc_42 VNB N_A_c_442_n 0.155475f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.035
cc_43 VNB N_A_M1033_g 0.0235825f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_44 VNB A 0.0230602f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_45 VNB N_VPWR_c_565_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Z_c_788_n 0.0105158f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=1.035
cc_47 VNB N_VGND_c_885_n 3.99129e-19 $X=-0.19 $Y=-0.24 $X2=1.675 $Y2=1.035
cc_48 VNB N_VGND_c_886_n 3.05427e-19 $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_49 VNB N_VGND_c_887_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.56
cc_50 VNB N_VGND_c_888_n 3.01744e-19 $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.96
cc_51 VNB N_VGND_c_889_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=2.59 $Y2=0.56
cc_52 VNB N_VGND_c_890_n 0.00520071f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=0.56
cc_53 VNB N_VGND_c_891_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=3.085 $Y2=1.035
cc_54 VNB N_VGND_c_892_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.96
cc_55 VNB N_VGND_c_893_n 0.0110228f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.56
cc_56 VNB N_VGND_c_894_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=3.43 $Y2=0.56
cc_57 VNB N_VGND_c_895_n 0.014319f $X=-0.19 $Y=-0.24 $X2=3.85 $Y2=0.96
cc_58 VNB N_VGND_c_896_n 0.0123936f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.035
cc_59 VNB N_VGND_c_897_n 0.0935303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_898_n 0.39278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_899_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_900_n 0.00436274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_901_n 0.00526505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_193_47#_c_1012_n 0.00608242f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.035
cc_65 VNB N_A_193_47#_c_1013_n 0.00299848f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_66 VNB N_A_193_47#_c_1014_n 0.00279976f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_67 VNB N_A_193_47#_c_1015_n 0.0102574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VPB N_TE_M1023_g 0.025505f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_69 VPB N_TE_c_135_n 0.01029f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.035
cc_70 VPB TE 0.0127315f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_71 VPB N_A_27_47#_c_274_n 0.0174982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_275_n 0.00892157f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.96
cc_73 VPB N_A_27_47#_c_276_n 0.00858091f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_74 VPB N_A_27_47#_c_277_n 0.0140273f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_75 VPB N_A_27_47#_c_278_n 0.00892095f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.96
cc_76 VPB N_A_27_47#_c_279_n 0.0140273f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_77 VPB N_A_27_47#_c_280_n 0.00892157f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.96
cc_78 VPB N_A_27_47#_c_281_n 0.0140273f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_79 VPB N_A_27_47#_c_282_n 0.00892095f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.96
cc_80 VPB N_A_27_47#_c_283_n 0.0140273f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_81 VPB N_A_27_47#_c_284_n 0.00892157f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.96
cc_82 VPB N_A_27_47#_c_285_n 0.0140273f $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.56
cc_83 VPB N_A_27_47#_c_286_n 0.00892095f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=0.96
cc_84 VPB N_A_27_47#_c_287_n 0.0140273f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=0.56
cc_85 VPB N_A_27_47#_c_288_n 0.0146322f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.96
cc_86 VPB N_A_27_47#_c_289_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.775 $Y2=1.035
cc_87 VPB N_A_27_47#_c_290_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.035
cc_88 VPB N_A_27_47#_c_291_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.85 $Y2=0.96
cc_89 VPB N_A_27_47#_c_292_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.85 $Y2=0.56
cc_90 VPB N_A_27_47#_c_293_n 0.00391059f $X=-0.19 $Y=1.305 $X2=3.85 $Y2=0.56
cc_91 VPB N_A_27_47#_c_294_n 0.0215363f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.035
cc_92 VPB N_A_27_47#_c_295_n 0.0198678f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.142
cc_93 VPB N_A_27_47#_c_296_n 0.0168153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_27_47#_c_272_n 0.0133223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_47#_c_273_n 0.00101273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_M1002_g 0.0187449f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_97 VPB N_A_M1007_g 0.0176224f $X=-0.19 $Y=1.305 $X2=1.255 $Y2=1.035
cc_98 VPB N_A_M1017_g 0.0191533f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_99 VPB N_A_M1018_g 0.0191843f $X=-0.19 $Y=1.305 $X2=2.245 $Y2=1.035
cc_100 VPB N_A_M1022_g 0.0181338f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=0.56
cc_101 VPB N_A_M1025_g 0.0181338f $X=-0.19 $Y=1.305 $X2=3.775 $Y2=1.035
cc_102 VPB N_A_M1026_g 0.0191843f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=1.035
cc_103 VPB N_A_c_442_n 0.0167135f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.035
cc_104 VPB N_A_M1029_g 0.0263683f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.142
cc_105 VPB N_VPWR_c_566_n 0.0066501f $X=-0.19 $Y=1.305 $X2=1.675 $Y2=1.035
cc_106 VPB N_VPWR_c_567_n 3.14017e-19 $X=-0.19 $Y=1.305 $X2=1.75 $Y2=0.56
cc_107 VPB N_VPWR_c_568_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.56
cc_108 VPB N_VPWR_c_569_n 3.01744e-19 $X=-0.19 $Y=1.305 $X2=2.59 $Y2=0.96
cc_109 VPB N_VPWR_c_570_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.035
cc_110 VPB N_VPWR_c_571_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=0.56
cc_111 VPB N_VPWR_c_572_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.355 $Y2=1.035
cc_112 VPB N_VPWR_c_573_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.96
cc_113 VPB N_VPWR_c_574_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.56
cc_114 VPB N_VPWR_c_575_n 0.0150576f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.035
cc_115 VPB N_VPWR_c_576_n 0.0153895f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.035
cc_116 VPB N_VPWR_c_577_n 0.0124915f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=1.035
cc_117 VPB N_VPWR_c_578_n 0.0916214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_565_n 0.0528486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_580_n 0.00565587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_581_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_582_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_215_309#_c_686_n 0.00133077f $X=-0.19 $Y=1.305 $X2=2.935
+ $Y2=1.035
cc_123 VPB N_A_215_309#_c_687_n 0.00821273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_215_309#_c_688_n 0.0367644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB Z 0.00218571f $X=-0.19 $Y=1.305 $X2=3.085 $Y2=1.035
cc_126 VPB Z 0.00223196f $X=-0.19 $Y=1.305 $X2=3.43 $Y2=0.56
cc_127 VPB Z 0.00223815f $X=-0.19 $Y=1.305 $X2=3.505 $Y2=1.035
cc_128 VPB N_Z_c_792_n 0.0026552f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_129 VPB N_Z_c_793_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_130 VPB N_Z_c_794_n 0.00218965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 TE N_A_27_47#_M1023_s 0.00429701f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_132 N_TE_c_139_n N_A_27_47#_c_275_n 0.014005f $X=1.675 $Y=1.035 $X2=0 $Y2=0
cc_133 N_TE_c_152_n N_A_27_47#_c_276_n 0.014005f $X=1.33 $Y=1.035 $X2=0 $Y2=0
cc_134 N_TE_c_141_n N_A_27_47#_c_278_n 0.014005f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_135 N_TE_c_143_n N_A_27_47#_c_280_n 0.014005f $X=2.515 $Y=1.035 $X2=0 $Y2=0
cc_136 N_TE_c_145_n N_A_27_47#_c_282_n 0.014005f $X=2.935 $Y=1.035 $X2=0 $Y2=0
cc_137 N_TE_c_147_n N_A_27_47#_c_284_n 0.014005f $X=3.355 $Y=1.035 $X2=0 $Y2=0
cc_138 N_TE_c_149_n N_A_27_47#_c_286_n 0.014005f $X=3.775 $Y=1.035 $X2=0 $Y2=0
cc_139 N_TE_c_153_n N_A_27_47#_c_289_n 0.014005f $X=1.75 $Y=1.035 $X2=0 $Y2=0
cc_140 N_TE_c_154_n N_A_27_47#_c_290_n 0.014005f $X=2.17 $Y=1.035 $X2=0 $Y2=0
cc_141 N_TE_c_155_n N_A_27_47#_c_291_n 0.014005f $X=2.59 $Y=1.035 $X2=0 $Y2=0
cc_142 N_TE_c_156_n N_A_27_47#_c_292_n 0.014005f $X=3.01 $Y=1.035 $X2=0 $Y2=0
cc_143 N_TE_c_157_n N_A_27_47#_c_293_n 0.014005f $X=3.43 $Y=1.035 $X2=0 $Y2=0
cc_144 N_TE_c_133_n N_A_27_47#_c_270_n 0.0150211f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_145 N_TE_c_134_n N_A_27_47#_c_270_n 3.34655e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_146 N_TE_c_135_n N_A_27_47#_c_270_n 0.00303485f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_147 N_TE_c_136_n N_A_27_47#_c_270_n 0.00161437f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_148 TE N_A_27_47#_c_270_n 0.019129f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_149 N_TE_c_133_n N_A_27_47#_c_271_n 0.00680774f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_150 N_TE_c_134_n N_A_27_47#_c_271_n 0.00300693f $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_151 N_TE_c_135_n N_A_27_47#_c_271_n 0.0014487f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_152 N_TE_c_136_n N_A_27_47#_c_271_n 0.00302911f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_153 N_TE_M1023_g N_A_27_47#_c_296_n 0.0379477f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_154 N_TE_c_134_n N_A_27_47#_c_296_n 5.69379e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_155 N_TE_c_135_n N_A_27_47#_c_296_n 0.00191321f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_156 TE N_A_27_47#_c_296_n 0.0421802f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_157 N_TE_c_137_n N_A_27_47#_c_272_n 0.0139399f $X=1.255 $Y=1.035 $X2=0 $Y2=0
cc_158 N_TE_c_139_n N_A_27_47#_c_272_n 0.0083577f $X=1.675 $Y=1.035 $X2=0 $Y2=0
cc_159 N_TE_c_141_n N_A_27_47#_c_272_n 0.008352f $X=2.095 $Y=1.035 $X2=0 $Y2=0
cc_160 N_TE_c_143_n N_A_27_47#_c_272_n 0.0083577f $X=2.515 $Y=1.035 $X2=0 $Y2=0
cc_161 N_TE_c_145_n N_A_27_47#_c_272_n 0.008352f $X=2.935 $Y=1.035 $X2=0 $Y2=0
cc_162 N_TE_c_147_n N_A_27_47#_c_272_n 0.0083577f $X=3.355 $Y=1.035 $X2=0 $Y2=0
cc_163 N_TE_c_149_n N_A_27_47#_c_272_n 0.0145953f $X=3.775 $Y=1.035 $X2=0 $Y2=0
cc_164 N_TE_c_151_n N_A_27_47#_c_272_n 0.00686545f $X=0.89 $Y=1.035 $X2=0 $Y2=0
cc_165 N_TE_c_152_n N_A_27_47#_c_272_n 0.0058582f $X=1.33 $Y=1.035 $X2=0 $Y2=0
cc_166 N_TE_c_153_n N_A_27_47#_c_272_n 0.0051004f $X=1.75 $Y=1.035 $X2=0 $Y2=0
cc_167 N_TE_c_154_n N_A_27_47#_c_272_n 0.0051004f $X=2.17 $Y=1.035 $X2=0 $Y2=0
cc_168 N_TE_c_155_n N_A_27_47#_c_272_n 0.0051004f $X=2.59 $Y=1.035 $X2=0 $Y2=0
cc_169 N_TE_c_156_n N_A_27_47#_c_272_n 0.0051004f $X=3.01 $Y=1.035 $X2=0 $Y2=0
cc_170 N_TE_c_157_n N_A_27_47#_c_272_n 0.0051004f $X=3.43 $Y=1.035 $X2=0 $Y2=0
cc_171 N_TE_c_149_n N_A_27_47#_c_273_n 0.00670028f $X=3.775 $Y=1.035 $X2=0 $Y2=0
cc_172 N_TE_c_134_n N_A_27_47#_c_340_n 0.0120485f $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_173 N_TE_c_135_n N_A_27_47#_c_340_n 0.0115132f $X=0.545 $Y=1.035 $X2=0 $Y2=0
cc_174 N_TE_c_151_n N_A_27_47#_c_340_n 0.00442816f $X=0.89 $Y=1.035 $X2=0 $Y2=0
cc_175 TE N_A_27_47#_c_340_n 0.025787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_176 N_TE_M1023_g N_VPWR_c_566_n 0.0113741f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_177 N_TE_M1023_g N_VPWR_c_575_n 0.0046653f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_178 N_TE_M1023_g N_VPWR_c_565_n 0.00523707f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_179 N_TE_M1023_g N_A_215_309#_c_689_n 0.00545173f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_TE_M1023_g N_A_215_309#_c_686_n 6.87579e-19 $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_181 N_TE_c_137_n N_A_215_309#_c_686_n 0.00101624f $X=1.255 $Y=1.035 $X2=0
+ $Y2=0
cc_182 N_TE_c_141_n N_A_215_309#_c_692_n 2.11158e-19 $X=2.095 $Y=1.035 $X2=0
+ $Y2=0
cc_183 N_TE_c_145_n N_A_215_309#_c_693_n 2.11158e-19 $X=2.935 $Y=1.035 $X2=0
+ $Y2=0
cc_184 N_TE_c_149_n N_A_215_309#_c_694_n 2.11158e-19 $X=3.775 $Y=1.035 $X2=0
+ $Y2=0
cc_185 N_TE_c_133_n N_VGND_c_885_n 0.00856801f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_186 N_TE_c_134_n N_VGND_c_885_n 5.1499e-19 $X=0.815 $Y=1.035 $X2=0 $Y2=0
cc_187 N_TE_c_136_n N_VGND_c_885_n 0.00735324f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_188 N_TE_c_138_n N_VGND_c_885_n 5.57248e-19 $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_189 N_TE_c_136_n N_VGND_c_886_n 5.5023e-19 $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_190 N_TE_c_138_n N_VGND_c_886_n 0.00691072f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_191 N_TE_c_140_n N_VGND_c_886_n 0.00685342f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_192 N_TE_c_142_n N_VGND_c_886_n 5.54209e-19 $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_193 N_TE_c_140_n N_VGND_c_887_n 5.54209e-19 $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_194 N_TE_c_142_n N_VGND_c_887_n 0.00685342f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_195 N_TE_c_144_n N_VGND_c_887_n 0.00685342f $X=2.59 $Y=0.96 $X2=0 $Y2=0
cc_196 N_TE_c_146_n N_VGND_c_887_n 5.54209e-19 $X=3.01 $Y=0.96 $X2=0 $Y2=0
cc_197 N_TE_c_144_n N_VGND_c_888_n 5.54209e-19 $X=2.59 $Y=0.96 $X2=0 $Y2=0
cc_198 N_TE_c_146_n N_VGND_c_888_n 0.00685342f $X=3.01 $Y=0.96 $X2=0 $Y2=0
cc_199 N_TE_c_148_n N_VGND_c_888_n 0.00685342f $X=3.43 $Y=0.96 $X2=0 $Y2=0
cc_200 N_TE_c_150_n N_VGND_c_888_n 5.54209e-19 $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_201 N_TE_c_148_n N_VGND_c_889_n 0.00341689f $X=3.43 $Y=0.96 $X2=0 $Y2=0
cc_202 N_TE_c_150_n N_VGND_c_889_n 0.00341689f $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_203 N_TE_c_148_n N_VGND_c_890_n 5.54817e-19 $X=3.43 $Y=0.96 $X2=0 $Y2=0
cc_204 N_TE_c_150_n N_VGND_c_890_n 0.0079747f $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_205 N_TE_c_140_n N_VGND_c_891_n 0.00341689f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_206 N_TE_c_142_n N_VGND_c_891_n 0.00341689f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_207 N_TE_c_144_n N_VGND_c_893_n 0.00341689f $X=2.59 $Y=0.96 $X2=0 $Y2=0
cc_208 N_TE_c_146_n N_VGND_c_893_n 0.00341689f $X=3.01 $Y=0.96 $X2=0 $Y2=0
cc_209 N_TE_c_133_n N_VGND_c_895_n 0.00341689f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_210 N_TE_c_136_n N_VGND_c_896_n 0.0046653f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_211 N_TE_c_138_n N_VGND_c_896_n 0.00341689f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_212 N_TE_c_133_n N_VGND_c_898_n 0.0050171f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_213 N_TE_c_136_n N_VGND_c_898_n 0.00802193f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_214 N_TE_c_138_n N_VGND_c_898_n 0.00408046f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_215 N_TE_c_140_n N_VGND_c_898_n 0.0040262f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_216 N_TE_c_142_n N_VGND_c_898_n 0.0040262f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_217 N_TE_c_144_n N_VGND_c_898_n 0.0040262f $X=2.59 $Y=0.96 $X2=0 $Y2=0
cc_218 N_TE_c_146_n N_VGND_c_898_n 0.0040262f $X=3.01 $Y=0.96 $X2=0 $Y2=0
cc_219 N_TE_c_148_n N_VGND_c_898_n 0.0040262f $X=3.43 $Y=0.96 $X2=0 $Y2=0
cc_220 N_TE_c_150_n N_VGND_c_898_n 0.0040262f $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_221 N_TE_c_136_n N_A_193_47#_c_1016_n 0.0043107f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_222 N_TE_c_138_n N_A_193_47#_c_1017_n 0.0103667f $X=1.33 $Y=0.96 $X2=0 $Y2=0
cc_223 N_TE_c_139_n N_A_193_47#_c_1017_n 0.00179137f $X=1.675 $Y=1.035 $X2=0
+ $Y2=0
cc_224 N_TE_c_140_n N_A_193_47#_c_1017_n 0.0104925f $X=1.75 $Y=0.96 $X2=0 $Y2=0
cc_225 N_TE_c_136_n N_A_193_47#_c_1020_n 0.00161811f $X=0.89 $Y=0.96 $X2=0 $Y2=0
cc_226 N_TE_c_137_n N_A_193_47#_c_1020_n 0.00227361f $X=1.255 $Y=1.035 $X2=0
+ $Y2=0
cc_227 N_TE_c_142_n N_A_193_47#_c_1022_n 0.0105367f $X=2.17 $Y=0.96 $X2=0 $Y2=0
cc_228 N_TE_c_143_n N_A_193_47#_c_1022_n 0.00179137f $X=2.515 $Y=1.035 $X2=0
+ $Y2=0
cc_229 N_TE_c_144_n N_A_193_47#_c_1022_n 0.0105367f $X=2.59 $Y=0.96 $X2=0 $Y2=0
cc_230 N_TE_c_146_n N_A_193_47#_c_1025_n 0.0105367f $X=3.01 $Y=0.96 $X2=0 $Y2=0
cc_231 N_TE_c_147_n N_A_193_47#_c_1025_n 0.00179137f $X=3.355 $Y=1.035 $X2=0
+ $Y2=0
cc_232 N_TE_c_148_n N_A_193_47#_c_1025_n 0.0105367f $X=3.43 $Y=0.96 $X2=0 $Y2=0
cc_233 N_TE_c_150_n N_A_193_47#_c_1012_n 0.0126397f $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_234 N_TE_c_150_n N_A_193_47#_c_1013_n 0.00362209f $X=3.85 $Y=0.96 $X2=0 $Y2=0
cc_235 N_TE_c_141_n N_A_193_47#_c_1030_n 0.00186022f $X=2.095 $Y=1.035 $X2=0
+ $Y2=0
cc_236 N_TE_c_145_n N_A_193_47#_c_1031_n 0.00186022f $X=2.935 $Y=1.035 $X2=0
+ $Y2=0
cc_237 N_TE_c_149_n N_A_193_47#_c_1032_n 0.00186022f $X=3.775 $Y=1.035 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_c_294_n N_A_M1002_g 0.0169129f $X=4.35 $Y=1.395 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_272_n N_A_c_442_n 0.00353496f $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_273_n N_A_c_442_n 0.0169129f $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_296_n N_VPWR_M1023_d 0.00535662f $X=0.687 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_242 N_A_27_47#_c_274_n N_VPWR_c_566_n 0.00230982f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_296_n N_VPWR_c_566_n 0.0238531f $X=0.687 $Y=1.785 $X2=0
+ $Y2=0
cc_244 N_A_27_47#_c_274_n N_VPWR_c_567_n 0.0109235f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_277_n N_VPWR_c_567_n 0.0104025f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_279_n N_VPWR_c_567_n 6.14905e-19 $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_277_n N_VPWR_c_568_n 6.14905e-19 $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_279_n N_VPWR_c_568_n 0.0104025f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_281_n N_VPWR_c_568_n 0.0104025f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_283_n N_VPWR_c_568_n 6.14905e-19 $X=3.09 $Y=1.47 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_281_n N_VPWR_c_569_n 6.14905e-19 $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_283_n N_VPWR_c_569_n 0.0104025f $X=3.09 $Y=1.47 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_285_n N_VPWR_c_569_n 0.0104025f $X=3.51 $Y=1.47 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_287_n N_VPWR_c_569_n 6.14905e-19 $X=3.93 $Y=1.47 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_285_n N_VPWR_c_570_n 6.14905e-19 $X=3.51 $Y=1.47 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_287_n N_VPWR_c_570_n 0.0104025f $X=3.93 $Y=1.47 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_288_n N_VPWR_c_570_n 0.0116531f $X=4.35 $Y=1.47 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_281_n N_VPWR_c_571_n 0.0046653f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_283_n N_VPWR_c_571_n 0.0046653f $X=3.09 $Y=1.47 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_285_n N_VPWR_c_573_n 0.0046653f $X=3.51 $Y=1.47 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_287_n N_VPWR_c_573_n 0.0046653f $X=3.93 $Y=1.47 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_295_n N_VPWR_c_575_n 0.0176305f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_274_n N_VPWR_c_576_n 0.0046653f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_277_n N_VPWR_c_577_n 0.0046653f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_279_n N_VPWR_c_577_n 0.0046653f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_288_n N_VPWR_c_578_n 0.0046653f $X=4.35 $Y=1.47 $X2=0 $Y2=0
cc_267 N_A_27_47#_M1023_s N_VPWR_c_565_n 0.00238524f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_274_n N_VPWR_c_565_n 0.00934473f $X=1.41 $Y=1.47 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_277_n N_VPWR_c_565_n 0.00789179f $X=1.83 $Y=1.47 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_279_n N_VPWR_c_565_n 0.00789179f $X=2.25 $Y=1.47 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_281_n N_VPWR_c_565_n 0.00789179f $X=2.67 $Y=1.47 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_283_n N_VPWR_c_565_n 0.00789179f $X=3.09 $Y=1.47 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_285_n N_VPWR_c_565_n 0.00789179f $X=3.51 $Y=1.47 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_287_n N_VPWR_c_565_n 0.00789179f $X=3.93 $Y=1.47 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_288_n N_VPWR_c_565_n 0.00804845f $X=4.35 $Y=1.47 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_295_n N_VPWR_c_565_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_296_n N_VPWR_c_565_n 0.00671954f $X=0.687 $Y=1.785 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_296_n N_A_215_309#_c_689_n 0.0168242f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_279 N_A_27_47#_c_274_n N_A_215_309#_c_696_n 0.0155912f $X=1.41 $Y=1.47 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_275_n N_A_215_309#_c_696_n 0.00197697f $X=1.755 $Y=1.395
+ $X2=0 $Y2=0
cc_281 N_A_27_47#_c_277_n N_A_215_309#_c_696_n 0.0142192f $X=1.83 $Y=1.47 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_272_n N_A_215_309#_c_696_n 0.0323847f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_296_n N_A_215_309#_c_686_n 0.0132199f $X=0.687 $Y=1.785
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_272_n N_A_215_309#_c_686_n 0.0143803f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_279_n N_A_215_309#_c_702_n 0.0142634f $X=2.25 $Y=1.47 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_280_n N_A_215_309#_c_702_n 0.00197697f $X=2.595 $Y=1.395
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_281_n N_A_215_309#_c_702_n 0.0142634f $X=2.67 $Y=1.47 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_272_n N_A_215_309#_c_702_n 0.0321432f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_283_n N_A_215_309#_c_706_n 0.0142634f $X=3.09 $Y=1.47 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_284_n N_A_215_309#_c_706_n 0.00197697f $X=3.435 $Y=1.395
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_285_n N_A_215_309#_c_706_n 0.0142634f $X=3.51 $Y=1.47 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_272_n N_A_215_309#_c_706_n 0.0321432f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_287_n N_A_215_309#_c_710_n 0.0143019f $X=3.93 $Y=1.47 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_288_n N_A_215_309#_c_710_n 0.0143232f $X=4.35 $Y=1.47 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_294_n N_A_215_309#_c_710_n 0.0021442f $X=4.35 $Y=1.395 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_272_n N_A_215_309#_c_710_n 0.0476181f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_278_n N_A_215_309#_c_692_n 0.00209962f $X=2.175 $Y=1.395
+ $X2=0 $Y2=0
cc_298 N_A_27_47#_c_272_n N_A_215_309#_c_692_n 0.0106208f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_282_n N_A_215_309#_c_693_n 0.00209962f $X=3.015 $Y=1.395
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_272_n N_A_215_309#_c_693_n 0.0106208f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_286_n N_A_215_309#_c_694_n 0.00209962f $X=3.855 $Y=1.395
+ $X2=0 $Y2=0
cc_302 N_A_27_47#_c_272_n N_A_215_309#_c_694_n 0.0106208f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_294_n Z 0.00124898f $X=4.35 $Y=1.395 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_272_n Z 0.027927f $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_273_n Z 2.33571e-19 $X=4.29 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_270_n N_VGND_M1030_d 0.00310523f $X=0.597 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_307 N_A_27_47#_c_271_n N_VGND_M1030_d 9.5711e-19 $X=0.597 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_308 N_A_27_47#_c_270_n N_VGND_c_885_n 0.00918217f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_340_n N_VGND_c_885_n 0.004225f $X=0.687 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_269_n N_VGND_c_895_n 0.0173297f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_270_n N_VGND_c_895_n 0.00235711f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_M1030_s N_VGND_c_898_n 0.00230206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_269_n N_VGND_c_898_n 0.00980382f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_270_n N_VGND_c_898_n 0.00499131f $X=0.597 $Y=0.825 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_272_n N_A_193_47#_c_1017_n 0.0408222f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_c_270_n N_A_193_47#_c_1020_n 0.00897896f $X=0.597 $Y=0.825
+ $X2=0 $Y2=0
cc_317 N_A_27_47#_c_272_n N_A_193_47#_c_1020_n 0.0135368f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_272_n N_A_193_47#_c_1022_n 0.0408222f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_272_n N_A_193_47#_c_1025_n 0.0408222f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_294_n N_A_193_47#_c_1012_n 7.32088e-19 $X=4.35 $Y=1.395
+ $X2=0 $Y2=0
cc_321 N_A_27_47#_c_272_n N_A_193_47#_c_1012_n 0.0720833f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_273_n N_A_193_47#_c_1012_n 0.00706393f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_272_n N_A_193_47#_c_1030_n 0.0132296f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_272_n N_A_193_47#_c_1031_n 0.0132296f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_272_n N_A_193_47#_c_1032_n 0.0132296f $X=4.29 $Y=1.16 $X2=0
+ $Y2=0
cc_326 N_A_M1002_g N_VPWR_c_570_n 0.00102044f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A_M1002_g N_VPWR_c_578_n 0.00357877f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_M1007_g N_VPWR_c_578_n 0.00357877f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_M1017_g N_VPWR_c_578_n 0.00357877f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_M1018_g N_VPWR_c_578_n 0.00357877f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_331 N_A_M1022_g N_VPWR_c_578_n 0.00357877f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_332 N_A_M1025_g N_VPWR_c_578_n 0.00357877f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_333 N_A_M1026_g N_VPWR_c_578_n 0.00357877f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A_M1029_g N_VPWR_c_578_n 0.00357877f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_M1002_g N_VPWR_c_565_n 0.00538183f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_M1007_g N_VPWR_c_565_n 0.00522516f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_M1017_g N_VPWR_c_565_n 0.00522516f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_338 N_A_M1018_g N_VPWR_c_565_n 0.00522516f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_M1022_g N_VPWR_c_565_n 0.00522516f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_340 N_A_M1025_g N_VPWR_c_565_n 0.00522516f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_341 N_A_M1026_g N_VPWR_c_565_n 0.00522516f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_342 N_A_M1029_g N_VPWR_c_565_n 0.00621986f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_343 N_A_M1002_g N_A_215_309#_c_720_n 0.0112878f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_M1007_g N_A_215_309#_c_720_n 0.0112437f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_345 N_A_M1017_g N_A_215_309#_c_722_n 0.0112585f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_346 N_A_M1018_g N_A_215_309#_c_722_n 0.0112585f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_347 N_A_M1022_g N_A_215_309#_c_724_n 0.0112878f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A_M1025_g N_A_215_309#_c_724_n 0.0112878f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_349 N_A_M1026_g N_A_215_309#_c_687_n 0.0112878f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_350 N_A_M1029_g N_A_215_309#_c_687_n 0.0112878f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_351 N_A_c_442_n N_A_215_309#_c_688_n 0.00562759f $X=7.765 $Y=1.015 $X2=0
+ $Y2=0
cc_352 N_A_M1029_g N_A_215_309#_c_688_n 0.00628807f $X=7.765 $Y=1.985 $X2=0
+ $Y2=0
cc_353 A N_A_215_309#_c_688_n 0.0253648f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_354 N_A_c_433_n N_Z_c_788_n 0.00662588f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A_M1006_g N_Z_c_788_n 0.00955084f $X=5.665 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_M1011_g N_Z_c_788_n 0.00955084f $X=6.085 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_c_438_n N_Z_c_788_n 0.00955084f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A_c_439_n N_Z_c_788_n 0.00955084f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A_M1032_g N_Z_c_788_n 0.00955084f $X=7.345 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_c_442_n N_Z_c_788_n 0.0117461f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_361 N_A_M1033_g N_Z_c_788_n 0.0115423f $X=7.765 $Y=0.56 $X2=0 $Y2=0
cc_362 A N_Z_c_788_n 0.181633f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_363 N_A_c_432_n N_Z_c_807_n 0.00369523f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_c_433_n N_Z_c_807_n 0.00273142f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A_c_432_n Z 0.00761361f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A_M1002_g Z 0.012805f $X=4.825 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_c_433_n Z 0.00447935f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A_M1007_g Z 0.0151729f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_369 N_A_M1006_g Z 9.23891e-19 $X=5.665 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_M1017_g Z 0.00136258f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A_c_442_n Z 0.0238164f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_372 A Z 0.0204219f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_373 N_A_M1017_g Z 0.00142036f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A_M1018_g Z 0.00142036f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_375 N_A_c_442_n Z 0.0019843f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_376 A Z 0.0242306f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_377 N_A_M1022_g Z 0.0013397f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_378 N_A_M1025_g Z 0.0013397f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_379 N_A_c_442_n Z 0.00222344f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_380 A Z 0.0270806f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_381 N_A_M1018_g Z 5.55259e-19 $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_382 N_A_M1022_g Z 0.00687627f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_383 N_A_M1025_g Z 0.00688691f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_384 N_A_M1026_g Z 5.55478e-19 $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_385 N_A_M1026_g Z 0.0013397f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_386 N_A_c_442_n Z 0.00206069f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_387 N_A_M1029_g Z 0.00275184f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_388 A Z 0.0270809f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_389 N_A_M1025_g Z 5.55478e-19 $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_390 N_A_M1026_g Z 0.00688691f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_391 N_A_M1029_g Z 0.00599632f $X=7.765 $Y=1.985 $X2=0 $Y2=0
cc_392 N_A_M1007_g N_Z_c_792_n 0.00792131f $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_393 N_A_M1017_g N_Z_c_792_n 0.0107189f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_394 N_A_c_442_n N_Z_c_792_n 0.00202711f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_395 A N_Z_c_792_n 0.020892f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_396 N_A_M1018_g N_Z_c_793_n 0.0107189f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_397 N_A_M1022_g N_Z_c_793_n 0.0107189f $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_398 N_A_c_442_n N_Z_c_793_n 0.00198252f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_399 A N_Z_c_793_n 0.036625f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_400 N_A_M1025_g N_Z_c_794_n 0.0107189f $X=6.925 $Y=1.985 $X2=0 $Y2=0
cc_401 N_A_M1026_g N_Z_c_794_n 0.0107189f $X=7.345 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A_c_442_n N_Z_c_794_n 0.00198252f $X=7.765 $Y=1.015 $X2=0 $Y2=0
cc_403 A N_Z_c_794_n 0.036625f $X=7.99 $Y=1.105 $X2=0 $Y2=0
cc_404 N_A_M1007_g N_Z_c_848_n 5.53432e-19 $X=5.245 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A_M1017_g N_Z_c_848_n 0.00700222f $X=5.665 $Y=1.985 $X2=0 $Y2=0
cc_406 N_A_M1018_g N_Z_c_848_n 0.00700222f $X=6.085 $Y=1.985 $X2=0 $Y2=0
cc_407 N_A_M1022_g N_Z_c_848_n 5.53432e-19 $X=6.505 $Y=1.985 $X2=0 $Y2=0
cc_408 N_A_c_432_n N_VGND_c_890_n 0.00295671f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A_c_432_n N_VGND_c_897_n 0.00357877f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A_c_433_n N_VGND_c_897_n 0.00357877f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A_M1006_g N_VGND_c_897_n 0.00357877f $X=5.665 $Y=0.56 $X2=0 $Y2=0
cc_412 N_A_M1011_g N_VGND_c_897_n 0.00357877f $X=6.085 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A_c_438_n N_VGND_c_897_n 0.00357877f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A_c_439_n N_VGND_c_897_n 0.00357877f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A_M1032_g N_VGND_c_897_n 0.00357877f $X=7.345 $Y=0.56 $X2=0 $Y2=0
cc_416 N_A_M1033_g N_VGND_c_897_n 0.00357877f $X=7.765 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A_c_432_n N_VGND_c_898_n 0.00664112f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_418 N_A_c_433_n N_VGND_c_898_n 0.00522516f $X=5.245 $Y=0.995 $X2=0 $Y2=0
cc_419 N_A_M1006_g N_VGND_c_898_n 0.00522516f $X=5.665 $Y=0.56 $X2=0 $Y2=0
cc_420 N_A_M1011_g N_VGND_c_898_n 0.00522516f $X=6.085 $Y=0.56 $X2=0 $Y2=0
cc_421 N_A_c_438_n N_VGND_c_898_n 0.00522516f $X=6.505 $Y=0.995 $X2=0 $Y2=0
cc_422 N_A_c_439_n N_VGND_c_898_n 0.00522516f $X=6.925 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A_M1032_g N_VGND_c_898_n 0.00522516f $X=7.345 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A_M1033_g N_VGND_c_898_n 0.00621986f $X=7.765 $Y=0.56 $X2=0 $Y2=0
cc_425 N_A_c_432_n N_A_193_47#_c_1015_n 0.014178f $X=4.825 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A_c_433_n N_A_193_47#_c_1015_n 0.00866372f $X=5.245 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_A_M1006_g N_A_193_47#_c_1015_n 0.00866705f $X=5.665 $Y=0.56 $X2=0 $Y2=0
cc_428 N_A_M1011_g N_A_193_47#_c_1015_n 0.00866705f $X=6.085 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A_c_438_n N_A_193_47#_c_1015_n 0.00866705f $X=6.505 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_c_439_n N_A_193_47#_c_1015_n 0.00866705f $X=6.925 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A_M1032_g N_A_193_47#_c_1015_n 0.00866705f $X=7.345 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A_c_442_n N_A_193_47#_c_1015_n 3.01257e-19 $X=7.765 $Y=1.015 $X2=0
+ $Y2=0
cc_433 N_A_M1033_g N_A_193_47#_c_1015_n 0.00866705f $X=7.765 $Y=0.56 $X2=0 $Y2=0
cc_434 N_VPWR_c_565_n N_A_215_309#_M1000_d 0.00386369f $X=8.05 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_435 N_VPWR_c_565_n N_A_215_309#_M1001_d 0.00562358f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_565_n N_A_215_309#_M1008_d 0.00562358f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_565_n N_A_215_309#_M1013_d 0.00562358f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_565_n N_A_215_309#_M1027_d 0.00429477f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_565_n N_A_215_309#_M1007_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_565_n N_A_215_309#_M1018_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_565_n N_A_215_309#_M1025_s 0.0021521f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_565_n N_A_215_309#_M1029_s 0.00209324f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_566_n N_A_215_309#_c_689_n 0.0240954f $X=0.68 $Y=2.34 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_576_n N_A_215_309#_c_689_n 0.0144177f $X=1.455 $Y=2.72 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_565_n N_A_215_309#_c_689_n 0.00801045f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_446 N_VPWR_M1000_s N_A_215_309#_c_696_n 0.00318028f $X=1.485 $Y=1.545 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_567_n N_A_215_309#_c_696_n 0.0170258f $X=1.62 $Y=2.02 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_577_n N_A_215_309#_c_745_n 0.0113958f $X=2.295 $Y=2.72 $X2=0
+ $Y2=0
cc_449 N_VPWR_c_565_n N_A_215_309#_c_745_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_450 N_VPWR_M1005_s N_A_215_309#_c_702_n 0.00318028f $X=2.325 $Y=1.545 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_568_n N_A_215_309#_c_702_n 0.0170258f $X=2.46 $Y=2.02 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_571_n N_A_215_309#_c_749_n 0.0113958f $X=3.135 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_565_n N_A_215_309#_c_749_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_M1009_s N_A_215_309#_c_706_n 0.00318028f $X=3.165 $Y=1.545 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_569_n N_A_215_309#_c_706_n 0.0170258f $X=3.3 $Y=2.02 $X2=0 $Y2=0
cc_456 N_VPWR_c_573_n N_A_215_309#_c_753_n 0.0113958f $X=3.975 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_565_n N_A_215_309#_c_753_n 0.00646998f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_M1024_s N_A_215_309#_c_710_n 0.00328966f $X=4.005 $Y=1.545 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_570_n N_A_215_309#_c_710_n 0.0170258f $X=4.14 $Y=2.02 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_578_n N_A_215_309#_c_720_n 0.0358391f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_565_n N_A_215_309#_c_720_n 0.0234424f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_578_n N_A_215_309#_c_759_n 0.0153344f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_565_n N_A_215_309#_c_759_n 0.00866514f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_578_n N_A_215_309#_c_722_n 0.0358391f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_565_n N_A_215_309#_c_722_n 0.0234424f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_578_n N_A_215_309#_c_724_n 0.0358391f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_565_n N_A_215_309#_c_724_n 0.0234424f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_578_n N_A_215_309#_c_687_n 0.0571736f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_565_n N_A_215_309#_c_687_n 0.0351832f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_578_n N_A_215_309#_c_767_n 0.0114668f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_565_n N_A_215_309#_c_767_n 0.006547f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_472 N_VPWR_c_578_n N_A_215_309#_c_769_n 0.0114668f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_565_n N_A_215_309#_c_769_n 0.006547f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_474 N_VPWR_c_578_n N_A_215_309#_c_771_n 0.0114668f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_565_n N_A_215_309#_c_771_n 0.006547f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_476 N_VPWR_c_565_n N_Z_M1002_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_477 N_VPWR_c_565_n N_Z_M1017_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_478 N_VPWR_c_565_n N_Z_M1022_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_479 N_VPWR_c_565_n N_Z_M1026_d 0.00216833f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_480 N_A_215_309#_c_720_n N_Z_M1002_d 0.00312348f $X=5.37 $Y=2.38 $X2=0 $Y2=0
cc_481 N_A_215_309#_c_722_n N_Z_M1017_d 0.00312752f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_482 N_A_215_309#_c_724_n N_Z_M1022_d 0.00312348f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_483 N_A_215_309#_c_687_n N_Z_M1026_d 0.00312348f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_484 N_A_215_309#_c_720_n Z 0.015949f $X=5.37 $Y=2.38 $X2=0 $Y2=0
cc_485 N_A_215_309#_c_724_n Z 0.015949f $X=7.05 $Y=2.38 $X2=0 $Y2=0
cc_486 N_A_215_309#_c_688_n Z 0.00877121f $X=8.042 $Y=2.295 $X2=0 $Y2=0
cc_487 N_A_215_309#_c_687_n Z 0.015949f $X=7.89 $Y=2.38 $X2=0 $Y2=0
cc_488 N_A_215_309#_M1007_s N_Z_c_792_n 0.00165831f $X=5.32 $Y=1.485 $X2=0 $Y2=0
cc_489 N_A_215_309#_c_782_p N_Z_c_792_n 0.0126919f $X=5.455 $Y=1.96 $X2=0 $Y2=0
cc_490 N_A_215_309#_M1018_s N_Z_c_793_n 0.00165831f $X=6.16 $Y=1.485 $X2=0 $Y2=0
cc_491 N_A_215_309#_c_784_p N_Z_c_793_n 0.0126919f $X=6.295 $Y=1.96 $X2=0 $Y2=0
cc_492 N_A_215_309#_M1025_s N_Z_c_794_n 0.00165831f $X=7 $Y=1.485 $X2=0 $Y2=0
cc_493 N_A_215_309#_c_786_p N_Z_c_794_n 0.0126919f $X=7.135 $Y=1.96 $X2=0 $Y2=0
cc_494 N_A_215_309#_c_722_n N_Z_c_848_n 0.0156554f $X=6.21 $Y=2.38 $X2=0 $Y2=0
cc_495 N_Z_M1003_s N_VGND_c_898_n 0.00216833f $X=4.9 $Y=0.235 $X2=0 $Y2=0
cc_496 N_Z_M1006_s N_VGND_c_898_n 0.00216833f $X=5.74 $Y=0.235 $X2=0 $Y2=0
cc_497 N_Z_M1028_s N_VGND_c_898_n 0.00216833f $X=6.58 $Y=0.235 $X2=0 $Y2=0
cc_498 N_Z_M1032_s N_VGND_c_898_n 0.00216833f $X=7.42 $Y=0.235 $X2=0 $Y2=0
cc_499 N_Z_c_788_n N_A_193_47#_M1004_d 0.00338736f $X=7.555 $Y=0.76 $X2=0 $Y2=0
cc_500 N_Z_c_788_n N_A_193_47#_M1011_d 0.00307913f $X=7.555 $Y=0.76 $X2=0 $Y2=0
cc_501 N_Z_c_788_n N_A_193_47#_M1031_d 0.00307913f $X=7.555 $Y=0.76 $X2=0 $Y2=0
cc_502 N_Z_c_788_n N_A_193_47#_M1033_d 0.00531396f $X=7.555 $Y=0.76 $X2=0 $Y2=0
cc_503 N_Z_M1003_s N_A_193_47#_c_1015_n 0.00304479f $X=4.9 $Y=0.235 $X2=0 $Y2=0
cc_504 N_Z_M1006_s N_A_193_47#_c_1015_n 0.00305599f $X=5.74 $Y=0.235 $X2=0 $Y2=0
cc_505 N_Z_M1028_s N_A_193_47#_c_1015_n 0.00304849f $X=6.58 $Y=0.235 $X2=0 $Y2=0
cc_506 N_Z_M1032_s N_A_193_47#_c_1015_n 0.00305599f $X=7.42 $Y=0.235 $X2=0 $Y2=0
cc_507 N_Z_c_788_n N_A_193_47#_c_1015_n 0.152241f $X=7.555 $Y=0.76 $X2=0 $Y2=0
cc_508 N_Z_c_807_n N_A_193_47#_c_1015_n 0.0201274f $X=5.06 $Y=0.85 $X2=0 $Y2=0
cc_509 N_VGND_c_898_n N_A_193_47#_M1010_s 0.00498236f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_510 N_VGND_c_898_n N_A_193_47#_M1014_s 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_898_n N_A_193_47#_M1016_s 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_898_n N_A_193_47#_M1020_s 0.00254582f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_898_n N_A_193_47#_M1003_d 0.00210127f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_898_n N_A_193_47#_M1004_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_898_n N_A_193_47#_M1011_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_898_n N_A_193_47#_M1031_d 0.00215227f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_898_n N_A_193_47#_M1033_d 0.00225742f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_885_n N_A_193_47#_c_1016_n 0.0155846f $X=0.68 $Y=0.36 $X2=0
+ $Y2=0
cc_519 N_VGND_c_896_n N_A_193_47#_c_1016_n 0.011459f $X=1.375 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_898_n N_A_193_47#_c_1016_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_M1012_d N_A_193_47#_c_1017_n 0.00297022f $X=1.405 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_VGND_c_886_n N_A_193_47#_c_1017_n 0.0160613f $X=1.54 $Y=0.36 $X2=0
+ $Y2=0
cc_523 N_VGND_c_891_n N_A_193_47#_c_1017_n 0.00232396f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_896_n N_A_193_47#_c_1017_n 0.00232396f $X=1.375 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_898_n N_A_193_47#_c_1017_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_891_n N_A_193_47#_c_1080_n 0.0112554f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_898_n N_A_193_47#_c_1080_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_M1015_d N_A_193_47#_c_1022_n 0.00297022f $X=2.245 $Y=0.235 $X2=0
+ $Y2=0
cc_529 N_VGND_c_887_n N_A_193_47#_c_1022_n 0.0160613f $X=2.38 $Y=0.36 $X2=0
+ $Y2=0
cc_530 N_VGND_c_891_n N_A_193_47#_c_1022_n 0.00232396f $X=2.215 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_893_n N_A_193_47#_c_1022_n 0.00232396f $X=3.055 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_898_n N_A_193_47#_c_1022_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_893_n N_A_193_47#_c_1087_n 0.0112554f $X=3.055 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_898_n N_A_193_47#_c_1087_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_535 N_VGND_M1019_d N_A_193_47#_c_1025_n 0.00297022f $X=3.085 $Y=0.235 $X2=0
+ $Y2=0
cc_536 N_VGND_c_888_n N_A_193_47#_c_1025_n 0.0160613f $X=3.22 $Y=0.36 $X2=0
+ $Y2=0
cc_537 N_VGND_c_889_n N_A_193_47#_c_1025_n 0.00232396f $X=3.895 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_893_n N_A_193_47#_c_1025_n 0.00232396f $X=3.055 $Y=0 $X2=0 $Y2=0
cc_539 N_VGND_c_898_n N_A_193_47#_c_1025_n 0.00970544f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_889_n N_A_193_47#_c_1094_n 0.0112554f $X=3.895 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_898_n N_A_193_47#_c_1094_n 0.00644035f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_542 N_VGND_M1021_d N_A_193_47#_c_1012_n 0.00522868f $X=3.925 $Y=0.235 $X2=0
+ $Y2=0
cc_543 N_VGND_c_889_n N_A_193_47#_c_1012_n 0.00232396f $X=3.895 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_890_n N_A_193_47#_c_1012_n 0.0214727f $X=4.06 $Y=0.36 $X2=0
+ $Y2=0
cc_545 N_VGND_c_897_n N_A_193_47#_c_1012_n 0.00296166f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_546 N_VGND_c_898_n N_A_193_47#_c_1012_n 0.0103752f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_547 N_VGND_c_890_n N_A_193_47#_c_1013_n 0.0016142f $X=4.06 $Y=0.36 $X2=0
+ $Y2=0
cc_548 N_VGND_c_890_n N_A_193_47#_c_1014_n 0.0186164f $X=4.06 $Y=0.36 $X2=0
+ $Y2=0
cc_549 N_VGND_c_897_n N_A_193_47#_c_1014_n 0.0203543f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_898_n N_A_193_47#_c_1014_n 0.011309f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_897_n N_A_193_47#_c_1015_n 0.196043f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_898_n N_A_193_47#_c_1015_n 0.124805f $X=8.05 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a22o_1.pex.spice
* Created: Thu Aug 27 14:02:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A22O_1%B2 3 6 8 11 12 13
r26 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=1.325
r27 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.41 $Y2=0.995
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r29 8 12 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.41 $Y2=1.175
r30 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.985
+ $X2=0.47 $Y2=1.325
r31 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%B1 3 6 8 9 13 15
c41 6 0 1.7212e-19 $X=0.89 $Y=1.985
r42 17 23 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=1.13 $Y=1.075
+ $X2=1.13 $Y2=1.18
r43 14 23 10.5628 $w=2.08e-07 $l=2e-07 $layer=LI1_cond $X=0.93 $Y=1.18 $X2=1.13
+ $Y2=1.18
r44 13 16 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=1.325
r45 13 15 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.92 $Y2=0.995
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.93
+ $Y=1.16 $X2=0.93 $Y2=1.16
r47 9 23 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.13 $Y2=1.18
r48 8 17 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.13 $Y=0.85
+ $X2=1.13 $Y2=1.075
r49 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.985
+ $X2=0.89 $Y2=1.325
r50 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.56 $X2=0.85
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%A1 1 3 4 6 7 8
c37 8 0 1.98592e-19 $X=1.61 $Y=1.19
r38 14 18 0.716491 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=1.59 $Y=1.075
+ $X2=1.59 $Y2=1.18
r39 8 18 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=1.18 $X2=1.59
+ $Y2=1.18
r40 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.16 $X2=1.65 $Y2=1.16
r41 7 14 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.59 $Y=0.85
+ $X2=1.59 $Y2=1.075
r42 4 12 50.3657 $w=3.56e-07 $l=3.06186e-07 $layer=POLY_cond $X=1.82 $Y=1.41
+ $X2=1.695 $Y2=1.16
r43 4 6 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.82 $Y=1.41 $X2=1.82
+ $Y2=1.985
r44 1 12 38.8573 $w=3.56e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.79 $Y=0.995
+ $X2=1.695 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.79 $Y=0.995 $X2=1.79
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%A2 1 3 4 6 8 12
c40 12 0 6.73606e-20 $X=2.23 $Y=1.16
c41 4 0 1.98592e-19 $X=2.29 $Y=1.325
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.16 $X2=2.23 $Y2=1.16
r43 8 12 6.0456 $w=3.03e-07 $l=1.6e-07 $layer=LI1_cond $X=2.07 $Y=1.192 $X2=2.23
+ $Y2=1.192
r44 4 11 38.7751 $w=2.77e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.29 $Y=1.325
+ $X2=2.225 $Y2=1.16
r45 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.29 $Y=1.325 $X2=2.29
+ $Y2=1.985
r46 1 11 44.8654 $w=2.77e-07 $l=2.30217e-07 $layer=POLY_cond $X=2.29 $Y=0.96
+ $X2=2.225 $Y2=1.16
r47 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.29 $Y=0.96 $X2=2.29
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%A_27_297# 1 2 3 4 15 18 23 25 26 32 35 36 37
+ 38 41 42 44 49 50 53
c107 42 0 1.55628e-19 $X=2.71 $Y=1.16
c108 18 0 6.73606e-20 $X=2.75 $Y=1.985
r109 48 50 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=1.585
+ $X2=1.265 $Y2=1.585
r110 48 49 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=1.585
+ $X2=0.935 $Y2=1.585
r111 44 45 3.9534 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=0.257 $Y=2.34
+ $X2=0.257 $Y2=2.245
r112 42 54 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.16
+ $X2=2.76 $Y2=1.325
r113 42 53 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.16
+ $X2=2.76 $Y2=0.995
r114 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.16 $X2=2.71 $Y2=1.16
r115 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.71 $Y=1.48
+ $X2=2.71 $Y2=1.16
r116 38 51 11.7016 $w=2.31e-07 $l=2.28637e-07 $layer=LI1_cond $X=2.71 $Y=0.905
+ $X2=2.66 $Y2=0.7
r117 38 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.71 $Y=0.905
+ $X2=2.71 $Y2=1.16
r118 36 51 2.5345 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=0.7
+ $X2=2.66 $Y2=0.7
r119 36 37 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.525 $Y=0.7
+ $X2=2.12 $Y2=0.7
r120 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.035 $Y=0.615
+ $X2=2.12 $Y2=0.7
r121 34 35 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.035 $Y=0.465
+ $X2=2.035 $Y2=0.615
r122 32 39 7.29036 $w=1.58e-07 $l=1.67929e-07 $layer=LI1_cond $X=2.595 $Y=1.6
+ $X2=2.71 $Y2=1.48
r123 32 50 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=2.595 $Y=1.6
+ $X2=1.265 $Y2=1.6
r124 28 31 27.4632 $w=2.08e-07 $l=5.2e-07 $layer=LI1_cond $X=1.06 $Y=0.36
+ $X2=1.58 $Y2=0.36
r125 26 34 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.95 $Y=0.36
+ $X2=2.035 $Y2=0.465
r126 26 31 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.95 $Y=0.36
+ $X2=1.58 $Y2=0.36
r127 25 49 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.345 $Y=1.54
+ $X2=0.935 $Y2=1.54
r128 23 45 26.4384 $w=2.53e-07 $l=5.85e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.245
r129 20 25 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=1.625
+ $X2=0.345 $Y2=1.54
r130 20 23 1.58178 $w=2.53e-07 $l=3.5e-08 $layer=LI1_cond $X=0.217 $Y=1.625
+ $X2=0.217 $Y2=1.66
r131 18 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.75 $Y=1.985
+ $X2=2.75 $Y2=1.325
r132 15 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.75 $Y=0.56
+ $X2=2.75 $Y2=0.995
r133 4 48 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=1.63
r134 3 44 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r135 3 23 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r136 2 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.455
+ $Y=0.235 $X2=1.58 $Y2=0.38
r137 1 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.235 $X2=1.06 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%A_109_297# 1 2 8 9 11 17
c26 9 0 1.7212e-19 $X=2.08 $Y=2.085
r27 16 17 35.4207 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=2.04 $Y=1.98
+ $X2=1.37 $Y2=1.98
r28 9 16 2.11255 $w=2.08e-07 $l=4e-08 $layer=LI1_cond $X=2.08 $Y=1.98 $X2=2.04
+ $Y2=1.98
r29 9 11 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.08 $Y=2.085
+ $X2=2.08 $Y2=2.3
r30 8 14 7.23718 $w=3.12e-07 $l=1.57003e-07 $layer=LI1_cond $X=0.825 $Y=1.985
+ $X2=0.68 $Y2=1.96
r31 8 17 30.2227 $w=1.98e-07 $l=5.45e-07 $layer=LI1_cond $X=0.825 $Y=1.985
+ $X2=1.37 $Y2=1.985
r32 2 16 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.04 $Y2=1.96
r33 2 11 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.485 $X2=2.04 $Y2=2.3
r34 1 14 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%VPWR 1 2 9 11 15 17 19 29 30 33 36
c47 15 0 8.13529e-20 $X=2.54 $Y=2.02
r48 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r52 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r53 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.58 $Y2=2.72
r54 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 26 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 21 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r58 19 33 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.607 $Y2=2.72
r59 19 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.43 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 17 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r61 17 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r62 13 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.72
r63 13 15 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=2.58 $Y=2.635
+ $X2=2.58 $Y2=2.02
r64 12 33 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.607 $Y2=2.72
r65 11 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.58 $Y2=2.72
r66 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=1.785 $Y2=2.72
r67 7 33 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.72
r68 7 9 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.607 $Y=2.635
+ $X2=1.607 $Y2=2.34
r69 2 15 300 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=2 $X=2.365
+ $Y=1.485 $X2=2.54 $Y2=2.02
r70 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=2.195 $X2=1.61 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%X 1 2 10 13 14 30
r16 19 30 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.005 $Y=1.915
+ $X2=3.005 $Y2=1.87
r17 13 30 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.005 $Y=1.85
+ $X2=3.005 $Y2=1.87
r18 13 14 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.005 $Y=1.935
+ $X2=3.005 $Y2=2.21
r19 13 19 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.005 $Y=1.935
+ $X2=3.005 $Y2=1.915
r20 11 13 50.6043 $w=2.78e-07 $l=1.2e-06 $layer=LI1_cond $X=3.05 $Y=0.585
+ $X2=3.05 $Y2=1.785
r21 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0.42
+ $X2=3.05 $Y2=0.585
r22 8 10 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.96 $Y=0.42 $X2=3.05
+ $Y2=0.42
r23 2 13 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.825
+ $Y=1.485 $X2=2.96 $Y2=1.96
r24 1 8 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.235 $X2=2.96 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A22O_1%VGND 1 2 7 9 13 15 17 27 28 34
c41 13 0 7.4275e-20 $X=2.54 $Y=0.36
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r43 28 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r44 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r45 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.54
+ $Y2=0
r46 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.99
+ $Y2=0
r47 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r48 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r49 21 24 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r50 20 23 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r51 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 18 31 5.99367 $w=1.7e-07 $l=2.73e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.272
+ $Y2=0
r53 18 20 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.69
+ $Y2=0
r54 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.54
+ $Y2=0
r55 17 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.07
+ $Y2=0
r56 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r59 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.36
r60 7 31 2.85413 $w=4.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.272 $Y2=0
r61 7 9 8.28054 $w=4.53e-07 $l=3.15e-07 $layer=LI1_cond $X=0.317 $Y=0.085
+ $X2=0.317 $Y2=0.4
r62 2 13 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.235 $X2=2.54 $Y2=0.36
r63 1 9 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends


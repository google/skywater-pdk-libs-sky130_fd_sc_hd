# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415000 1.075000 3.220000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.075000 4.480000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.715000 1.075000 5.860000 1.625000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.080000 1.725000 1.285000 ;
        RECT 1.175000 1.075000 1.505000 1.080000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.825000 1.285000 ;
        RECT 0.145000 1.285000 0.325000 1.625000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.955000 0.845000 2.125000 ;
        RECT 0.595000 1.455000 2.180000 1.625000 ;
        RECT 0.595000 1.625000 0.765000 1.955000 ;
        RECT 1.355000 0.655000 3.100000 0.825000 ;
        RECT 1.435000 1.625000 1.605000 2.125000 ;
        RECT 1.965000 0.825000 2.180000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.595000  0.085000 0.765000 0.545000 ;
        RECT 4.555000  0.085000 4.890000 0.465000 ;
        RECT 5.560000  0.085000 5.885000 0.885000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 2.270000 2.255000 2.940000 2.635000 ;
        RECT 3.550000 2.255000 4.220000 2.635000 ;
        RECT 4.765000 2.255000 5.435000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.295000 0.425000 0.465000 ;
      RECT 0.175000 0.465000 0.345000 0.715000 ;
      RECT 0.175000 0.715000 1.185000 0.885000 ;
      RECT 0.175000 1.795000 0.345000 2.295000 ;
      RECT 0.175000 2.295000 2.025000 2.465000 ;
      RECT 0.935000 0.295000 2.115000 0.465000 ;
      RECT 1.015000 0.465000 1.185000 0.715000 ;
      RECT 1.015000 1.795000 1.185000 2.295000 ;
      RECT 1.855000 1.795000 2.025000 1.915000 ;
      RECT 1.855000 1.915000 5.805000 2.085000 ;
      RECT 1.855000 2.085000 2.025000 2.295000 ;
      RECT 2.350000 0.295000 4.370000 0.465000 ;
      RECT 3.180000 1.795000 3.350000 1.915000 ;
      RECT 3.180000 2.085000 3.350000 2.465000 ;
      RECT 3.620000 0.635000 5.390000 0.805000 ;
      RECT 4.390000 1.795000 4.560000 1.915000 ;
      RECT 4.390000 2.085000 4.560000 2.465000 ;
      RECT 5.060000 0.275000 5.390000 0.635000 ;
      RECT 5.635000 1.795000 5.805000 1.915000 ;
      RECT 5.635000 2.085000 5.805000 2.465000 ;
  END
END sky130_fd_sc_hd__a32oi_2

* File: sky130_fd_sc_hd__or3b_2.pex.spice
* Created: Tue Sep  1 19:28:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR3B_2%C_N 3 7 9 10 17
r28 14 17 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r29 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.16
+ $X2=0.255 $Y2=1.53
r30 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r31 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r32 5 7 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=2.01
r33 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r34 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%A_176_21# 1 2 3 10 12 15 17 19 22 26 29 30 33
+ 35 39 42 44 45 49 54
r103 47 49 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.915 $Y=1.71
+ $X2=3.05 $Y2=1.71
r104 42 49 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.05 $Y=1.495
+ $X2=3.05 $Y2=1.71
r105 41 45 4.27425 $w=2.12e-07 $l=1.39929e-07 $layer=LI1_cond $X=3.05 $Y=0.825
+ $X2=2.982 $Y2=0.715
r106 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.05 $Y=0.825
+ $X2=3.05 $Y2=1.495
r107 37 45 4.27425 $w=2.12e-07 $l=1.21861e-07 $layer=LI1_cond $X=2.957 $Y=0.605
+ $X2=2.982 $Y2=0.715
r108 37 39 6.10117 $w=2.53e-07 $l=1.35e-07 $layer=LI1_cond $X=2.957 $Y=0.605
+ $X2=2.957 $Y2=0.47
r109 36 44 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.16 $Y=0.74
+ $X2=2.075 $Y2=0.78
r110 35 45 2.15711 $w=1.7e-07 $l=1.64024e-07 $layer=LI1_cond $X=2.83 $Y=0.74
+ $X2=2.982 $Y2=0.715
r111 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.83 $Y=0.74
+ $X2=2.16 $Y2=0.74
r112 31 44 1.34256 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.655
+ $X2=2.075 $Y2=0.78
r113 31 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.075 $Y=0.655
+ $X2=2.075 $Y2=0.47
r114 30 43 15.5991 $w=1.85e-07 $l=2.42384e-07 $layer=LI1_cond $X=1.595 $Y=0.82
+ $X2=1.36 $Y2=0.835
r115 29 44 5.16603 $w=1.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.99 $Y=0.82
+ $X2=2.075 $Y2=0.78
r116 29 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.99 $Y=0.82
+ $X2=1.595 $Y2=0.82
r117 27 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.36 $Y=1.16
+ $X2=1.375 $Y2=1.16
r118 27 51 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.36 $Y=1.16
+ $X2=0.955 $Y2=1.16
r119 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.36
+ $Y=1.16 $X2=1.36 $Y2=1.16
r120 24 43 1.22693 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.36 $Y=0.935 $X2=1.36
+ $Y2=0.835
r121 24 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.36 $Y=0.935
+ $X2=1.36 $Y2=1.16
r122 20 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.16
r123 20 22 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.985
r124 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=1.16
r125 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.375 $Y=0.995
+ $X2=1.375 $Y2=0.56
r126 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r127 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r128 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.16
r129 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r130 3 47 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.485 $X2=2.915 $Y2=1.685
r131 2 39 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.265 $X2=2.915 $Y2=0.47
r132 1 33 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.265 $X2=2.075 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%A 3 7 9 10 14 15
c45 7 0 1.45794e-19 $X=1.865 $Y=1.695
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=1.16 $X2=1.865 $Y2=1.16
r47 9 10 7.60125 $w=5.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.962 $Y=1.19
+ $X2=1.962 $Y2=1.53
r48 9 15 0.670698 $w=5.33e-07 $l=3e-08 $layer=LI1_cond $X=1.962 $Y=1.19
+ $X2=1.962 $Y2=1.16
r49 5 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=1.16
r50 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.865 $Y=1.325
+ $X2=1.865 $Y2=1.695
r51 1 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=0.995
+ $X2=1.865 $Y2=1.16
r52 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.865 $Y=0.995
+ $X2=1.865 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%B 3 6 7 8 12
c30 8 0 1.45794e-19 $X=2.91 $Y=2.125
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=2.28 $X2=2.285 $Y2=2.28
r32 7 8 22.0885 $w=2.38e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=2.245
+ $X2=2.995 $Y2=2.245
r33 7 13 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=2.535 $Y=2.245
+ $X2=2.285 $Y2=2.245
r34 3 6 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.285 $Y=0.475
+ $X2=2.285 $Y2=1.695
r35 1 12 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.285 $Y=2.145
+ $X2=2.285 $Y2=2.28
r36 1 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.285 $Y=2.145
+ $X2=2.285 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%A_27_47# 1 2 9 13 17 19 20 21 24 27 30 33 35
+ 36 37 41 42
c100 27 0 9.56717e-20 $X=2.49 $Y=1.87
r101 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.16 $X2=2.705 $Y2=1.16
r102 38 41 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.575 $Y=1.16
+ $X2=2.705 $Y2=1.16
r103 36 37 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.55 $Y=1.912
+ $X2=1.72 $Y2=1.912
r104 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=1.16
r105 29 30 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.575 $Y=1.325
+ $X2=2.575 $Y2=1.785
r106 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.49 $Y=1.87
+ $X2=2.575 $Y2=1.785
r107 27 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.49 $Y=1.87
+ $X2=1.72 $Y2=1.87
r108 26 35 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.765 $Y=1.955
+ $X2=0.68 $Y2=1.925
r109 26 36 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.765 $Y=1.955
+ $X2=1.55 $Y2=1.955
r110 24 35 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.68 $Y=1.81
+ $X2=0.68 $Y2=1.925
r111 23 24 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.68 $Y=0.905
+ $X2=0.68 $Y2=1.81
r112 22 33 1.45362 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.925
+ $X2=0.215 $Y2=1.925
r113 21 35 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=1.925
+ $X2=0.68 $Y2=1.925
r114 21 22 12.5266 $w=2.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=1.925
+ $X2=0.345 $Y2=1.925
r115 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.68 $Y2=0.905
r116 19 20 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.345 $Y2=0.82
r117 15 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.345 $Y2=0.82
r118 15 17 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.215 $Y=0.735
+ $X2=0.215 $Y2=0.455
r119 11 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.16
r120 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.705 $Y=1.325
+ $X2=2.705 $Y2=1.695
r121 7 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=1.16
r122 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.705 $Y=0.995
+ $X2=2.705 $Y2=0.475
r123 2 33 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.8 $X2=0.26 $Y2=1.975
r124 1 17 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%VPWR 1 2 9 13 15 17 22 32 33 36 39
c47 2 0 9.56717e-20 $X=1.45 $Y=1.485
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r49 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r52 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r54 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r55 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=1.59 $Y2=2.72
r56 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r58 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 23 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.91 $Y=2.72 $X2=0.73
+ $Y2=2.72
r61 23 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=1.59 $Y2=2.72
r63 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 17 36 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.73
+ $Y2=2.72
r65 17 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=2.72 $X2=0.23
+ $Y2=2.72
r66 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.635
+ $X2=1.59 $Y2=2.72
r69 11 13 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.59 $Y=2.635
+ $X2=1.59 $Y2=2.295
r70 7 36 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r71 7 9 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.295
r72 2 13 600 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.485 $X2=1.59 $Y2=2.295
r73 1 9 600 $w=1.7e-07 $l=5.86536e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.8 $X2=0.745 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%X 1 2 8 11 13
r30 13 18 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.155 $Y=0.43
+ $X2=1.02 $Y2=0.43
r31 13 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0.595
+ $X2=1.02 $Y2=0.43
r32 8 13 49.0479 $w=2.03e-07 $l=9e-07 $layer=LI1_cond $X=1.02 $Y=1.495 $X2=1.02
+ $Y2=0.595
r33 8 11 7.84479 $w=2.03e-07 $l=1.45e-07 $layer=LI1_cond $X=1.02 $Y=1.597
+ $X2=1.165 $Y2=1.597
r34 2 11 600 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.615
r35 1 13 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.165 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__OR3B_2%VGND 1 2 3 12 16 20 23 24 26 27 28 37 43 44
+ 47
r60 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r61 44 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r62 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r63 41 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.66 $Y=0 $X2=2.495
+ $Y2=0
r64 41 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.66 $Y=0 $X2=2.99
+ $Y2=0
r65 40 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r66 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r67 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.495
+ $Y2=0
r68 37 39 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.07
+ $Y2=0
r69 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r70 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r71 28 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r72 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 26 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.15
+ $Y2=0
r74 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.605
+ $Y2=0
r75 25 39 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=2.07
+ $Y2=0
r76 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.605
+ $Y2=0
r77 23 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r78 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r79 22 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=1.15
+ $Y2=0
r80 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r81 18 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.495 $Y2=0
r82 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.495 $Y=0.085
+ $X2=2.495 $Y2=0.4
r83 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0
r84 14 16 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0.4
r85 10 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r86 10 12 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.4
r87 3 20 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.265 $X2=2.495 $Y2=0.4
r88 2 16 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.605 $Y2=0.4
r89 1 12 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.4
.ends


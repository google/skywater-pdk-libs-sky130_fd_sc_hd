# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.990000 1.075000 5.895000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.780000 1.075000 4.820000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.885000 1.285000 ;
        RECT 0.605000 1.285000 0.885000 1.705000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.255000 1.385000 0.725000 ;
        RECT 1.055000 0.725000 2.225000 0.905000 ;
        RECT 1.055000 0.905000 1.455000 1.445000 ;
        RECT 1.055000 1.445000 2.225000 1.705000 ;
        RECT 1.895000 0.255000 2.225000 0.725000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.715000  0.085000 0.885000 0.905000 ;
        RECT 1.555000  0.085000 1.725000 0.555000 ;
        RECT 2.395000  0.085000 2.565000 0.555000 ;
        RECT 4.175000  0.085000 4.345000 0.555000 ;
        RECT 5.015000  0.085000 5.185000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.635000 2.215000 0.965000 2.635000 ;
        RECT 1.475000 2.215000 1.805000 2.635000 ;
        RECT 2.315000 2.215000 2.645000 2.635000 ;
        RECT 3.200000 2.135000 3.450000 2.635000 ;
        RECT 4.935000 1.835000 5.265000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.265000 0.545000 0.855000 ;
      RECT 0.085000 0.855000 0.255000 1.455000 ;
      RECT 0.085000 1.455000 0.435000 1.875000 ;
      RECT 0.085000 1.875000 2.565000 2.045000 ;
      RECT 0.085000 2.045000 0.435000 2.465000 ;
      RECT 1.625000 1.075000 2.565000 1.275000 ;
      RECT 2.395000 0.725000 3.585000 0.895000 ;
      RECT 2.395000 0.895000 2.565000 1.075000 ;
      RECT 2.395000 1.445000 2.905000 1.615000 ;
      RECT 2.395000 1.615000 2.565000 1.875000 ;
      RECT 2.735000 1.075000 3.135000 1.245000 ;
      RECT 2.735000 1.245000 2.905000 1.445000 ;
      RECT 2.805000 0.255000 4.005000 0.475000 ;
      RECT 2.815000 1.795000 4.380000 1.965000 ;
      RECT 2.815000 1.965000 2.985000 2.465000 ;
      RECT 3.235000 0.645000 3.585000 0.725000 ;
      RECT 3.395000 0.895000 3.585000 1.795000 ;
      RECT 3.685000 2.135000 3.925000 2.295000 ;
      RECT 3.685000 2.295000 4.765000 2.465000 ;
      RECT 3.755000 0.475000 4.005000 0.725000 ;
      RECT 3.755000 0.725000 5.710000 0.905000 ;
      RECT 4.135000 1.445000 4.380000 1.795000 ;
      RECT 4.135000 1.965000 4.380000 2.125000 ;
      RECT 4.515000 0.255000 4.845000 0.725000 ;
      RECT 4.595000 1.455000 5.710000 1.665000 ;
      RECT 4.595000 1.665000 4.765000 2.295000 ;
      RECT 5.355000 0.265000 5.710000 0.725000 ;
      RECT 5.435000 1.665000 5.710000 2.465000 ;
  END
END sky130_fd_sc_hd__o21ba_4

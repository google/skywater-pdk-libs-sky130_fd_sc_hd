* File: sky130_fd_sc_hd__dfxbp_2.spice
* Created: Tue Sep  1 19:04:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__dfxbp_2.pex.spice"
.subckt sky130_fd_sc_hd__dfxbp_2  VNB VPB CLK D VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_CLK_M1028_g N_A_27_47#_M1028_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_193_47#_M1020_d N_A_27_47#_M1020_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_381_47#_M1006_d N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0875538 AS=0.1092 PD=0.893846 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1009 N_A_466_413#_M1009_d N_A_27_47#_M1009_g N_A_381_47#_M1006_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0621 AS=0.0750462 PD=0.705 PS=0.766154 NRD=0 NRS=43.332 M=1
+ R=2.4 SA=75000.7 SB=75003.3 A=0.054 P=1.02 MULT=1
MM1016 A_592_47# N_A_193_47#_M1016_g N_A_466_413#_M1009_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0642462 AS=0.0621 PD=0.706154 PS=0.705 NRD=41.148 NRS=23.328 M=1
+ R=2.4 SA=75001.2 SB=75002.8 A=0.054 P=1.02 MULT=1
MM1026 N_VGND_M1026_d N_A_634_159#_M1026_g A_592_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0958472 AS=0.0749538 PD=0.859811 PS=0.823846 NRD=0 NRS=35.268 M=1 R=2.8
+ SA=75001.5 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1013 N_A_634_159#_M1013_d N_A_466_413#_M1013_g N_VGND_M1026_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.126592 AS=0.146053 PD=1.2736 PS=1.31019 NRD=0 NRS=30.936
+ M=1 R=4.26667 SA=75001.4 SB=75001 A=0.096 P=1.58 MULT=1
MM1031 N_A_891_413#_M1031_d N_A_193_47#_M1031_g N_A_634_159#_M1013_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0684 AS=0.071208 PD=0.74 PS=0.7164 NRD=3.324 NRS=24.996 M=1
+ R=2.4 SA=75002.8 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1004 A_1017_47# N_A_27_47#_M1004_g N_A_891_413#_M1031_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0684 PD=0.687692 PS=0.74 NRD=38.076 NRS=30 M=1 R=2.4
+ SA=75003.4 SB=75000.7 A=0.054 P=1.02 MULT=1
MM1011 N_VGND_M1011_d N_A_1059_315#_M1011_g A_1017_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_891_413#_M1015_g N_A_1059_315#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1015_d N_A_1059_315#_M1021_g N_Q_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1022_d N_A_1059_315#_M1022_g N_Q_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_1059_315#_M1002_g N_A_1589_47#_M1002_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=17.136 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1002_d N_A_1589_47#_M1003_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.121799 AS=0.08775 PD=1.19673 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_1589_47#_M1005_g N_Q_N_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.17225 AS=0.08775 PD=1.83 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_M1017_g N_A_27_47#_M1017_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_381_47#_M1023_d N_D_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.05775 AS=0.1092 PD=0.695 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_466_413#_M1012_d N_A_193_47#_M1012_g N_A_381_47#_M1023_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06825 AS=0.05775 PD=0.745 PS=0.695 NRD=14.0658 NRS=0 M=1
+ R=2.8 SA=75000.6 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1001 A_561_413# N_A_27_47#_M1001_g N_A_466_413#_M1012_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07665 AS=0.06825 PD=0.785 PS=0.745 NRD=59.7895 NRS=7.0329 M=1
+ R=2.8 SA=75001.1 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1029 N_VPWR_M1029_d N_A_634_159#_M1029_g A_561_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.128423 AS=0.07665 PD=0.904615 PS=0.785 NRD=111.384 NRS=59.7895 M=1 R=2.8
+ SA=75001.6 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_A_634_159#_M1008_d N_A_466_413#_M1008_g N_VPWR_M1029_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.140385 AS=0.229327 PD=1.37821 PS=1.61538 NRD=0 NRS=0 M=1
+ R=5 SA=75001.4 SB=75001 A=0.1125 P=1.8 MULT=1
MM1024 N_A_891_413#_M1024_d N_A_27_47#_M1024_g N_A_634_159#_M1008_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0567 AS=0.0786154 PD=0.69 PS=0.771795 NRD=0 NRS=23.443 M=1
+ R=2.8 SA=75002.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 A_975_413# N_A_193_47#_M1018_g N_A_891_413#_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.0567 PD=0.84 PS=0.69 NRD=72.693 NRS=0 M=1 R=2.8
+ SA=75003.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_1059_315#_M1007_g A_975_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0882 PD=1.37 PS=0.84 NRD=0 NRS=72.693 M=1 R=2.8 SA=75003.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_891_413#_M1025_g N_A_1059_315#_M1025_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0.9653 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1014 N_VPWR_M1025_d N_A_1059_315#_M1014_g N_Q_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_1059_315#_M1019_g N_Q_M1014_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.2
+ A=0.15 P=2.3 MULT=1
MM1010 N_VPWR_M1010_d N_A_1059_315#_M1010_g N_A_1589_47#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.120195 AS=0.1664 PD=1.04195 PS=1.8 NRD=18.4589 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1010_d N_A_1589_47#_M1027_g N_Q_N_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.187805 AS=0.135 PD=1.62805 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1030_d N_A_1589_47#_M1030_g N_Q_N_M1027_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.135 PD=2.53 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_98 VNB 0 1.97281e-19 $X=0.145 $Y=-0.085
c_204 VPB 0 2.47358e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__dfxbp_2.pxi.spice"
*
.ends
*
*

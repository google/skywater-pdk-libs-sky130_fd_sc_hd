* File: sky130_fd_sc_hd__a21boi_1.pex.spice
* Created: Tue Sep  1 18:51:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A21BOI_1%B1_N 1 2 3 5 6 8 13 15 16 20
r36 15 16 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16
+ $X2=0.22 $Y2=1.53
r37 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r38 11 20 145.524 $w=2.7e-07 $l=6.55e-07 $layer=POLY_cond $X=0.24 $Y=1.815
+ $X2=0.24 $Y2=1.16
r39 11 13 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.24 $Y=1.89
+ $X2=0.475 $Y2=1.89
r40 9 20 56.6543 $w=2.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=0.905
+ $X2=0.24 $Y2=1.16
r41 6 8 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.765 $Y=0.755
+ $X2=0.765 $Y2=0.445
r42 3 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.965
+ $X2=0.475 $Y2=1.89
r43 3 5 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.475 $Y=1.965
+ $X2=0.475 $Y2=2.275
r44 2 9 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.375 $Y=0.83
+ $X2=0.24 $Y2=0.905
r45 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.69 $Y=0.83
+ $X2=0.765 $Y2=0.755
r46 1 2 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=0.69 $Y=0.83
+ $X2=0.375 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%A_27_413# 1 2 7 11 13 15 17 21 25 26 28 35
+ 38 39
c67 25 0 1.83237e-19 $X=0.685 $Y=1.335
c68 17 0 1.96819e-19 $X=1.425 $Y=1.285
c69 11 0 1.36517e-19 $X=1.255 $Y=0.56
r70 37 38 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.63 $Y=0.715
+ $X2=0.63 $Y2=1.165
r71 35 37 9.81916 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=0.555 $Y=0.45
+ $X2=0.555 $Y2=0.715
r72 29 39 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=0.72 $Y=1.44
+ $X2=0.72 $Y2=1.285
r73 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.44 $X2=0.72 $Y2=1.44
r74 26 28 13.7276 $w=3.38e-07 $l=4.05e-07 $layer=LI1_cond $X=0.685 $Y=1.845
+ $X2=0.685 $Y2=1.44
r75 25 38 6.97447 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.685 $Y=1.335
+ $X2=0.685 $Y2=1.165
r76 25 28 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=0.685 $Y=1.335
+ $X2=0.685 $Y2=1.44
r77 19 26 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.225 $Y=1.945
+ $X2=0.685 $Y2=1.945
r78 19 21 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=2.27
r79 16 17 56.3681 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=1.255 $Y=1.285
+ $X2=1.425 $Y2=1.285
r80 13 17 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.425 $Y=1.385
+ $X2=1.425 $Y2=1.285
r81 13 15 192.8 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.425 $Y=1.385 $X2=1.425
+ $Y2=1.985
r82 9 16 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.255 $Y=1.185
+ $X2=1.255 $Y2=1.285
r83 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.255 $Y=1.185
+ $X2=1.255 $Y2=0.56
r84 8 39 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.855 $Y=1.285
+ $X2=0.72 $Y2=1.285
r85 7 16 24.8683 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.18 $Y=1.285 $X2=1.255
+ $Y2=1.285
r86 7 8 107.763 $w=2e-07 $l=3.25e-07 $layer=POLY_cond $X=1.18 $Y=1.285 $X2=0.855
+ $Y2=1.285
r87 2 21 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.27
r88 1 35 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.425
+ $Y=0.235 $X2=0.55 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%A1 3 6 8 9 10 15 17
c38 10 0 4.81425e-19 $X=2.07 $Y=1.19
c39 6 0 8.25831e-20 $X=1.855 $Y=1.985
r40 18 26 3.72573 $w=2.1e-07 $l=1.75e-07 $layer=LI1_cond $X=2.05 $Y=0.995
+ $X2=2.05 $Y2=1.17
r41 16 26 6.42075 $w=3.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.855 $Y=1.17
+ $X2=2.05 $Y2=1.17
r42 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.855 $Y2=0.995
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.16 $X2=1.855 $Y2=1.16
r44 10 26 0.658539 $w=3.48e-07 $l=2e-08 $layer=LI1_cond $X=2.07 $Y=1.17 $X2=2.05
+ $Y2=1.17
r45 9 18 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=2.05 $Y=0.85
+ $X2=2.05 $Y2=0.995
r46 8 9 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=2.05 $Y=0.51 $X2=2.05
+ $Y2=0.85
r47 4 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.325
+ $X2=1.855 $Y2=1.16
r48 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.855 $Y=1.325
+ $X2=1.855 $Y2=1.985
r49 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.845 $Y=0.56
+ $X2=1.845 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%A2 1 3 6 8 14
c24 8 0 1.34131e-20 $X=2.53 $Y=1.19
c25 6 0 1.48089e-19 $X=2.285 $Y=1.985
r26 12 14 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.285 $Y=1.16
+ $X2=2.485 $Y2=1.16
r27 10 12 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.275 $Y=1.16
+ $X2=2.285 $Y2=1.16
r28 8 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.16 $X2=2.485 $Y2=1.16
r29 4 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.325
+ $X2=2.285 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.285 $Y=1.325
+ $X2=2.285 $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 30 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.235 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 23 25 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 15 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.72
r59 11 13 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.07 $Y=2.635
+ $X2=2.07 $Y2=2.02
r60 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.635 $X2=0.69
+ $Y2=2.72
r61 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=2.635
+ $X2=0.69 $Y2=2.34
r62 2 13 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.485 $X2=2.07 $Y2=2.02
r63 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.065 $X2=0.69 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%Y 1 2 8 9 10 11 12 13 35
c36 35 0 6.917e-20 $X=1.457 $Y=1.195
r37 34 35 9.48845 $w=2.98e-07 $l=2.47e-07 $layer=LI1_cond $X=1.21 $Y=1.195
+ $X2=1.457 $Y2=1.195
r38 19 34 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.21 $Y=1.345
+ $X2=1.21 $Y2=1.195
r39 13 41 9.75371 $w=4.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.55 $Y=0.51
+ $X2=1.55 $Y2=0.795
r40 12 29 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.21 $Y=2.21 $X2=1.21
+ $Y2=2.31
r41 11 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.21 $Y=1.87
+ $X2=1.21 $Y2=2.21
r42 11 23 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.21 $Y=1.87 $X2=1.21
+ $Y2=1.63
r43 10 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.21 $Y=1.53 $X2=1.21
+ $Y2=1.63
r44 10 19 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.21 $Y=1.53
+ $X2=1.21 $Y2=1.345
r45 9 34 2.30489 $w=2.98e-07 $l=6e-08 $layer=LI1_cond $X=1.15 $Y=1.195 $X2=1.21
+ $Y2=1.195
r46 8 35 1.94584 $w=2.45e-07 $l=1.5e-07 $layer=LI1_cond $X=1.457 $Y=1.045
+ $X2=1.457 $Y2=1.195
r47 8 41 11.7596 $w=2.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.457 $Y=1.045
+ $X2=1.457 $Y2=0.795
r48 2 29 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=2.31
r49 2 23 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.21 $Y2=1.63
r50 1 13 182 $w=1.7e-07 $l=4.20862e-07 $layer=licon1_NDIFF $count=1 $X=1.33
+ $Y=0.235 $X2=1.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%A_300_297# 1 2 9 11 12 15
r16 13 15 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.5 $Y=1.725
+ $X2=2.5 $Y2=1.95
r17 11 13 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.415 $Y=1.625
+ $X2=2.5 $Y2=1.725
r18 11 12 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=2.415 $Y=1.625
+ $X2=1.735 $Y2=1.625
r19 7 12 6.82232 $w=2e-07 $l=1.39642e-07 $layer=LI1_cond $X=1.64 $Y=1.725
+ $X2=1.735 $Y2=1.625
r20 7 9 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.64 $Y=1.725 $X2=1.64
+ $Y2=1.95
r21 2 15 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.485 $X2=2.5 $Y2=1.95
r22 1 9 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.485 $X2=1.64 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HD__A21BOI_1%VGND 1 2 9 11 13 15 17 22 28 32
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r37 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r38 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r39 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r40 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r41 23 28 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.04
+ $Y2=0
r42 23 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=2.07
+ $Y2=0
r43 22 31 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.542
+ $Y2=0
r44 22 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.07
+ $Y2=0
r45 20 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r46 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 17 28 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=1.04
+ $Y2=0
r48 17 19 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.925 $Y=0 $X2=0.69
+ $Y2=0
r49 15 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r50 11 31 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.542 $Y2=0
r51 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.38
r52 7 28 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.04 $Y=0.085
+ $X2=1.04 $Y2=0
r53 7 9 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.04 $Y=0.085
+ $X2=1.04 $Y2=0.36
r54 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.35
+ $Y=0.235 $X2=2.49 $Y2=0.38
r55 1 9 91 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=2 $X=0.84
+ $Y=0.235 $X2=1.04 $Y2=0.36
.ends


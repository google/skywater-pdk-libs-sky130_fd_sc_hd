* File: sky130_fd_sc_hd__inv_4.pex.spice
* Created: Tue Sep  1 19:10:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__INV_4%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 32
+ 37 48
c77 13 0 5.55636e-20 $X=0.94 $Y=1.985
r78 46 48 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.57 $Y=1.16
+ $X2=1.78 $Y2=1.16
r79 44 46 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.36 $Y=1.16
+ $X2=1.57 $Y2=1.16
r80 43 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=1.36 $Y2=1.16
r81 42 43 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=1.16
+ $X2=0.94 $Y2=1.16
r82 37 42 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.445 $Y=1.16
+ $X2=0.52 $Y2=1.16
r83 37 39 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.445 $Y=1.16
+ $X2=0.27 $Y2=1.16
r84 32 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.57
+ $Y=1.16 $X2=1.57 $Y2=1.16
r85 31 32 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.57
+ $Y2=1.2
r86 30 31 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=1.2 $X2=1.15
+ $Y2=1.2
r87 29 30 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.23 $Y=1.2 $X2=0.69
+ $Y2=1.2
r88 29 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r89 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.16
r90 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.985
r91 22 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=0.995
+ $X2=1.78 $Y2=1.16
r92 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.78 $Y=0.995
+ $X2=1.78 $Y2=0.56
r93 18 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.16
r94 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.36 $Y=1.325
+ $X2=1.36 $Y2=1.985
r95 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=1.16
r96 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.36 $Y=0.995
+ $X2=1.36 $Y2=0.56
r97 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=0.94 $Y2=1.16
r98 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=0.94 $Y2=1.985
r99 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.16
r100 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r101 4 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.325
+ $X2=0.52 $Y2=1.16
r102 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.52 $Y=1.325
+ $X2=0.52 $Y2=1.985
r103 1 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__INV_4%VPWR 1 2 3 10 12 18 20 22 24 26 31 40 44
r35 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 35 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r38 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 32 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.15 $Y2=2.72
r41 32 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 31 43 3.64249 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=2.102 $Y2=2.72
r43 31 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 30 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r46 27 37 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r47 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 26 29 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r50 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 24 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 20 43 3.2727 $w=2.1e-07 $l=1.27609e-07 $layer=LI1_cond $X=2.01 $Y=2.635
+ $X2=2.102 $Y2=2.72
r53 20 22 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.01 $Y=2.635
+ $X2=2.01 $Y2=2.34
r54 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=2.635
+ $X2=1.15 $Y2=2.72
r55 16 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.15 $Y=2.635
+ $X2=1.15 $Y2=2
r56 12 15 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=0.262 $Y=1.66
+ $X2=0.262 $Y2=2.34
r57 10 37 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.197 $Y2=2.72
r58 10 15 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.262 $Y2=2.34
r59 3 22 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.485 $X2=1.99 $Y2=2.34
r60 2 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=1.485 $X2=1.15 $Y2=2
r61 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=2.34
r62 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__INV_4%Y 1 2 3 4 15 17 19 21 22 27 31 35 36 37 56
c66 37 0 5.55636e-20 $X=2.07 $Y=1.53
r67 55 56 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=1.59
+ $X2=1.405 $Y2=1.59
r68 44 55 27.2603 $w=1.88e-07 $l=4.67e-07 $layer=LI1_cond $X=2.037 $Y=1.59
+ $X2=1.57 $Y2=1.59
r69 37 44 1.92632 $w=1.88e-07 $l=3.3e-08 $layer=LI1_cond $X=2.07 $Y=1.59
+ $X2=2.037 $Y2=1.59
r70 37 44 1.08721 $w=2.63e-07 $l=2.5e-08 $layer=LI1_cond $X=2.037 $Y=1.47
+ $X2=2.037 $Y2=1.495
r71 36 37 12.1768 $w=2.63e-07 $l=2.8e-07 $layer=LI1_cond $X=2.037 $Y=1.19
+ $X2=2.037 $Y2=1.47
r72 35 43 2.03333 $w=1.78e-07 $l=3.3e-08 $layer=LI1_cond $X=2.07 $Y=0.815
+ $X2=2.037 $Y2=0.815
r73 35 36 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=2.037 $Y=0.92
+ $X2=2.037 $Y2=1.19
r74 35 43 0.652326 $w=2.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.037 $Y=0.92
+ $X2=2.037 $Y2=0.905
r75 31 55 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.57 $Y=2.34
+ $X2=1.57 $Y2=1.685
r76 25 43 28.7747 $w=1.78e-07 $l=4.67e-07 $layer=LI1_cond $X=1.57 $Y=0.815
+ $X2=2.037 $Y2=0.815
r77 25 27 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.57 $Y=0.725
+ $X2=1.57 $Y2=0.42
r78 24 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r79 24 56 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=1.405 $Y2=1.58
r80 21 25 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.815
+ $X2=1.57 $Y2=0.815
r81 21 22 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.405 $Y=0.815
+ $X2=0.895 $Y2=0.815
r82 17 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665 $X2=0.73
+ $Y2=1.58
r83 17 19 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.34
r84 13 22 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.895 $Y2=0.815
r85 13 15 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.73 $Y2=0.42
r86 4 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.485 $X2=1.57 $Y2=1.66
r87 4 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.485 $X2=1.57 $Y2=2.34
r88 3 34 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.485 $X2=0.73 $Y2=1.66
r89 3 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.485 $X2=0.73 $Y2=2.34
r90 2 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.57 $Y2=0.42
r91 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__INV_4%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r38 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r39 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r40 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r41 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r43 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r44 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.61
+ $Y2=0
r45 29 41 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.102
+ $Y2=0
r46 29 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.61
+ $Y2=0
r47 28 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r48 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r49 25 35 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r50 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r51 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.15
+ $Y2=0
r52 24 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.69
+ $Y2=0
r53 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r54 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r55 18 41 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.102 $Y2=0
r56 18 20 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=2.03 $Y=0.085 $X2=2.03
+ $Y2=0.385
r57 14 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r58 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.38
r59 10 35 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.197 $Y2=0
r60 10 12 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.262 $Y2=0.38
r61 3 20 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.235 $X2=1.99 $Y2=0.385
r62 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.15 $Y2=0.38
r63 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends


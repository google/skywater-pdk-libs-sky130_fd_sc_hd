* File: sky130_fd_sc_hd__nand2b_1.spice
* Created: Thu Aug 27 14:29:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand2b_1.pex.spice"
.subckt sky130_fd_sc_hd__nand2b_1  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_N_M1005_g N_A_27_93#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=37.812 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_206_47# N_B_M1001_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.121799 PD=0.92 PS=1.19673 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75000.5
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1000 N_Y_M1000_d N_A_27_93#_M1000_g A_206_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=14.76 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_27_93#_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.1092 PD=0.789718 PS=1.36 NRD=70.4866 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.205282 PD=1.27 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.4 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_93#_M1003_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.135 PD=2.53 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.8
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__nand2b_1.pxi.spice"
*
.ends
*
*

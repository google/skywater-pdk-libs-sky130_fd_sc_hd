* File: sky130_fd_sc_hd__a41oi_2.spice
* Created: Thu Aug 27 14:06:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a41oi_2.pex.spice"
.subckt sky130_fd_sc_hd__a41oi_2  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_B1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1000_d N_B1_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_317_47#_M1008_d N_A1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1011 N_A_317_47#_M1011_d N_A1_M1011_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1015 N_A_317_47#_M1011_d N_A2_M1015_g N_A_567_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_317_47#_M1016_d N_A2_M1016_g N_A_567_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_757_47#_M1005_d N_A3_M1005_g N_A_567_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1012 N_A_757_47#_M1012_d N_A3_M1012_g N_A_567_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 N_A_757_47#_M1012_d N_A4_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_757_47#_M1007_d N_A4_M1007_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_149_297#_M1006_d N_B1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75004.5 A=0.15 P=2.3 MULT=1
MM1018 N_A_149_297#_M1018_d N_B1_M1018_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.1 A=0.15 P=2.3 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_149_297#_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75003.6 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1002_d N_A1_M1019_g N_A_149_297#_M1019_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1010 N_A_149_297#_M1019_s N_A2_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1017 N_A_149_297#_M1017_d N_A2_M1017_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.135 PD=1.29 PS=1.27 NRD=2.9353 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A3_M1001_g N_A_149_297#_M1017_d VPB PHIGHVT L=0.15 W=1
+ AD=0.385 AS=0.145 PD=1.77 PS=1.29 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75002.7
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1013 N_VPWR_M1001_d N_A3_M1013_g N_A_149_297#_M1013_s VPB PHIGHVT L=0.15 W=1
+ AD=0.385 AS=0.135 PD=1.77 PS=1.27 NRD=12.7853 NRS=0 M=1 R=6.66667 SA=75003.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1004 N_A_149_297#_M1013_s N_A4_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.1
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1009 N_A_149_297#_M1009_d N_A4_M1009_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hd__a41oi_2.pxi.spice"
*
.ends
*
*

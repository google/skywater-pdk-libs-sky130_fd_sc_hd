* File: sky130_fd_sc_hd__o221ai_4.spice.pex
* Created: Thu Aug 27 14:37:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O221AI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 39 40
r59 38 40 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.51 $Y=1.16
+ $X2=1.75 $Y2=1.16
r60 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.51
+ $Y=1.16 $X2=1.51 $Y2=1.16
r61 36 38 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.33 $Y=1.16 $X2=1.51
+ $Y2=1.16
r62 35 36 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.91 $Y=1.16
+ $X2=1.33 $Y2=1.16
r63 33 35 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.49 $Y=1.16
+ $X2=0.91 $Y2=1.16
r64 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r65 29 39 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=1.51 $Y2=1.175
r66 29 34 36.8773 $w=1.98e-07 $l=6.65e-07 $layer=LI1_cond $X=1.155 $Y=1.175
+ $X2=0.49 $Y2=1.175
r67 25 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.16
r68 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.75 $Y=1.325
+ $X2=1.75 $Y2=1.985
r69 22 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=1.16
r70 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.75 $Y=0.995
+ $X2=1.75 $Y2=0.56
r71 18 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.16
r72 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.33 $Y=1.325
+ $X2=1.33 $Y2=1.985
r73 15 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=1.16
r74 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.56
r75 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.16
r76 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.91 $Y=1.325
+ $X2=0.91 $Y2=1.985
r77 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=1.16
r78 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.91 $Y=0.995
+ $X2=0.91 $Y2=0.56
r79 4 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.16
r80 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325 $X2=0.49
+ $Y2=1.985
r81 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.16
r82 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 30 31 32
+ 35 36 38 39 50
c111 35 0 1.93193e-19 $X=5.63 $Y=1.16
c112 32 0 1.61784e-19 $X=4.505 $Y=1.58
c113 30 0 1.07404e-19 $X=4.42 $Y=1.495
r114 48 50 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.415 $Y=1.16
+ $X2=3.53 $Y2=1.16
r115 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.16 $X2=3.415 $Y2=1.16
r116 46 48 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=3.11 $Y=1.16
+ $X2=3.415 $Y2=1.16
r117 44 46 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=3.11 $Y2=1.16
r118 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r119 41 44 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.69 $Y=1.16
+ $X2=2.735 $Y2=1.16
r120 39 49 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.415 $Y2=1.175
r121 39 45 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=2.735 $Y2=1.175
r122 38 49 51.0182 $w=1.98e-07 $l=9.2e-07 $layer=LI1_cond $X=4.335 $Y=1.175
+ $X2=3.415 $Y2=1.175
r123 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=1.16 $X2=5.63 $Y2=1.16
r124 33 35 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.63 $Y=1.495
+ $X2=5.63 $Y2=1.16
r125 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.465 $Y=1.58
+ $X2=5.63 $Y2=1.495
r126 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.465 $Y=1.58
+ $X2=4.505 $Y2=1.58
r127 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.42 $Y=1.495
+ $X2=4.505 $Y2=1.58
r128 29 38 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.42 $Y=1.275
+ $X2=4.335 $Y2=1.175
r129 29 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.42 $Y=1.275
+ $X2=4.42 $Y2=1.495
r130 25 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.16
r131 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.63 $Y=1.325
+ $X2=5.63 $Y2=1.985
r132 22 36 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=1.16
r133 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.63 $Y=0.995
+ $X2=5.63 $Y2=0.56
r134 18 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.16
r135 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.53 $Y=1.325
+ $X2=3.53 $Y2=1.985
r136 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=1.16
r137 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=0.56
r138 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.16
r139 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.985
r140 8 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=1.16
r141 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.11 $Y=0.995
+ $X2=3.11 $Y2=0.56
r142 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.16
r143 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.69 $Y=1.325
+ $X2=2.69 $Y2=1.985
r144 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.69 $Y2=1.16
r145 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.69 $Y=0.995
+ $X2=2.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 37 38
c75 37 0 1.20766e-19 $X=5.15 $Y=1.16
c76 6 0 1.61784e-19 $X=3.95 $Y=1.985
r77 36 38 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.15 $Y=1.16 $X2=5.21
+ $Y2=1.16
r78 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.15
+ $Y=1.16 $X2=5.15 $Y2=1.16
r79 34 36 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=5.15 $Y2=1.16
r80 33 34 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.37 $Y=1.16
+ $X2=4.79 $Y2=1.16
r81 31 33 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.95 $Y=1.16
+ $X2=4.37 $Y2=1.16
r82 29 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=1.16
+ $X2=5.15 $Y2=1.16
r83 25 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.16
r84 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.21 $Y=1.325
+ $X2=5.21 $Y2=1.985
r85 22 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=1.16
r86 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.21 $Y=0.995
+ $X2=5.21 $Y2=0.56
r87 18 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.16
r88 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.79 $Y=1.325
+ $X2=4.79 $Y2=1.985
r89 15 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=1.16
r90 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.79 $Y=0.995
+ $X2=4.79 $Y2=0.56
r91 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.16
r92 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.37 $Y=1.325
+ $X2=4.37 $Y2=1.985
r93 8 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=1.16
r94 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.37 $Y=0.995
+ $X2=4.37 $Y2=0.56
r95 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.325
+ $X2=3.95 $Y2=1.16
r96 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.95 $Y=1.325 $X2=3.95
+ $Y2=1.985
r97 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=1.16
r98 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995 $X2=3.95
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 31 32 34
+ 35 36 37 42 51 52
c128 8 0 2.92312e-20 $X=8.23 $Y=0.995
c129 1 0 2.92312e-20 $X=6.13 $Y=0.995
r130 50 52 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9 $Y=1.16 $X2=9.07
+ $Y2=1.16
r131 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9 $Y=1.16
+ $X2=9 $Y2=1.16
r132 48 50 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=8.65 $Y=1.16 $X2=9
+ $Y2=1.16
r133 42 51 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=8.535 $Y=1.175
+ $X2=9 $Y2=1.175
r134 41 48 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=8.32 $Y=1.16
+ $X2=8.65 $Y2=1.16
r135 41 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.32 $Y=1.16 $X2=8.23
+ $Y2=1.16
r136 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.32
+ $Y=1.16 $X2=8.32 $Y2=1.16
r137 38 42 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=8.42 $Y=1.175
+ $X2=8.535 $Y2=1.175
r138 38 40 3.99067 $w=2e-07 $l=1.33e-07 $layer=LI1_cond $X=8.42 $Y=1.175
+ $X2=8.287 $Y2=1.175
r139 36 40 3.0005 $w=2.65e-07 $l=1e-07 $layer=LI1_cond $X=8.287 $Y=1.275
+ $X2=8.287 $Y2=1.175
r140 36 37 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=8.287 $Y=1.275
+ $X2=8.287 $Y2=1.445
r141 34 37 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=8.155 $Y=1.53
+ $X2=8.287 $Y2=1.445
r142 34 35 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=8.155 $Y=1.53
+ $X2=6.295 $Y2=1.53
r143 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.13
+ $Y=1.16 $X2=6.13 $Y2=1.16
r144 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.13 $Y=1.445
+ $X2=6.295 $Y2=1.53
r145 29 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.13 $Y=1.445
+ $X2=6.13 $Y2=1.16
r146 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.07 $Y=1.325
+ $X2=9.07 $Y2=1.16
r147 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.07 $Y=1.325
+ $X2=9.07 $Y2=1.985
r148 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.07 $Y=0.995
+ $X2=9.07 $Y2=1.16
r149 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.07 $Y=0.995
+ $X2=9.07 $Y2=0.56
r150 18 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.16
r151 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.65 $Y=1.325
+ $X2=8.65 $Y2=1.985
r152 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=1.16
r153 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.65 $Y=0.995
+ $X2=8.65 $Y2=0.56
r154 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.16
r155 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.23 $Y=1.325
+ $X2=8.23 $Y2=1.985
r156 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=1.16
r157 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.23 $Y=0.995
+ $X2=8.23 $Y2=0.56
r158 4 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.16
r159 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.13 $Y=1.325
+ $X2=6.13 $Y2=1.985
r160 1 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=1.16
r161 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=0.995
+ $X2=6.13 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 35 41
c83 22 0 2.92312e-20 $X=7.81 $Y=0.995
r84 39 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=7.66 $Y=1.16
+ $X2=7.81 $Y2=1.16
r85 37 39 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.39 $Y=1.16
+ $X2=7.66 $Y2=1.16
r86 36 37 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.97 $Y=1.16
+ $X2=7.39 $Y2=1.16
r87 35 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.66
+ $Y=1.16 $X2=7.66 $Y2=1.16
r88 34 36 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.64 $Y=1.16
+ $X2=6.97 $Y2=1.16
r89 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.64
+ $Y=1.16 $X2=6.64 $Y2=1.16
r90 31 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.55 $Y=1.16 $X2=6.64
+ $Y2=1.16
r91 29 35 0.259574 $w=1.408e-06 $l=3e-08 $layer=LI1_cond $X=7.18 $Y=1.19
+ $X2=7.18 $Y2=1.16
r92 25 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=1.325
+ $X2=7.81 $Y2=1.16
r93 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.81 $Y=1.325
+ $X2=7.81 $Y2=1.985
r94 22 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=0.995
+ $X2=7.81 $Y2=1.16
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.81 $Y=0.995
+ $X2=7.81 $Y2=0.56
r96 18 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.16
r97 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.39 $Y=1.325
+ $X2=7.39 $Y2=1.985
r98 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=0.995
+ $X2=7.39 $Y2=1.16
r99 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.39 $Y=0.995
+ $X2=7.39 $Y2=0.56
r100 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.16
r101 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.97 $Y=1.325
+ $X2=6.97 $Y2=1.985
r102 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=1.16
r103 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.97 $Y=0.995
+ $X2=6.97 $Y2=0.56
r104 4 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.325
+ $X2=6.55 $Y2=1.16
r105 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.55 $Y=1.325
+ $X2=6.55 $Y2=1.985
r106 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=1.16
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 44 46
+ 51 52 54 55 57 58 59 61 87 95 100 103 106
c136 5 0 7.93326e-20 $X=5.705 $Y=1.485
r137 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r138 102 103 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.48 $Y=2.465
+ $X2=2.605 $Y2=2.465
r139 98 102 7.21165 $w=6.78e-07 $l=4.1e-07 $layer=LI1_cond $X=2.07 $Y=2.465
+ $X2=2.48 $Y2=2.465
r140 98 100 11.9076 $w=6.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.07 $Y=2.465
+ $X2=1.835 $Y2=2.465
r141 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r143 90 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r144 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r145 87 105 3.87948 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=9.407 $Y2=2.72
r146 87 89 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=8.97 $Y2=2.72
r147 86 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r148 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r149 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r150 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=8.05 $Y2=2.72
r151 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r153 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r154 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=5.75 $Y2=2.72
r155 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=5.75 $Y2=2.72
r156 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r157 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r158 74 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 73 103 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.605 $Y2=2.72
r160 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r161 70 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r162 70 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r163 69 100 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.835 $Y2=2.72
r164 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r165 67 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.12 $Y2=2.72
r166 67 69 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.245 $Y=2.72
+ $X2=1.61 $Y2=2.72
r167 65 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r168 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r169 62 92 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r170 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.69 $Y2=2.72
r171 61 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=1.12 $Y2=2.72
r172 61 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.995 $Y=2.72
+ $X2=0.69 $Y2=2.72
r173 59 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r174 59 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r175 57 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.05 $Y2=2.72
r176 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.44 $Y2=2.72
r177 56 89 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.97 $Y2=2.72
r178 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.44 $Y2=2.72
r179 54 79 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.755 $Y=2.72
+ $X2=5.75 $Y2=2.72
r180 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.755 $Y=2.72
+ $X2=5.88 $Y2=2.72
r181 53 82 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=6.21 $Y2=2.72
r182 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.005 $Y=2.72
+ $X2=5.88 $Y2=2.72
r183 51 73 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.195 $Y=2.72
+ $X2=2.99 $Y2=2.72
r184 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.195 $Y=2.72
+ $X2=3.32 $Y2=2.72
r185 50 76 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=3.45 $Y2=2.72
r186 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=3.32 $Y2=2.72
r187 46 49 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=9.28 $Y=1.62
+ $X2=9.28 $Y2=2.3
r188 44 105 3.26369 $w=2.5e-07 $l=1.64085e-07 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.407 $Y2=2.72
r189 44 49 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.28 $Y2=2.3
r190 40 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=2.635
+ $X2=8.44 $Y2=2.72
r191 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.44 $Y=2.635
+ $X2=8.44 $Y2=2.3
r192 36 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=2.635
+ $X2=5.88 $Y2=2.72
r193 36 38 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=5.88 $Y=2.635
+ $X2=5.88 $Y2=2.35
r194 32 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=2.635
+ $X2=3.32 $Y2=2.72
r195 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.32 $Y=2.635
+ $X2=3.32 $Y2=2.3
r196 28 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=2.72
r197 28 30 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.12 $Y=2.635
+ $X2=1.12 $Y2=1.99
r198 24 27 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=1.65
+ $X2=0.28 $Y2=2.33
r199 22 92 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.202 $Y2=2.72
r200 22 27 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=2.33
r201 7 49 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=2.3
r202 7 46 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=9.145
+ $Y=1.485 $X2=9.28 $Y2=1.62
r203 6 42 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.485 $X2=8.44 $Y2=2.3
r204 5 38 600 $w=1.7e-07 $l=9.48472e-07 $layer=licon1_PDIFF $count=1 $X=5.705
+ $Y=1.485 $X2=5.88 $Y2=2.35
r205 4 34 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.485 $X2=3.32 $Y2=2.3
r206 3 102 300 $w=1.7e-07 $l=1.09455e-06 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.485 $X2=2.48 $Y2=2.3
r207 2 30 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=0.985
+ $Y=1.485 $X2=1.12 $Y2=1.99
r208 1 27 400 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.33
r209 1 24 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%Y 1 2 3 4 5 6 7 8 25 33 38 41 44 45 48 49
+ 51 53 54 57 59 64 67 69 74
r130 74 79 25.9312 $w=2.47e-07 $l=5.25e-07 $layer=LI1_cond $X=6.235 $Y=1.955
+ $X2=6.76 $Y2=1.955
r131 69 72 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.6 $Y=1.87 $X2=7.6
+ $Y2=1.96
r132 63 64 6.9243 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.16 $Y=1.98
+ $X2=4.285 $Y2=1.98
r133 60 63 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=1.98 $X2=4.16
+ $Y2=1.98
r134 58 59 8.12479 $w=5.08e-07 $l=1.03e-07 $layer=LI1_cond $X=2.022 $Y=1.7
+ $X2=2.125 $Y2=1.7
r135 56 58 11.3041 $w=5.08e-07 $l=4.82e-07 $layer=LI1_cond $X=1.54 $Y=1.7
+ $X2=2.022 $Y2=1.7
r136 56 57 8.64074 $w=5.08e-07 $l=1.25e-07 $layer=LI1_cond $X=1.54 $Y=1.7
+ $X2=1.415 $Y2=1.7
r137 54 79 7.36982 $w=2.47e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.885 $Y=1.87
+ $X2=6.76 $Y2=1.955
r138 53 69 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.475 $Y=1.87
+ $X2=7.6 $Y2=1.87
r139 53 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.475 $Y=1.87
+ $X2=6.885 $Y2=1.87
r140 52 67 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.085 $Y=1.92
+ $X2=4.98 $Y2=1.92
r141 51 74 14.5318 $w=2.47e-07 $l=2.86967e-07 $layer=LI1_cond $X=5.965 $Y=1.92
+ $X2=6.235 $Y2=1.955
r142 51 52 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=5.965 $Y=1.92
+ $X2=5.085 $Y2=1.92
r143 49 67 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.875 $Y=1.92
+ $X2=4.98 $Y2=1.92
r144 49 64 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.875 $Y=1.92
+ $X2=4.285 $Y2=1.92
r145 48 60 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.08 $Y=1.835
+ $X2=4.08 $Y2=1.98
r146 47 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=4.08 $Y2=1.835
r147 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.995 $Y=1.53
+ $X2=4.08 $Y2=1.615
r148 45 59 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=3.995 $Y=1.53
+ $X2=2.125 $Y2=1.53
r149 44 58 6.13047 $w=2.05e-07 $l=2.55e-07 $layer=LI1_cond $X=2.022 $Y=1.445
+ $X2=2.022 $Y2=1.7
r150 43 44 31.3792 $w=2.03e-07 $l=5.8e-07 $layer=LI1_cond $X=2.022 $Y=0.865
+ $X2=2.022 $Y2=1.445
r151 39 56 4.91917 $w=2.5e-07 $l=2.55e-07 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.54 $Y2=1.7
r152 39 41 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.54 $Y=1.955
+ $X2=1.54 $Y2=1.96
r153 38 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.825 $Y=1.53
+ $X2=1.415 $Y2=1.53
r154 33 35 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.7 $Y=1.62 $X2=0.7
+ $Y2=2.3
r155 31 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.7 $Y=1.615
+ $X2=0.825 $Y2=1.53
r156 31 33 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.7 $Y=1.615 $X2=0.7
+ $Y2=1.62
r157 27 30 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=0.7 $Y=0.755
+ $X2=1.54 $Y2=0.755
r158 25 43 6.82754 $w=2.2e-07 $l=1.52709e-07 $layer=LI1_cond $X=1.92 $Y=0.755
+ $X2=2.022 $Y2=0.865
r159 25 30 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=1.92 $Y=0.755
+ $X2=1.54 $Y2=0.755
r160 8 72 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=7.465
+ $Y=1.485 $X2=7.6 $Y2=1.96
r161 7 79 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.485 $X2=6.76 $Y2=1.96
r162 6 67 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5 $Y2=1.96
r163 5 63 600 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.485 $X2=4.16 $Y2=1.96
r164 4 56 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.62
r165 4 41 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.405
+ $Y=1.485 $X2=1.54 $Y2=1.96
r166 3 35 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=2.3
r167 3 33 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.7 $Y2=1.62
r168 2 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.405
+ $Y=0.235 $X2=1.54 $Y2=0.73
r169 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A_553_297# 1 2 3 4 15 17 18 24 29 30 32 33
c39 4 0 1.13861e-19 $X=5.285 $Y=1.485
c40 3 0 1.07404e-19 $X=4.445 $Y=1.485
r41 32 33 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.42 $Y=2.32
+ $X2=5.255 $Y2=2.32
r42 30 33 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=5.255 $Y2=2.38
r43 28 30 6.9243 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.58 $Y=2.32
+ $X2=4.705 $Y2=2.32
r44 28 29 6.9243 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.58 $Y=2.32
+ $X2=4.455 $Y2=2.32
r45 24 29 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.825 $Y=2.38
+ $X2=4.455 $Y2=2.38
r46 20 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.72 $Y=2.295
+ $X2=3.825 $Y2=2.38
r47 20 22 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=3.72 $Y=2.295
+ $X2=3.72 $Y2=1.96
r48 19 22 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=3.72 $Y=1.955
+ $X2=3.72 $Y2=1.96
r49 17 19 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.615 $Y=1.87
+ $X2=3.72 $Y2=1.955
r50 17 18 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.615 $Y=1.87
+ $X2=3.025 $Y2=1.87
r51 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.9 $Y=1.955
+ $X2=3.025 $Y2=1.87
r52 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.9 $Y=1.955 $X2=2.9
+ $Y2=1.96
r53 4 32 600 $w=1.7e-07 $l=9.30054e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.42 $Y2=2.35
r54 3 28 600 $w=1.7e-07 $l=9.30054e-07 $layer=licon1_PDIFF $count=1 $X=4.445
+ $Y=1.485 $X2=4.58 $Y2=2.35
r55 2 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.605
+ $Y=1.485 $X2=3.74 $Y2=1.96
r56 1 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.765
+ $Y=1.485 $X2=2.9 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A_1241_297# 1 2 3 4 13 15 21 22 25 29 34 36
r49 36 38 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.18 $Y=2.3 $X2=7.18
+ $Y2=2.38
r50 32 34 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=2.32
+ $X2=6.505 $Y2=2.32
r51 27 40 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=1.955
+ $X2=8.86 $Y2=1.87
r52 27 29 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.86 $Y=1.955
+ $X2=8.86 $Y2=1.96
r53 23 40 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=1.785
+ $X2=8.86 $Y2=1.87
r54 23 25 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=1.785
+ $X2=8.86 $Y2=1.62
r55 21 40 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.735 $Y=1.87
+ $X2=8.86 $Y2=1.87
r56 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.735 $Y=1.87
+ $X2=8.145 $Y2=1.87
r57 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.02 $Y=2.295
+ $X2=8.02 $Y2=1.96
r58 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.02 $Y=1.955
+ $X2=8.145 $Y2=1.87
r59 17 20 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.02 $Y=1.955
+ $X2=8.02 $Y2=1.96
r60 16 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.305 $Y=2.38
+ $X2=7.18 $Y2=2.38
r61 15 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.895 $Y=2.38
+ $X2=8.02 $Y2=2.295
r62 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.895 $Y=2.38
+ $X2=7.305 $Y2=2.38
r63 13 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.055 $Y=2.38
+ $X2=7.18 $Y2=2.38
r64 13 34 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=7.055 $Y=2.38
+ $X2=6.505 $Y2=2.38
r65 4 29 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=1.96
r66 4 25 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.485 $X2=8.86 $Y2=1.62
r67 3 20 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.885
+ $Y=1.485 $X2=8.02 $Y2=1.96
r68 2 36 600 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.485 $X2=7.18 $Y2=2.3
r69 1 32 600 $w=1.7e-07 $l=9.30054e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.34 $Y2=2.35
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A_27_47# 1 2 3 4 5 6 7 22 24 38
r46 36 38 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=4.58 $Y=0.365
+ $X2=5.42 $Y2=0.365
r47 34 36 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=3.74 $Y=0.365
+ $X2=4.58 $Y2=0.365
r48 32 34 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=2.9 $Y=0.365
+ $X2=3.74 $Y2=0.365
r49 30 32 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=1.96 $Y=0.365
+ $X2=2.9 $Y2=0.365
r50 28 30 44.0024 $w=2.18e-07 $l=8.4e-07 $layer=LI1_cond $X=1.12 $Y=0.365
+ $X2=1.96 $Y2=0.365
r51 26 41 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.365
+ $X2=0.24 $Y2=0.365
r52 26 28 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=0.365 $Y=0.365
+ $X2=1.12 $Y2=0.365
r53 22 41 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.24 $Y=0.475
+ $X2=0.24 $Y2=0.365
r54 22 24 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=0.475
+ $X2=0.24 $Y2=0.73
r55 7 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.235 $X2=5.42 $Y2=0.39
r56 6 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.58 $Y2=0.39
r57 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.74 $Y2=0.39
r58 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.235 $X2=2.9 $Y2=0.39
r59 3 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.235 $X2=1.96 $Y2=0.39
r60 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.235 $X2=1.12 $Y2=0.39
r61 1 41 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
r62 1 24 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%A_471_47# 1 2 3 4 5 6 7 8 9 40 42 46 48 52
+ 54 58 60 64 67 69 70 71 72
c131 72 0 2.92312e-20 $X=8.44 $Y=0.815
c132 71 0 2.92312e-20 $X=7.6 $Y=0.815
c133 70 0 2.92312e-20 $X=6.76 $Y=0.815
r134 62 64 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.28 $Y=0.725
+ $X2=9.28 $Y2=0.39
r135 61 72 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=0.815
+ $X2=8.44 $Y2=0.815
r136 60 62 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=9.115 $Y=0.815
+ $X2=9.28 $Y2=0.725
r137 60 61 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=9.115 $Y=0.815
+ $X2=8.605 $Y2=0.815
r138 56 72 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.44 $Y=0.725
+ $X2=8.44 $Y2=0.815
r139 56 58 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.44 $Y=0.725
+ $X2=8.44 $Y2=0.39
r140 55 71 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=7.765 $Y=0.82
+ $X2=7.6 $Y2=0.815
r141 54 72 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=8.44 $Y2=0.815
r142 54 55 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=7.765 $Y2=0.82
r143 50 71 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.6 $Y=0.725 $X2=7.6
+ $Y2=0.815
r144 50 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.6 $Y=0.725
+ $X2=7.6 $Y2=0.39
r145 49 70 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=0.815
+ $X2=6.76 $Y2=0.815
r146 48 71 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=0.815
+ $X2=7.6 $Y2=0.815
r147 48 49 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.435 $Y=0.815
+ $X2=6.925 $Y2=0.815
r148 44 70 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.76 $Y=0.725
+ $X2=6.76 $Y2=0.815
r149 44 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.76 $Y=0.725
+ $X2=6.76 $Y2=0.39
r150 42 70 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.595 $Y=0.82
+ $X2=6.76 $Y2=0.815
r151 42 69 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.595 $Y=0.82
+ $X2=6.085 $Y2=0.82
r152 38 69 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=0.775
+ $X2=6.085 $Y2=0.775
r153 38 67 21.4044 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=5.92 $Y=0.775
+ $X2=5.465 $Y2=0.775
r154 38 40 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.92 $Y=0.645
+ $X2=5.92 $Y2=0.39
r155 37 67 29.4701 $w=1.73e-07 $l=4.65e-07 $layer=LI1_cond $X=5 $Y=0.732
+ $X2=5.465 $Y2=0.732
r156 35 37 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=4.16 $Y=0.732 $X2=5
+ $Y2=0.732
r157 33 35 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=3.32 $Y=0.732
+ $X2=4.16 $Y2=0.732
r158 30 33 53.2364 $w=1.73e-07 $l=8.4e-07 $layer=LI1_cond $X=2.48 $Y=0.732
+ $X2=3.32 $Y2=0.732
r159 9 64 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.145
+ $Y=0.235 $X2=9.28 $Y2=0.39
r160 8 58 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.305
+ $Y=0.235 $X2=8.44 $Y2=0.39
r161 7 52 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.465
+ $Y=0.235 $X2=7.6 $Y2=0.39
r162 6 46 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.625
+ $Y=0.235 $X2=6.76 $Y2=0.39
r163 5 38 182 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.92 $Y2=0.73
r164 5 40 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=5.705
+ $Y=0.235 $X2=5.92 $Y2=0.39
r165 4 37 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5 $Y2=0.73
r166 3 35 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.16 $Y2=0.73
r167 2 33 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.235 $X2=3.32 $Y2=0.73
r168 1 30 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=2.355
+ $Y=0.235 $X2=2.48 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O221AI_4%VGND 1 2 3 4 15 17 21 25 29 31 32 34 35 37
+ 38 39 56 57 60
r116 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r117 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r118 54 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r119 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r120 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r121 51 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r122 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r123 48 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.265 $Y=0 $X2=7.18
+ $Y2=0
r124 48 50 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=7.59 $Y2=0
r125 47 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r126 46 47 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r127 42 46 390.139 $w=1.68e-07 $l=5.98e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=6.21
+ $Y2=0
r128 39 47 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=6.21
+ $Y2=0
r129 39 42 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r130 37 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.775 $Y=0
+ $X2=8.51 $Y2=0
r131 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.775 $Y=0 $X2=8.86
+ $Y2=0
r132 36 56 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.945 $Y=0
+ $X2=9.43 $Y2=0
r133 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.945 $Y=0 $X2=8.86
+ $Y2=0
r134 34 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.935 $Y=0 $X2=7.59
+ $Y2=0
r135 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=0 $X2=8.02
+ $Y2=0
r136 33 53 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=8.51 $Y2=0
r137 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.02
+ $Y2=0
r138 31 46 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.255 $Y=0 $X2=6.21
+ $Y2=0
r139 31 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=0 $X2=6.34
+ $Y2=0
r140 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0
r141 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.86 $Y=0.085
+ $X2=8.86 $Y2=0.39
r142 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0
r143 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.02 $Y=0.085
+ $X2=8.02 $Y2=0.39
r144 19 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0
r145 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0.39
r146 18 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=0 $X2=6.34
+ $Y2=0
r147 17 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=0 $X2=7.18
+ $Y2=0
r148 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.095 $Y=0
+ $X2=6.425 $Y2=0
r149 13 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=0.085
+ $X2=6.34 $Y2=0
r150 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.34 $Y=0.085
+ $X2=6.34 $Y2=0.39
r151 4 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.235 $X2=8.86 $Y2=0.39
r152 3 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.885
+ $Y=0.235 $X2=8.02 $Y2=0.39
r153 2 21 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.045
+ $Y=0.235 $X2=7.18 $Y2=0.39
r154 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.205
+ $Y=0.235 $X2=6.34 $Y2=0.39
.ends


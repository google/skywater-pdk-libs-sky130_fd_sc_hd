* File: sky130_fd_sc_hd__a22oi_1.pxi.spice
* Created: Thu Aug 27 14:02:50 2020
* 
x_PM_SKY130_FD_SC_HD__A22OI_1%B2 N_B2_M1007_g N_B2_M1004_g B2 B2 N_B2_c_52_n
+ N_B2_c_53_n PM_SKY130_FD_SC_HD__A22OI_1%B2
x_PM_SKY130_FD_SC_HD__A22OI_1%B1 N_B1_M1000_g N_B1_M1003_g B1 B1 N_B1_c_83_n
+ N_B1_c_84_n PM_SKY130_FD_SC_HD__A22OI_1%B1
x_PM_SKY130_FD_SC_HD__A22OI_1%A1 N_A1_M1001_g N_A1_M1006_g A1 A1 N_A1_c_123_n
+ N_A1_c_124_n A1 PM_SKY130_FD_SC_HD__A22OI_1%A1
x_PM_SKY130_FD_SC_HD__A22OI_1%A2 N_A2_M1002_g N_A2_M1005_g A2 N_A2_c_157_n
+ N_A2_c_158_n N_A2_c_159_n PM_SKY130_FD_SC_HD__A22OI_1%A2
x_PM_SKY130_FD_SC_HD__A22OI_1%Y N_Y_M1000_d N_Y_M1001_s N_Y_M1004_s N_Y_M1003_d
+ N_Y_c_193_n N_Y_c_194_n N_Y_c_195_n N_Y_c_190_n N_Y_c_196_n N_Y_c_235_n
+ N_Y_c_191_n N_Y_c_239_n N_Y_c_192_n N_Y_c_198_n N_Y_c_207_n Y Y Y N_Y_c_200_n
+ PM_SKY130_FD_SC_HD__A22OI_1%Y
x_PM_SKY130_FD_SC_HD__A22OI_1%A_109_297# N_A_109_297#_M1004_d
+ N_A_109_297#_M1006_d N_A_109_297#_c_281_n N_A_109_297#_c_282_n
+ N_A_109_297#_c_284_n PM_SKY130_FD_SC_HD__A22OI_1%A_109_297#
x_PM_SKY130_FD_SC_HD__A22OI_1%VPWR N_VPWR_M1006_s N_VPWR_M1005_d N_VPWR_c_309_n
+ N_VPWR_c_310_n N_VPWR_c_311_n VPWR N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_308_n PM_SKY130_FD_SC_HD__A22OI_1%VPWR
x_PM_SKY130_FD_SC_HD__A22OI_1%VGND N_VGND_M1007_s N_VGND_M1002_d N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n VGND N_VGND_c_352_n
+ N_VGND_c_353_n PM_SKY130_FD_SC_HD__A22OI_1%VGND
cc_1 VNB B2 0.024374f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_2 VNB N_B2_c_52_n 0.0254443f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_3 VNB N_B2_c_53_n 0.0175319f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_4 VNB B1 0.00533903f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_5 VNB B1 0.00528218f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_B1_c_83_n 0.0240214f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_7 VNB N_B1_c_84_n 0.0190064f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_8 VNB A1 0.00444945f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_9 VNB N_A1_c_123_n 0.0307265f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_10 VNB N_A1_c_124_n 0.0188105f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=0.995
cc_11 VNB A1 0.00192528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_c_157_n 0.022195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_158_n 0.00302548f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_14 VNB N_A2_c_159_n 0.0190295f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_15 VNB N_Y_c_190_n 0.0145699f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_16 VNB N_Y_c_191_n 0.00785825f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_192_n 0.021962f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_308_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_348_n 0.0119082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_349_n 0.0184558f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_21 VNB N_VGND_c_350_n 0.0123324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_351_n 0.0149926f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_23 VNB N_VGND_c_352_n 0.0415342f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=0.85
cc_24 VNB N_VGND_c_353_n 0.163698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_B2_M1004_g 0.0252917f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_26 VPB N_B2_c_52_n 0.00474892f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_27 VPB N_B1_M1003_g 0.0253102f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_28 VPB N_B1_c_83_n 0.00485592f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_29 VPB N_A1_M1006_g 0.0245208f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_30 VPB N_A1_c_123_n 0.00718746f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_31 VPB N_A2_M1005_g 0.0223895f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_32 VPB N_A2_c_157_n 0.00424854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A2_c_158_n 0.00116599f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_34 VPB N_Y_c_193_n 0.0110511f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_35 VPB N_Y_c_194_n 0.00746643f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_36 VPB N_Y_c_195_n 0.025859f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.325
cc_37 VPB N_Y_c_196_n 0.0092337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_Y_c_192_n 0.00919843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_198_n 0.00250932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB Y 0.0232628f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_Y_c_200_n 8.28086e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_109_297#_c_281_n 0.00808846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_109_297#_c_282_n 5.01725e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_44 VPB N_VPWR_c_309_n 0.00572125f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_45 VPB N_VPWR_c_310_n 0.0115786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_311_n 0.0045947f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_47 VPB N_VPWR_c_312_n 0.0358463f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=0.85
cc_48 VPB N_VPWR_c_313_n 0.0149232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_314_n 0.00578832f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_308_n 0.0476202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_B2_M1004_g N_B1_M1003_g 0.0436634f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_52 B2 B1 0.010577f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_53 B2 B1 0.0161017f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_54 N_B2_c_52_n B1 6.83135e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_55 B2 N_B1_c_83_n 7.05986e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_56 N_B2_c_52_n N_B1_c_83_n 0.0338773f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_57 B2 N_B1_c_84_n 0.00195579f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_58 N_B2_c_53_n N_B1_c_84_n 0.0338773f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_59 N_B2_M1004_g N_Y_c_193_n 0.0017138f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_60 B2 N_Y_c_193_n 0.0266308f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_61 N_B2_c_52_n N_Y_c_193_n 0.00296763f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B2_M1004_g N_Y_c_194_n 7.12665e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_63 N_B2_M1004_g N_Y_c_195_n 0.00966083f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_64 N_B2_c_53_n N_Y_c_190_n 7.24737e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_65 N_B2_M1004_g N_Y_c_207_n 0.00819053f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_66 N_B2_M1004_g Y 0.00901884f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_67 B2 Y 0.0113279f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_68 N_B2_M1004_g N_VPWR_c_312_n 0.00357835f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_69 N_B2_M1004_g N_VPWR_c_308_n 0.00620759f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_70 B2 N_VGND_M1007_s 0.00240421f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_71 B2 N_VGND_c_349_n 0.0300914f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_72 N_B2_c_52_n N_VGND_c_349_n 4.51734e-19 $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B2_c_53_n N_VGND_c_349_n 0.0212578f $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_74 B2 N_VGND_c_353_n 0.00275279f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_B2_c_53_n N_VGND_c_353_n 7.20442e-19 $X=0.41 $Y=0.995 $X2=0 $Y2=0
cc_76 B1 A1 0.0240915f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_77 N_B1_c_83_n A1 2.15452e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_78 B1 N_A1_c_123_n 2.99118e-19 $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_79 B1 N_A1_c_123_n 8.24852e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_80 N_B1_c_83_n N_A1_c_123_n 0.00824835f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_81 B1 A1 0.0130934f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_82 N_B1_c_83_n A1 5.81957e-19 $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_83 B1 N_Y_M1000_d 0.00596846f $X=1.07 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_84 N_B1_M1003_g N_Y_c_195_n 0.00147562f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_85 B1 N_Y_c_190_n 0.0191219f $X=1.07 $Y=0.765 $X2=0 $Y2=0
cc_86 B1 N_Y_c_190_n 0.00374973f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 N_B1_c_83_n N_Y_c_190_n 0.00137136f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B1_c_84_n N_Y_c_190_n 0.00810253f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_M1003_g N_Y_c_198_n 0.00179258f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_90 N_B1_M1003_g N_Y_c_207_n 0.0066112f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_91 N_B1_M1003_g Y 0.012932f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_92 B1 Y 0.0346852f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B1_c_83_n Y 0.00350026f $X=0.93 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B1_M1003_g N_Y_c_200_n 9.76525e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_95 N_B1_M1003_g N_A_109_297#_c_281_n 0.0144566f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_A_109_297#_c_284_n 0.00207757f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_97 N_B1_M1003_g N_VPWR_c_309_n 0.00247143f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_98 N_B1_M1003_g N_VPWR_c_312_n 0.00357877f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_VPWR_c_308_n 0.00657948f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B1_c_84_n N_VGND_c_349_n 0.00296089f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_101 N_B1_c_84_n N_VGND_c_352_n 0.0042613f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_84_n N_VGND_c_353_n 0.0081372f $X=0.92 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A1_M1006_g N_A2_M1005_g 0.042874f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_104 N_A1_c_123_n N_A2_c_157_n 0.0378724f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_105 A1 N_A2_c_158_n 0.00388011f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_106 N_A1_c_123_n N_A2_c_158_n 0.00326379f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_107 A1 N_A2_c_158_n 0.0158715f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_108 N_A1_c_124_n N_A2_c_159_n 0.0378724f $X=1.712 $Y=0.995 $X2=0 $Y2=0
cc_109 A1 N_Y_M1001_s 0.0036585f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_110 A1 N_Y_c_190_n 0.0158418f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A1_c_123_n N_Y_c_190_n 6.49925e-19 $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_c_124_n N_Y_c_190_n 0.0122623f $X=1.712 $Y=0.995 $X2=0 $Y2=0
cc_113 A1 N_Y_c_190_n 0.00295871f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_114 N_A1_M1006_g N_Y_c_196_n 0.00661917f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A1_c_123_n Y 0.00560998f $X=1.675 $Y=1.16 $X2=0 $Y2=0
cc_116 A1 Y 0.0254603f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_117 N_A1_M1006_g N_Y_c_200_n 0.0098405f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A1_M1006_g N_A_109_297#_c_281_n 0.00282228f $X=1.83 $Y=1.985 $X2=0
+ $Y2=0
cc_119 N_A1_M1006_g N_A_109_297#_c_282_n 0.0127274f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_120 N_A1_M1006_g N_VPWR_c_309_n 0.0110212f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_121 N_A1_M1006_g N_VPWR_c_313_n 0.00273041f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A1_M1006_g N_VPWR_c_308_n 0.00339032f $X=1.83 $Y=1.985 $X2=0 $Y2=0
cc_123 N_A1_c_124_n N_VGND_c_352_n 0.00357877f $X=1.712 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A1_c_124_n N_VGND_c_353_n 0.00641668f $X=1.712 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A2_c_159_n N_Y_c_190_n 0.0055472f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_M1005_g N_Y_c_196_n 0.016464f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_127 N_A2_c_157_n N_Y_c_196_n 0.00269153f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A2_c_158_n N_Y_c_196_n 0.0216323f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A2_c_159_n N_Y_c_235_n 0.00673349f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A2_c_157_n N_Y_c_191_n 0.00304803f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A2_c_158_n N_Y_c_191_n 0.0130625f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A2_c_159_n N_Y_c_191_n 0.0109928f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A2_c_158_n N_Y_c_239_n 0.0072757f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_159_n N_Y_c_239_n 0.00134585f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A2_M1005_g N_Y_c_192_n 0.00523374f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_136 N_A2_c_157_n N_Y_c_192_n 0.00755993f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A2_c_158_n N_Y_c_192_n 0.0247426f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A2_c_159_n N_Y_c_192_n 0.00536692f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_M1005_g N_VPWR_c_309_n 0.00119769f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A2_M1005_g N_VPWR_c_311_n 0.00316907f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A2_M1005_g N_VPWR_c_313_n 0.00585385f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A2_M1005_g N_VPWR_c_308_n 0.0115941f $X=2.25 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A2_c_159_n N_VGND_c_351_n 0.00951416f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A2_c_159_n N_VGND_c_352_n 0.00423331f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A2_c_159_n N_VGND_c_353_n 0.0066759f $X=2.25 $Y=0.995 $X2=0 $Y2=0
cc_146 N_Y_c_207_n N_A_109_297#_M1004_d 0.00312752f $X=0.935 $Y=2.36 $X2=-0.19
+ $Y2=-0.24
cc_147 Y N_A_109_297#_M1004_d 0.00166529f $X=1.615 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_148 N_Y_c_196_n N_A_109_297#_M1006_d 0.00373815f $X=2.505 $Y=1.58 $X2=0 $Y2=0
cc_149 N_Y_M1003_d N_A_109_297#_c_281_n 0.00642559f $X=0.965 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_Y_c_198_n N_A_109_297#_c_281_n 0.0190248f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_151 N_Y_c_207_n N_A_109_297#_c_281_n 0.00597442f $X=0.935 $Y=2.36 $X2=0 $Y2=0
cc_152 Y N_A_109_297#_c_281_n 0.0317057f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_153 N_Y_c_196_n N_A_109_297#_c_282_n 0.01198f $X=2.505 $Y=1.58 $X2=0 $Y2=0
cc_154 Y N_A_109_297#_c_282_n 0.00883438f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_155 N_Y_c_200_n N_A_109_297#_c_282_n 0.0165653f $X=1.84 $Y=1.555 $X2=0 $Y2=0
cc_156 N_Y_c_207_n N_A_109_297#_c_284_n 0.0118327f $X=0.935 $Y=2.36 $X2=0 $Y2=0
cc_157 Y N_A_109_297#_c_284_n 0.0257775f $X=1.615 $Y=1.53 $X2=0 $Y2=0
cc_158 Y N_VPWR_M1006_s 0.00200719f $X=1.615 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_159 N_Y_c_200_n N_VPWR_M1006_s 0.00169526f $X=1.84 $Y=1.555 $X2=-0.19
+ $Y2=-0.24
cc_160 N_Y_c_196_n N_VPWR_M1005_d 0.00623784f $X=2.505 $Y=1.58 $X2=0 $Y2=0
cc_161 N_Y_c_198_n N_VPWR_c_309_n 0.018382f $X=1.1 $Y=2.34 $X2=0 $Y2=0
cc_162 N_Y_c_196_n N_VPWR_c_311_n 0.019004f $X=2.505 $Y=1.58 $X2=0 $Y2=0
cc_163 N_Y_c_194_n N_VPWR_c_312_n 0.021178f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_164 N_Y_c_207_n N_VPWR_c_312_n 0.0481435f $X=0.935 $Y=2.36 $X2=0 $Y2=0
cc_165 N_Y_M1004_s N_VPWR_c_308_n 0.00209319f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_166 N_Y_M1003_d N_VPWR_c_308_n 0.00209344f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_167 N_Y_c_194_n N_VPWR_c_308_n 0.0124992f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_168 N_Y_c_207_n N_VPWR_c_308_n 0.030037f $X=0.935 $Y=2.36 $X2=0 $Y2=0
cc_169 N_Y_c_191_n N_VGND_M1002_d 0.00799132f $X=2.505 $Y=0.74 $X2=0 $Y2=0
cc_170 N_Y_c_192_n N_VGND_M1002_d 0.00108013f $X=2.59 $Y=1.495 $X2=0 $Y2=0
cc_171 N_Y_c_190_n N_VGND_c_349_n 0.0137634f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_172 N_Y_c_191_n N_VGND_c_350_n 7.81766e-19 $X=2.505 $Y=0.74 $X2=0 $Y2=0
cc_173 N_Y_c_191_n N_VGND_c_351_n 0.0249844f $X=2.505 $Y=0.74 $X2=0 $Y2=0
cc_174 N_Y_c_190_n N_VGND_c_352_n 0.0783673f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_175 N_Y_c_191_n N_VGND_c_352_n 0.00254364f $X=2.505 $Y=0.74 $X2=0 $Y2=0
cc_176 N_Y_M1000_d N_VGND_c_353_n 0.00209344f $X=0.925 $Y=0.235 $X2=0 $Y2=0
cc_177 N_Y_M1001_s N_VGND_c_353_n 0.00209344f $X=1.495 $Y=0.235 $X2=0 $Y2=0
cc_178 N_Y_c_190_n N_VGND_c_353_n 0.0478016f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_179 N_Y_c_191_n N_VGND_c_353_n 0.00702372f $X=2.505 $Y=0.74 $X2=0 $Y2=0
cc_180 N_Y_c_190_n A_381_47# 9.3379e-19 $X=1.945 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_181 N_Y_c_239_n A_381_47# 0.00149057f $X=2.125 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_182 N_A_109_297#_c_282_n N_VPWR_M1006_s 0.00529516f $X=1.955 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_183 N_A_109_297#_c_281_n N_VPWR_c_309_n 0.00258466f $X=1.065 $Y=1.94 $X2=0
+ $Y2=0
cc_184 N_A_109_297#_c_282_n N_VPWR_c_309_n 0.0169644f $X=1.955 $Y=1.935 $X2=0
+ $Y2=0
cc_185 N_A_109_297#_c_281_n N_VPWR_c_312_n 0.00287351f $X=1.065 $Y=1.94 $X2=0
+ $Y2=0
cc_186 N_A_109_297#_c_282_n N_VPWR_c_313_n 0.00540695f $X=1.955 $Y=1.935 $X2=0
+ $Y2=0
cc_187 N_A_109_297#_M1004_d N_VPWR_c_308_n 0.00216833f $X=0.545 $Y=1.485 $X2=0
+ $Y2=0
cc_188 N_A_109_297#_M1006_d N_VPWR_c_308_n 0.00458694f $X=1.905 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_109_297#_c_281_n N_VPWR_c_308_n 0.00506273f $X=1.065 $Y=1.94 $X2=0
+ $Y2=0
cc_190 N_A_109_297#_c_282_n N_VPWR_c_308_n 0.0102394f $X=1.955 $Y=1.935 $X2=0
+ $Y2=0
cc_191 N_VGND_c_353_n A_109_47# 0.00897221f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_192 N_VGND_c_353_n A_381_47# 0.00168632f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

* File: sky130_fd_sc_hd__nand4bb_1.pxi.spice
* Created: Tue Sep  1 19:17:16 2020
* 
x_PM_SKY130_FD_SC_HD__NAND4BB_1%B_N N_B_N_M1011_g N_B_N_M1003_g B_N B_N
+ N_B_N_c_73_n N_B_N_c_74_n N_B_N_c_75_n PM_SKY130_FD_SC_HD__NAND4BB_1%B_N
x_PM_SKY130_FD_SC_HD__NAND4BB_1%D N_D_M1005_g N_D_M1008_g D N_D_c_103_n
+ N_D_c_104_n PM_SKY130_FD_SC_HD__NAND4BB_1%D
x_PM_SKY130_FD_SC_HD__NAND4BB_1%C N_C_M1009_g N_C_M1000_g C C N_C_c_137_n
+ N_C_c_138_n PM_SKY130_FD_SC_HD__NAND4BB_1%C
x_PM_SKY130_FD_SC_HD__NAND4BB_1%A_27_93# N_A_27_93#_M1011_s N_A_27_93#_M1003_s
+ N_A_27_93#_M1007_g N_A_27_93#_M1002_g N_A_27_93#_c_172_n N_A_27_93#_c_186_n
+ N_A_27_93#_c_195_n N_A_27_93#_c_196_n N_A_27_93#_c_173_n N_A_27_93#_c_174_n
+ N_A_27_93#_c_175_n N_A_27_93#_c_181_n N_A_27_93#_c_176_n N_A_27_93#_c_177_n
+ PM_SKY130_FD_SC_HD__NAND4BB_1%A_27_93#
x_PM_SKY130_FD_SC_HD__NAND4BB_1%A_496_21# N_A_496_21#_M1001_d
+ N_A_496_21#_M1010_d N_A_496_21#_c_254_n N_A_496_21#_M1006_g
+ N_A_496_21#_M1004_g N_A_496_21#_c_255_n N_A_496_21#_c_256_n
+ N_A_496_21#_c_257_n N_A_496_21#_c_264_n N_A_496_21#_c_265_n
+ N_A_496_21#_c_266_n N_A_496_21#_c_258_n N_A_496_21#_c_259_n
+ N_A_496_21#_c_268_n PM_SKY130_FD_SC_HD__NAND4BB_1%A_496_21#
x_PM_SKY130_FD_SC_HD__NAND4BB_1%A_N N_A_N_M1001_g N_A_N_M1010_g A_N A_N A_N
+ N_A_N_c_322_n PM_SKY130_FD_SC_HD__NAND4BB_1%A_N
x_PM_SKY130_FD_SC_HD__NAND4BB_1%VPWR N_VPWR_M1003_d N_VPWR_M1000_d
+ N_VPWR_M1004_d N_VPWR_M1010_s N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n VPWR N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_353_n
+ N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n
+ PM_SKY130_FD_SC_HD__NAND4BB_1%VPWR
x_PM_SKY130_FD_SC_HD__NAND4BB_1%Y N_Y_M1006_d N_Y_M1008_d N_Y_M1002_d
+ N_Y_c_411_n N_Y_c_438_n N_Y_c_413_n N_Y_c_442_n Y Y Y Y Y N_Y_c_409_n
+ PM_SKY130_FD_SC_HD__NAND4BB_1%Y
x_PM_SKY130_FD_SC_HD__NAND4BB_1%VGND N_VGND_M1011_d N_VGND_M1001_s
+ N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n VGND
+ N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n N_VGND_c_457_n
+ PM_SKY130_FD_SC_HD__NAND4BB_1%VGND
cc_1 VNB N_B_N_c_73_n 0.026375f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_2 VNB N_B_N_c_74_n 0.00189996f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_3 VNB N_B_N_c_75_n 0.023136f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=0.995
cc_4 VNB D 0.00214691f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_5 VNB N_D_c_103_n 0.023866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_D_c_104_n 0.0203687f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_7 VNB C 7.87809e-19 $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_8 VNB N_C_c_137_n 0.0238372f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_9 VNB N_C_c_138_n 0.0175769f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=0.995
cc_10 VNB N_A_27_93#_c_172_n 0.00835494f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_11 VNB N_A_27_93#_c_173_n 0.00366705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_93#_c_174_n 0.0208034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_93#_c_175_n 0.0222415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_93#_c_176_n 0.0187525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_93#_c_177_n 0.01662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_496_21#_c_254_n 0.0202414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_496_21#_c_255_n 0.00838112f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=0.995
cc_18 VNB N_A_496_21#_c_256_n 0.00734112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_496_21#_c_257_n 0.0341261f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.19
cc_20 VNB N_A_496_21#_c_258_n 0.0375948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_496_21#_c_259_n 0.0121406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_N_M1001_g 0.0390961f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.675
cc_23 VNB A_N 0.0135725f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_24 VNB N_A_N_c_322_n 0.0246449f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_25 VNB N_VPWR_c_353_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB Y 0.00650928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_409_n 0.00710857f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_450_n 0.0104748f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.445
cc_29 VNB N_VGND_c_451_n 0.00832856f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_30 VNB N_VGND_c_452_n 0.0554535f $X=-0.19 $Y=-0.24 $X2=0.562 $Y2=1.325
cc_31 VNB N_VGND_c_453_n 0.00546079f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.16
cc_32 VNB N_VGND_c_454_n 0.0183994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_455_n 0.0183371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_456_n 0.230994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_457_n 0.00583833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_B_N_M1003_g 0.0581483f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_37 VPB N_B_N_c_73_n 0.00667871f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_38 VPB N_B_N_c_74_n 0.00405826f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_39 VPB N_D_M1008_g 0.0216276f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_40 VPB D 0.00303832f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_41 VPB N_D_c_103_n 0.00638136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_C_M1000_g 0.0212784f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_43 VPB C 8.33727e-19 $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.105
cc_44 VPB N_C_c_137_n 0.00505337f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_45 VPB N_A_27_93#_M1002_g 0.0208468f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=1.16
cc_46 VPB N_A_27_93#_c_173_n 0.00133929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_93#_c_174_n 0.00452473f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_93#_c_181_n 0.0190218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_93#_c_176_n 0.0359949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_496_21#_M1004_g 0.0232687f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=1.16
cc_51 VPB N_A_496_21#_c_255_n 5.40718e-19 $X=-0.19 $Y=1.305 $X2=0.562 $Y2=0.995
cc_52 VPB N_A_496_21#_c_256_n 0.00824115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_496_21#_c_257_n 0.0183624f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.19
cc_54 VPB N_A_496_21#_c_264_n 0.0157202f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.53
cc_55 VPB N_A_496_21#_c_265_n 0.00299094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_496_21#_c_266_n 0.0199642f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_496_21#_c_258_n 0.027959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_496_21#_c_268_n 0.0144617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_N_M1010_g 0.0680414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB A_N 0.00718991f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_61 VPB N_A_N_c_322_n 0.00443941f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=1.325
cc_62 VPB N_VPWR_c_354_n 0.00771155f $X=-0.19 $Y=1.305 $X2=0.562 $Y2=0.995
cc_63 VPB N_VPWR_c_355_n 0.00561441f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.19
cc_64 VPB N_VPWR_c_356_n 0.0196034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_357_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_358_n 0.0177718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_359_n 0.0184056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_353_n 0.0439291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_361_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_362_n 0.0194443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_363_n 0.024447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB Y 0.00336441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 N_B_N_M1003_g N_D_M1008_g 0.0232757f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_74 N_B_N_c_73_n D 2.70739e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_N_c_74_n D 0.0183643f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B_N_c_73_n N_D_c_103_n 0.0213919f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_77 N_B_N_c_74_n N_D_c_103_n 0.00733422f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_N_c_75_n N_D_c_104_n 0.0149036f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_N_c_73_n N_A_27_93#_c_172_n 0.0045695f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B_N_c_74_n N_A_27_93#_c_172_n 0.0274682f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B_N_c_75_n N_A_27_93#_c_172_n 0.0101641f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_82 N_B_N_c_75_n N_A_27_93#_c_186_n 4.86756e-19 $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_83 N_B_N_c_75_n N_A_27_93#_c_175_n 0.00902738f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_84 N_B_N_M1003_g N_A_27_93#_c_181_n 0.0075345f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_85 N_B_N_c_74_n N_A_27_93#_c_176_n 0.0438443f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_86 N_B_N_c_75_n N_A_27_93#_c_176_n 0.0273301f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_87 N_B_N_c_74_n N_VPWR_M1003_d 0.00418201f $X=0.595 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_88 N_B_N_M1003_g N_VPWR_c_354_n 0.00897037f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_89 N_B_N_c_73_n N_VPWR_c_354_n 5.2965e-19 $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_N_c_74_n N_VPWR_c_354_n 0.0157054f $X=0.595 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B_N_M1003_g N_VPWR_c_358_n 0.00541359f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_92 N_B_N_M1003_g N_VPWR_c_353_n 0.0108468f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_93 N_B_N_c_75_n N_VGND_c_450_n 0.00411685f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B_N_c_75_n N_VGND_c_454_n 0.00395103f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B_N_c_75_n N_VGND_c_456_n 0.00512902f $X=0.562 $Y=0.995 $X2=0 $Y2=0
cc_96 N_D_M1008_g N_C_M1000_g 0.0104726f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_97 D C 0.0185021f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 N_D_c_103_n C 8.22137e-19 $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_99 N_D_c_104_n C 6.64262e-19 $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_100 D N_C_c_137_n 0.00145882f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_101 N_D_c_103_n N_C_c_137_n 0.02083f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_102 N_D_c_104_n N_C_c_138_n 0.0260674f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_103 D N_A_27_93#_c_172_n 0.0231391f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_104 N_D_c_103_n N_A_27_93#_c_172_n 0.00457738f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_105 N_D_c_104_n N_A_27_93#_c_172_n 0.0139732f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_106 N_D_c_104_n N_A_27_93#_c_186_n 0.00465857f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_107 D N_A_27_93#_c_195_n 0.00167888f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_108 N_D_c_104_n N_A_27_93#_c_196_n 0.00491518f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_109 N_D_c_104_n N_A_27_93#_c_175_n 5.6862e-19 $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_110 N_D_M1008_g N_VPWR_c_354_n 0.00345838f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_111 N_D_M1008_g N_VPWR_c_356_n 0.00585385f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_112 N_D_M1008_g N_VPWR_c_353_n 0.0110469f $X=1.015 $Y=1.985 $X2=0 $Y2=0
cc_113 D N_Y_c_411_n 0.0151807f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_114 N_D_c_103_n N_Y_c_411_n 0.00110539f $X=1.135 $Y=1.16 $X2=0 $Y2=0
cc_115 N_D_c_104_n N_VGND_c_450_n 0.00463453f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_116 N_D_c_104_n N_VGND_c_452_n 0.00432695f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_117 N_D_c_104_n N_VGND_c_456_n 0.00746381f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_118 N_C_M1000_g N_A_27_93#_M1002_g 0.0222819f $X=1.555 $Y=1.985 $X2=0 $Y2=0
cc_119 C N_A_27_93#_c_172_n 0.0108569f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_120 N_C_c_138_n N_A_27_93#_c_172_n 0.00188341f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_121 N_C_c_138_n N_A_27_93#_c_186_n 0.00335427f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_122 C N_A_27_93#_c_195_n 0.0113003f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_123 N_C_c_137_n N_A_27_93#_c_195_n 0.00173005f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_c_138_n N_A_27_93#_c_195_n 0.0128703f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_125 C N_A_27_93#_c_173_n 0.0297189f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_126 N_C_c_137_n N_A_27_93#_c_173_n 0.00201864f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_127 N_C_c_138_n N_A_27_93#_c_173_n 4.48825e-19 $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_128 C N_A_27_93#_c_174_n 3.82383e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_129 N_C_c_137_n N_A_27_93#_c_174_n 0.0205111f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_130 C N_A_27_93#_c_177_n 9.44339e-19 $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_131 N_C_c_138_n N_A_27_93#_c_177_n 0.0311585f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C_M1000_g N_VPWR_c_355_n 0.00323788f $X=1.555 $Y=1.985 $X2=0 $Y2=0
cc_133 N_C_M1000_g N_VPWR_c_356_n 0.00585385f $X=1.555 $Y=1.985 $X2=0 $Y2=0
cc_134 N_C_M1000_g N_VPWR_c_353_n 0.010942f $X=1.555 $Y=1.985 $X2=0 $Y2=0
cc_135 N_C_M1000_g N_Y_c_413_n 0.0139315f $X=1.555 $Y=1.985 $X2=0 $Y2=0
cc_136 C N_Y_c_413_n 0.0145466f $X=1.53 $Y=0.765 $X2=0 $Y2=0
cc_137 N_C_c_137_n N_Y_c_413_n 0.00241891f $X=1.635 $Y=1.16 $X2=0 $Y2=0
cc_138 N_C_c_138_n N_VGND_c_452_n 0.0037981f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C_c_138_n N_VGND_c_456_n 0.00586764f $X=1.625 $Y=0.995 $X2=0 $Y2=0
cc_140 C A_326_47# 0.00188159f $X=1.53 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_141 N_A_27_93#_c_195_n N_A_496_21#_c_254_n 6.94902e-19 $X=1.97 $Y=0.46 $X2=0
+ $Y2=0
cc_142 N_A_27_93#_c_173_n N_A_496_21#_c_254_n 0.00137816f $X=2.115 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_27_93#_c_177_n N_A_496_21#_c_254_n 0.0303834f $X=2.115 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A_27_93#_M1002_g N_A_496_21#_M1004_g 0.00998098f $X=2.055 $Y=1.985
+ $X2=0 $Y2=0
cc_145 N_A_27_93#_c_173_n N_A_496_21#_c_255_n 3.67712e-19 $X=2.115 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_27_93#_c_174_n N_A_496_21#_c_255_n 0.0181638f $X=2.115 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_27_93#_c_176_n N_VPWR_c_354_n 0.00891459f $X=0.255 $Y=2.065 $X2=0
+ $Y2=0
cc_148 N_A_27_93#_M1002_g N_VPWR_c_355_n 0.00323788f $X=2.055 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_27_93#_c_181_n N_VPWR_c_358_n 0.0214784f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_150 N_A_27_93#_M1003_s N_VPWR_c_353_n 0.00209319f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_151 N_A_27_93#_M1002_g N_VPWR_c_353_n 0.0108595f $X=2.055 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A_27_93#_c_181_n N_VPWR_c_353_n 0.0127291f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_153 N_A_27_93#_M1002_g N_VPWR_c_362_n 0.00585385f $X=2.055 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_27_93#_M1002_g N_Y_c_413_n 0.0133199f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_155 N_A_27_93#_c_173_n N_Y_c_413_n 0.0122334f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_27_93#_c_173_n Y 0.00740837f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_27_93#_c_174_n Y 7.20275e-19 $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_27_93#_M1002_g Y 0.00333298f $X=2.055 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_27_93#_c_174_n Y 0.00184632f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_93#_c_195_n N_Y_c_409_n 0.0166939f $X=1.97 $Y=0.46 $X2=0 $Y2=0
cc_161 N_A_27_93#_c_173_n N_Y_c_409_n 0.0607984f $X=2.115 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A_27_93#_c_177_n N_Y_c_409_n 0.0043541f $X=2.115 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_27_93#_c_172_n N_VGND_M1011_d 0.00324813f $X=1.08 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_164 N_A_27_93#_c_172_n N_VGND_c_450_n 0.0220971f $X=1.08 $Y=0.81 $X2=0 $Y2=0
cc_165 N_A_27_93#_c_172_n N_VGND_c_452_n 0.00223349f $X=1.08 $Y=0.81 $X2=0 $Y2=0
cc_166 N_A_27_93#_c_195_n N_VGND_c_452_n 0.033353f $X=1.97 $Y=0.46 $X2=0 $Y2=0
cc_167 N_A_27_93#_c_196_n N_VGND_c_452_n 0.00658159f $X=1.27 $Y=0.46 $X2=0 $Y2=0
cc_168 N_A_27_93#_c_177_n N_VGND_c_452_n 0.0037962f $X=2.115 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_27_93#_c_172_n N_VGND_c_454_n 0.00204328f $X=1.08 $Y=0.81 $X2=0 $Y2=0
cc_170 N_A_27_93#_c_175_n N_VGND_c_454_n 0.00855792f $X=0.26 $Y=0.61 $X2=0 $Y2=0
cc_171 N_A_27_93#_c_172_n N_VGND_c_456_n 0.00970366f $X=1.08 $Y=0.81 $X2=0 $Y2=0
cc_172 N_A_27_93#_c_195_n N_VGND_c_456_n 0.0330472f $X=1.97 $Y=0.46 $X2=0 $Y2=0
cc_173 N_A_27_93#_c_196_n N_VGND_c_456_n 0.00678673f $X=1.27 $Y=0.46 $X2=0 $Y2=0
cc_174 N_A_27_93#_c_175_n N_VGND_c_456_n 0.0111791f $X=0.26 $Y=0.61 $X2=0 $Y2=0
cc_175 N_A_27_93#_c_177_n N_VGND_c_456_n 0.00578073f $X=2.115 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_27_93#_c_172_n A_218_47# 0.00177717f $X=1.08 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_27_93#_c_186_n A_218_47# 0.00191111f $X=1.175 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_178 N_A_27_93#_c_195_n A_218_47# 0.00699751f $X=1.97 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_27_93#_c_196_n A_218_47# 0.00149154f $X=1.27 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_27_93#_c_195_n A_326_47# 0.00974868f $X=1.97 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_27_93#_c_195_n A_426_47# 0.00246129f $X=1.97 $Y=0.46 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_27_93#_c_173_n A_426_47# 0.00285793f $X=2.115 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_183 N_A_496_21#_c_258_n N_A_N_M1001_g 0.0075831f $X=3.932 $Y=1.835 $X2=0
+ $Y2=0
cc_184 N_A_496_21#_c_256_n N_A_N_M1010_g 0.0084326f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_496_21#_c_264_n N_A_N_M1010_g 0.0157863f $X=3.635 $Y=1.92 $X2=0 $Y2=0
cc_186 N_A_496_21#_c_266_n N_A_N_M1010_g 0.0138244f $X=3.8 $Y=2.34 $X2=0 $Y2=0
cc_187 N_A_496_21#_c_258_n N_A_N_M1010_g 0.0090754f $X=3.932 $Y=1.835 $X2=0
+ $Y2=0
cc_188 N_A_496_21#_c_256_n A_N 0.0320257f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_496_21#_c_257_n A_N 0.00240888f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_496_21#_c_264_n A_N 0.0158783f $X=3.635 $Y=1.92 $X2=0 $Y2=0
cc_191 N_A_496_21#_c_258_n A_N 0.0696303f $X=3.932 $Y=1.835 $X2=0 $Y2=0
cc_192 N_A_496_21#_c_259_n A_N 0.0012329f $X=3.932 $Y=0.4 $X2=0 $Y2=0
cc_193 N_A_496_21#_c_256_n N_A_N_c_322_n 4.06462e-19 $X=2.925 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_A_496_21#_c_257_n N_A_N_c_322_n 0.0122476f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_496_21#_c_264_n N_A_N_c_322_n 2.38579e-19 $X=3.635 $Y=1.92 $X2=0
+ $Y2=0
cc_196 N_A_496_21#_c_258_n N_A_N_c_322_n 0.00760283f $X=3.932 $Y=1.835 $X2=0
+ $Y2=0
cc_197 N_A_496_21#_c_259_n N_A_N_c_322_n 0.00158681f $X=3.932 $Y=0.4 $X2=0 $Y2=0
cc_198 N_A_496_21#_c_268_n N_A_N_c_322_n 0.00155347f $X=3.845 $Y=1.92 $X2=0
+ $Y2=0
cc_199 N_A_496_21#_c_256_n N_VPWR_M1004_d 0.00444277f $X=2.925 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_496_21#_c_265_n N_VPWR_M1004_d 0.00308347f $X=3.09 $Y=1.92 $X2=0
+ $Y2=0
cc_201 N_A_496_21#_c_264_n N_VPWR_c_359_n 0.00263605f $X=3.635 $Y=1.92 $X2=0
+ $Y2=0
cc_202 N_A_496_21#_c_266_n N_VPWR_c_359_n 0.0293931f $X=3.8 $Y=2.34 $X2=0 $Y2=0
cc_203 N_A_496_21#_M1010_d N_VPWR_c_353_n 0.0038413f $X=3.57 $Y=2.065 $X2=0
+ $Y2=0
cc_204 N_A_496_21#_M1004_g N_VPWR_c_353_n 0.0120721f $X=2.555 $Y=1.985 $X2=0
+ $Y2=0
cc_205 N_A_496_21#_c_264_n N_VPWR_c_353_n 0.00570629f $X=3.635 $Y=1.92 $X2=0
+ $Y2=0
cc_206 N_A_496_21#_c_265_n N_VPWR_c_353_n 0.0010988f $X=3.09 $Y=1.92 $X2=0 $Y2=0
cc_207 N_A_496_21#_c_266_n N_VPWR_c_353_n 0.0160845f $X=3.8 $Y=2.34 $X2=0 $Y2=0
cc_208 N_A_496_21#_M1004_g N_VPWR_c_362_n 0.00585385f $X=2.555 $Y=1.985 $X2=0
+ $Y2=0
cc_209 N_A_496_21#_M1004_g N_VPWR_c_363_n 0.00483063f $X=2.555 $Y=1.985 $X2=0
+ $Y2=0
cc_210 N_A_496_21#_c_264_n N_VPWR_c_363_n 0.0257452f $X=3.635 $Y=1.92 $X2=0
+ $Y2=0
cc_211 N_A_496_21#_c_265_n N_VPWR_c_363_n 0.0220845f $X=3.09 $Y=1.92 $X2=0 $Y2=0
cc_212 N_A_496_21#_c_266_n N_VPWR_c_363_n 0.0226992f $X=3.8 $Y=2.34 $X2=0 $Y2=0
cc_213 N_A_496_21#_M1004_g Y 0.012632f $X=2.555 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_496_21#_c_254_n Y 0.00503311f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_496_21#_M1004_g Y 0.0058588f $X=2.555 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_496_21#_c_255_n Y 0.00586216f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_496_21#_c_256_n Y 0.0368507f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_496_21#_c_257_n Y 0.00749692f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_496_21#_c_254_n N_Y_c_409_n 0.0129144f $X=2.555 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_496_21#_c_256_n N_Y_c_409_n 0.00765497f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_496_21#_c_257_n N_Y_c_409_n 0.00767749f $X=2.925 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_496_21#_c_254_n N_VGND_c_451_n 0.00244252f $X=2.555 $Y=0.995 $X2=0
+ $Y2=0
cc_223 N_A_496_21#_c_254_n N_VGND_c_452_n 0.00357668f $X=2.555 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_496_21#_c_259_n N_VGND_c_455_n 0.0284384f $X=3.932 $Y=0.4 $X2=0 $Y2=0
cc_225 N_A_496_21#_M1001_d N_VGND_c_456_n 0.00378406f $X=3.57 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_496_21#_c_254_n N_VGND_c_456_n 0.00677056f $X=2.555 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_496_21#_c_259_n N_VGND_c_456_n 0.0163938f $X=3.932 $Y=0.4 $X2=0 $Y2=0
cc_228 N_A_N_M1010_g N_VPWR_c_359_n 0.00348405f $X=3.495 $Y=2.275 $X2=0 $Y2=0
cc_229 N_A_N_M1010_g N_VPWR_c_353_n 0.00525527f $X=3.495 $Y=2.275 $X2=0 $Y2=0
cc_230 N_A_N_M1010_g N_VPWR_c_363_n 0.0110596f $X=3.495 $Y=2.275 $X2=0 $Y2=0
cc_231 N_A_N_M1001_g N_Y_c_409_n 0.005305f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_232 A_N N_Y_c_409_n 0.00423976f $X=3.39 $Y=0.765 $X2=0 $Y2=0
cc_233 N_A_N_M1001_g N_VGND_c_451_n 0.0104027f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_234 A_N N_VGND_c_451_n 0.00338613f $X=3.39 $Y=0.765 $X2=0 $Y2=0
cc_235 N_A_N_M1001_g N_VGND_c_455_n 0.0034938f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_236 A_N N_VGND_c_455_n 0.00261406f $X=3.39 $Y=0.765 $X2=0 $Y2=0
cc_237 N_A_N_M1001_g N_VGND_c_456_n 0.00529027f $X=3.495 $Y=0.445 $X2=0 $Y2=0
cc_238 A_N N_VGND_c_456_n 0.00449455f $X=3.39 $Y=0.765 $X2=0 $Y2=0
cc_239 N_VPWR_c_353_n N_Y_M1008_d 0.00519854f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_240 N_VPWR_c_353_n N_Y_M1002_d 0.00348872f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_241 N_VPWR_c_356_n N_Y_c_438_n 0.0212535f $X=1.64 $Y=2.72 $X2=0 $Y2=0
cc_242 N_VPWR_c_353_n N_Y_c_438_n 0.0126319f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_243 N_VPWR_M1000_d N_Y_c_413_n 0.00920526f $X=1.63 $Y=1.485 $X2=0 $Y2=0
cc_244 N_VPWR_c_355_n N_Y_c_413_n 0.0192006f $X=1.805 $Y=2 $X2=0 $Y2=0
cc_245 N_VPWR_c_353_n N_Y_c_442_n 0.0126214f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_246 N_VPWR_c_362_n N_Y_c_442_n 0.0197903f $X=2.68 $Y=2.49 $X2=0 $Y2=0
cc_247 N_Y_c_409_n N_VGND_c_451_n 0.0250766f $X=2.765 $Y=0.38 $X2=0 $Y2=0
cc_248 N_Y_c_409_n N_VGND_c_452_n 0.0311616f $X=2.765 $Y=0.38 $X2=0 $Y2=0
cc_249 N_Y_M1006_d N_VGND_c_456_n 0.00209319f $X=2.63 $Y=0.235 $X2=0 $Y2=0
cc_250 N_Y_c_409_n N_VGND_c_456_n 0.0187494f $X=2.765 $Y=0.38 $X2=0 $Y2=0
cc_251 Y A_426_47# 5.23065e-19 $X=2.535 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_252 N_Y_c_409_n A_426_47# 0.00576542f $X=2.765 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_253 N_VGND_c_456_n A_218_47# 0.00331341f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_254 N_VGND_c_456_n A_326_47# 0.00297467f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_255 N_VGND_c_456_n A_426_47# 0.0088023f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24

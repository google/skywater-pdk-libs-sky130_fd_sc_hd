* File: sky130_fd_sc_hd__fah_1.pex.spice
* Created: Thu Aug 27 14:21:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__FAH_1%A_67_199# 1 2 9 12 14 18 22 23 27
c61 23 0 3.1734e-19 $X=0.51 $Y=1.16
c62 14 0 1.66784e-19 $X=0.99 $Y=0.82
r63 23 28 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=1.325
r64 23 27 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=0.995
r65 22 25 16.5723 $w=3.46e-07 $l=6.28331e-07 $layer=LI1_cond $X=0.78 $Y=1.16
+ $X2=1.15 $Y2=1.63
r66 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r67 16 18 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.155 $Y=0.735
+ $X2=1.155 $Y2=0.38
r68 15 22 11.9884 $w=3.46e-07 $l=3.4e-07 $layer=LI1_cond $X=0.78 $Y=0.82
+ $X2=0.78 $Y2=1.16
r69 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.99 $Y=0.82
+ $X2=1.155 $Y2=0.735
r70 14 15 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0.82
+ $X2=0.78 $Y2=0.82
r71 12 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.985
+ $X2=0.49 $Y2=1.325
r72 9 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.56 $X2=0.47
+ $Y2=0.995
r73 2 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.485 $X2=1.15 $Y2=1.63
r74 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A 3 5 7 8 10 13 16 17 18 19
c60 19 0 1.70828e-19 $X=1.15 $Y=1.19
c61 16 0 1.66784e-19 $X=0.942 $Y=1.16
c62 5 0 4.97626e-20 $X=0.945 $Y=0.995
r63 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.16 $X2=1.175 $Y2=1.16
r64 17 22 111.037 $w=3.3e-07 $l=6.35e-07 $layer=POLY_cond $X=1.81 $Y=1.16
+ $X2=1.175 $Y2=1.16
r65 17 18 5.03009 $w=3.3e-07 $l=8.2e-08 $layer=POLY_cond $X=1.81 $Y=1.16
+ $X2=1.892 $Y2=1.16
r66 15 22 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=1.175 $Y2=1.16
r67 15 16 5.03009 $w=3.3e-07 $l=7.8e-08 $layer=POLY_cond $X=1.02 $Y=1.16
+ $X2=0.942 $Y2=1.16
r68 11 18 37.0704 $w=1.5e-07 $l=1.68953e-07 $layer=POLY_cond $X=1.9 $Y=1.325
+ $X2=1.892 $Y2=1.16
r69 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.9 $Y=1.325 $X2=1.9
+ $Y2=1.985
r70 8 18 37.0704 $w=1.5e-07 $l=1.68464e-07 $layer=POLY_cond $X=1.885 $Y=0.995
+ $X2=1.892 $Y2=1.16
r71 8 10 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.885 $Y=0.995
+ $X2=1.885 $Y2=0.565
r72 5 16 37.0704 $w=1.5e-07 $l=1.66493e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.942 $Y2=1.16
r73 5 7 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.555
r74 1 16 37.0704 $w=1.5e-07 $l=1.65997e-07 $layer=POLY_cond $X=0.94 $Y=1.325
+ $X2=0.942 $Y2=1.16
r75 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.94 $Y=1.325 $X2=0.94
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%B 3 5 7 8 9 10 12 15 19 21 23 24 29 32 34 35
+ 37 43 54 55 60
c176 55 0 1.1816e-19 $X=5.76 $Y=1.16
c177 54 0 5.3971e-20 $X=5.76 $Y=1.16
c178 29 0 6.36267e-20 $X=2.33 $Y=1.16
c179 19 0 1.516e-19 $X=5.485 $Y=2.03
c180 5 0 2.80009e-19 $X=2.565 $Y=0.995
r181 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.16 $X2=5.76 $Y2=1.16
r182 52 54 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=5.705 $Y=1.16
+ $X2=5.76 $Y2=1.16
r183 50 52 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.485 $Y=1.16
+ $X2=5.705 $Y2=1.16
r184 48 49 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.465 $Y=1.16
+ $X2=2.565 $Y2=1.16
r185 43 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.765 $Y=1.19
+ $X2=5.765 $Y2=1.19
r186 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.22 $Y=1.19
+ $X2=2.075 $Y2=1.19
r187 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.62 $Y=1.19
+ $X2=5.765 $Y2=1.19
r188 34 35 4.20791 $w=1.4e-07 $l=3.4e-06 $layer=MET1_cond $X=5.62 $Y=1.19
+ $X2=2.22 $Y2=1.19
r189 32 60 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.09 $Y=1.19
+ $X2=2.09 $Y2=1.175
r190 32 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.075 $Y=1.19
+ $X2=2.075 $Y2=1.19
r191 30 48 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.33 $Y=1.16
+ $X2=2.465 $Y2=1.16
r192 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.33
+ $Y=1.16 $X2=2.33 $Y2=1.16
r193 27 60 0.716491 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=2.19 $Y=1.175 $X2=2.09
+ $Y2=1.175
r194 27 29 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=2.19 $Y=1.175
+ $X2=2.33 $Y2=1.175
r195 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=0.995
+ $X2=5.705 $Y2=1.16
r196 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.705 $Y=0.995
+ $X2=5.705 $Y2=0.565
r197 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.325
+ $X2=5.485 $Y2=1.16
r198 17 19 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=5.485 $Y=1.325
+ $X2=5.485 $Y2=2.03
r199 13 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.16
r200 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.52 $Y=1.325
+ $X2=3.52 $Y2=1.905
r201 10 24 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.52 $Y2=1.16
r202 10 12 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.52 $Y=0.995
+ $X2=3.52 $Y2=0.555
r203 9 49 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.64 $Y=1.16
+ $X2=2.565 $Y2=1.16
r204 8 24 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.445 $Y=1.16
+ $X2=3.52 $Y2=1.16
r205 8 9 140.763 $w=3.3e-07 $l=8.05e-07 $layer=POLY_cond $X=3.445 $Y=1.16
+ $X2=2.64 $Y2=1.16
r206 5 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=0.995
+ $X2=2.565 $Y2=1.16
r207 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.565 $Y=0.995
+ $X2=2.565 $Y2=0.56
r208 1 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.465 $Y=1.325
+ $X2=2.465 $Y2=1.16
r209 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.465 $Y=1.325
+ $X2=2.465 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_508_297# 1 2 3 4 13 15 18 20 22 25 28 29 30
+ 33 38 39 40 42 44 45 48 50 51 52 53 62 67 75
c204 53 0 9.12361e-20 $X=4.595 $Y=1.53
c205 48 0 7.83819e-20 $X=7.28 $Y=0.68
c206 44 0 3.36117e-19 $X=7.195 $Y=1.01
c207 42 0 1.50384e-19 $X=7.135 $Y=1.955
c208 39 0 1.90878e-20 $X=7.05 $Y=2.04
c209 30 0 1.1816e-19 $X=4.982 $Y=1.16
r210 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.235
+ $Y=1.16 $X2=4.235 $Y2=1.16
r211 63 75 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.235 $Y=1.53
+ $X2=6.375 $Y2=1.53
r212 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.235 $Y=1.53
+ $X2=6.235 $Y2=1.53
r213 60 67 10.1896 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=4.302 $Y=1.53
+ $X2=4.302 $Y2=1.16
r214 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.45 $Y=1.53
+ $X2=4.45 $Y2=1.53
r215 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.535 $Y=1.53
+ $X2=2.535 $Y2=1.53
r216 53 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.595 $Y=1.53
+ $X2=4.45 $Y2=1.53
r217 52 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.09 $Y=1.53
+ $X2=6.235 $Y2=1.53
r218 52 53 1.85024 $w=1.4e-07 $l=1.495e-06 $layer=MET1_cond $X=6.09 $Y=1.53
+ $X2=4.595 $Y2=1.53
r219 51 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.68 $Y=1.53
+ $X2=2.535 $Y2=1.53
r220 50 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.305 $Y=1.53
+ $X2=4.45 $Y2=1.53
r221 50 51 2.01113 $w=1.4e-07 $l=1.625e-06 $layer=MET1_cond $X=4.305 $Y=1.53
+ $X2=2.68 $Y2=1.53
r222 45 56 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.69 $Y=1.58
+ $X2=2.535 $Y2=1.58
r223 43 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.195 $Y=0.765
+ $X2=7.195 $Y2=0.68
r224 43 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.195 $Y=0.765
+ $X2=7.195 $Y2=1.01
r225 41 44 9.58571 $w=2.1e-07 $l=1.92678e-07 $layer=LI1_cond $X=7.135 $Y=1.175
+ $X2=7.195 $Y2=1.01
r226 41 42 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.135 $Y=1.175
+ $X2=7.135 $Y2=1.955
r227 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.05 $Y=2.04
+ $X2=7.135 $Y2=1.955
r228 39 40 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.05 $Y=2.04
+ $X2=6.46 $Y2=2.04
r229 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.955
+ $X2=6.46 $Y2=2.04
r230 36 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.375 $Y=1.955
+ $X2=6.375 $Y2=1.62
r231 35 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=1.615
+ $X2=6.375 $Y2=1.53
r232 35 38 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.375 $Y=1.615
+ $X2=6.375 $Y2=1.62
r233 31 45 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.775 $Y=1.445
+ $X2=2.69 $Y2=1.58
r234 31 33 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.775 $Y=1.445
+ $X2=2.775 $Y2=0.76
r235 29 66 114.534 $w=3.3e-07 $l=6.55e-07 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=4.235 $Y2=1.16
r236 29 30 5.03009 $w=3.3e-07 $l=9.2e-08 $layer=POLY_cond $X=4.89 $Y=1.16
+ $X2=4.982 $Y2=1.16
r237 27 66 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.02 $Y=1.16
+ $X2=4.235 $Y2=1.16
r238 27 28 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.02 $Y=1.16
+ $X2=3.945 $Y2=1.16
r239 23 30 37.0704 $w=1.5e-07 $l=1.73767e-07 $layer=POLY_cond $X=5 $Y=1.325
+ $X2=4.982 $Y2=1.16
r240 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5 $Y=1.325 $X2=5
+ $Y2=1.905
r241 20 30 37.0704 $w=1.5e-07 $l=1.73292e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.982 $Y2=1.16
r242 20 22 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.965 $Y2=0.555
r243 16 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.325
+ $X2=3.945 $Y2=1.16
r244 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.945 $Y=1.325
+ $X2=3.945 $Y2=1.905
r245 13 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=1.16
r246 13 15 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=0.555
r247 4 38 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.485 $X2=6.375 $Y2=1.62
r248 3 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.485 $X2=2.675 $Y2=1.63
r249 2 48 182 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.245 $X2=7.28 $Y2=0.68
r250 1 33 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.235 $X2=2.775 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_719_47# 1 2 9 11 13 14 16 17 18 21 23 24 26
+ 27 29 36 38 39 40 41 44 48 50 51 58
c221 50 0 4.54121e-21 $X=9.005 $Y=0.85
c222 26 0 1.42541e-19 $X=8.88 $Y=0.96
c223 24 0 3.20242e-19 $X=6.615 $Y=1.16
c224 21 0 1.0618e-19 $X=8.955 $Y=1.995
c225 18 0 1.60603e-19 $X=8.525 $Y=1.035
c226 11 0 1.85346e-19 $X=6.645 $Y=0.995
r227 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.27
+ $Y=1.16 $X2=6.27 $Y2=1.16
r228 51 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.12
+ $Y=0.77 $X2=9.12 $Y2=0.77
r229 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.005 $Y=0.85
+ $X2=9.005 $Y2=0.85
r230 48 55 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.27 $Y=0.85
+ $X2=6.27 $Y2=1.16
r231 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.235 $Y=0.85
+ $X2=6.235 $Y2=0.85
r232 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.455 $Y=0.85
+ $X2=3.455 $Y2=0.85
r233 41 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.38 $Y=0.85
+ $X2=6.235 $Y2=0.85
r234 40 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.86 $Y=0.85
+ $X2=9.005 $Y2=0.85
r235 40 41 3.0693 $w=1.4e-07 $l=2.48e-06 $layer=MET1_cond $X=8.86 $Y=0.85
+ $X2=6.38 $Y2=0.85
r236 39 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.6 $Y=0.85
+ $X2=3.455 $Y2=0.85
r237 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.09 $Y=0.85
+ $X2=6.235 $Y2=0.85
r238 38 39 3.08168 $w=1.4e-07 $l=2.49e-06 $layer=MET1_cond $X=6.09 $Y=0.85
+ $X2=3.6 $Y2=0.85
r239 33 44 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.455 $Y=1.455
+ $X2=3.455 $Y2=0.85
r240 32 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.455 $Y=1.62
+ $X2=3.73 $Y2=1.62
r241 32 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.455 $Y=1.62
+ $X2=3.455 $Y2=1.455
r242 31 44 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.455 $Y=0.805
+ $X2=3.455 $Y2=0.85
r243 27 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=0.72
+ $X2=3.455 $Y2=0.805
r244 27 29 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.54 $Y=0.72
+ $X2=3.735 $Y2=0.72
r245 25 58 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=9.12 $Y=0.96
+ $X2=9.12 $Y2=0.77
r246 25 26 15.2969 $w=2.1e-07 $l=2.4e-07 $layer=POLY_cond $X=9.12 $Y=0.96
+ $X2=8.88 $Y2=0.96
r247 23 54 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.51 $Y=1.16
+ $X2=6.27 $Y2=1.16
r248 23 24 5.03009 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.51 $Y=1.16
+ $X2=6.615 $Y2=1.16
r249 19 26 15.2969 $w=2.1e-07 $l=1.83712e-07 $layer=POLY_cond $X=8.955 $Y=1.11
+ $X2=8.88 $Y2=0.96
r250 19 21 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=8.955 $Y=1.11
+ $X2=8.955 $Y2=1.995
r251 17 26 10.1846 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.88 $Y=1.035
+ $X2=8.88 $Y2=0.96
r252 17 18 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=8.88 $Y=1.035
+ $X2=8.525 $Y2=1.035
r253 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.45 $Y=0.96
+ $X2=8.525 $Y2=1.035
r254 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.45 $Y=0.96
+ $X2=8.45 $Y2=0.565
r255 11 24 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.645 $Y=0.995
+ $X2=6.615 $Y2=1.16
r256 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.645 $Y=0.995
+ $X2=6.645 $Y2=0.565
r257 7 24 37.0704 $w=1.5e-07 $l=1.79374e-07 $layer=POLY_cond $X=6.585 $Y=1.325
+ $X2=6.615 $Y2=1.16
r258 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.585 $Y=1.325
+ $X2=6.585 $Y2=1.905
r259 2 36 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.595
+ $Y=1.485 $X2=3.73 $Y2=1.62
r260 1 29 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.235 $X2=3.735 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_1008_47# 1 2 9 11 13 14 16 17 19 21 23 25 30
+ 31 32 33 34 36 37 39 44
c170 30 0 5.3971e-20 $X=5.21 $Y=2.145
r171 42 44 13.1786 $w=1.68e-07 $l=2.02e-07 $layer=LI1_cond $X=5.21 $Y=1.235
+ $X2=5.412 $Y2=1.235
r172 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.535
+ $Y=1.16 $X2=7.535 $Y2=1.16
r173 37 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.535 $Y=1.275
+ $X2=7.535 $Y2=1.16
r174 35 37 8.3945 $w=2.18e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.475 $Y=1.425
+ $X2=7.535 $Y2=1.275
r175 35 36 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.475 $Y=1.425
+ $X2=7.475 $Y2=2.295
r176 34 44 0.22998 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.412 $Y=1.15
+ $X2=5.412 $Y2=1.235
r177 33 47 10.9216 $w=1.85e-07 $l=1.68953e-07 $layer=LI1_cond $X=5.412 $Y=0.925
+ $X2=5.42 $Y2=0.76
r178 33 34 13.4889 $w=1.83e-07 $l=2.25e-07 $layer=LI1_cond $X=5.412 $Y=0.925
+ $X2=5.412 $Y2=1.15
r179 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=2.38
+ $X2=7.475 $Y2=2.295
r180 31 32 136.679 $w=1.68e-07 $l=2.095e-06 $layer=LI1_cond $X=7.39 $Y=2.38
+ $X2=5.295 $Y2=2.38
r181 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.21 $Y=2.295
+ $X2=5.295 $Y2=2.38
r182 28 30 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.21 $Y=2.295
+ $X2=5.21 $Y2=2.145
r183 27 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=1.32
+ $X2=5.21 $Y2=1.235
r184 27 30 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.21 $Y=1.32
+ $X2=5.21 $Y2=2.145
r185 25 40 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=7.935 $Y=1.16
+ $X2=7.535 $Y2=1.16
r186 25 26 62.3073 $w=2.05e-07 $l=2.65e-07 $layer=POLY_cond $X=8.05 $Y=1.16
+ $X2=8.05 $Y2=1.425
r187 22 40 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.145 $Y=1.16
+ $X2=7.535 $Y2=1.16
r188 22 23 5.03009 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=7.145 $Y=1.16
+ $X2=7.037 $Y2=1.16
r189 19 21 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.535 $Y=1.5
+ $X2=8.535 $Y2=1.995
r190 18 26 10.146 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=8.165 $Y=1.425
+ $X2=8.05 $Y2=1.425
r191 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.46 $Y=1.425
+ $X2=8.535 $Y2=1.5
r192 17 18 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=8.46 $Y=1.425
+ $X2=8.165 $Y2=1.425
r193 14 25 42.3552 $w=2.05e-07 $l=1.83916e-07 $layer=POLY_cond $X=8.01 $Y=0.995
+ $X2=8.05 $Y2=1.16
r194 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.01 $Y=0.995
+ $X2=8.01 $Y2=0.565
r195 11 23 37.0704 $w=1.5e-07 $l=1.80748e-07 $layer=POLY_cond $X=7.07 $Y=0.995
+ $X2=7.037 $Y2=1.16
r196 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.07 $Y=0.995
+ $X2=7.07 $Y2=0.565
r197 7 23 37.0704 $w=1.5e-07 $l=1.80291e-07 $layer=POLY_cond $X=7.005 $Y=1.325
+ $X2=7.037 $Y2=1.16
r198 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.005 $Y=1.325
+ $X2=7.005 $Y2=1.905
r199 2 30 600 $w=1.7e-07 $l=7.24362e-07 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=1.485 $X2=5.21 $Y2=2.145
r200 1 47 182 $w=1.7e-07 $l=6.94982e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.435 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%CI 3 6 10 12 13 15 19
c67 19 0 4.54121e-21 $X=9.687 $Y=0.995
c68 12 0 1.0618e-19 $X=9.777 $Y=1.2
c69 10 0 1.69007e-19 $X=9.64 $Y=1.16
r70 15 23 8.20727 $w=1.98e-07 $l=1.48e-07 $layer=LI1_cond $X=9.925 $Y=0.835
+ $X2=9.777 $Y2=0.835
r71 15 23 1.54897 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=9.777 $Y=0.935
+ $X2=9.777 $Y2=0.835
r72 13 15 7.96581 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=9.777 $Y=1.075
+ $X2=9.777 $Y2=0.935
r73 12 13 2.85067 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=9.777 $Y=1.2
+ $X2=9.777 $Y2=1.075
r74 10 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.687 $Y=1.16
+ $X2=9.687 $Y2=1.325
r75 10 19 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.687 $Y=1.16
+ $X2=9.687 $Y2=0.995
r76 9 12 6.31539 $w=2.48e-07 $l=1.37e-07 $layer=LI1_cond $X=9.64 $Y=1.2
+ $X2=9.777 $Y2=1.2
r77 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.64
+ $Y=1.16 $X2=9.64 $Y2=1.16
r78 6 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.795 $Y=1.985
+ $X2=9.795 $Y2=1.325
r79 3 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.78 $Y=0.565
+ $X2=9.78 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_1262_49# 1 2 3 4 5 18 21 23 28 29 32 35 37
+ 38 41 42 43 47 48 50 55 56 57 66
c174 56 0 1.60603e-19 $X=7.832 $Y=0.825
c175 47 0 4.26682e-20 $X=10.265 $Y=1.16
r176 56 57 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=7.875 $Y=0.825
+ $X2=7.875 $Y2=1.51
r177 50 53 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.435 $Y=0.34
+ $X2=6.435 $Y2=0.485
r178 48 67 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=10.277 $Y=1.16
+ $X2=10.277 $Y2=1.325
r179 48 66 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=10.277 $Y=1.16
+ $X2=10.277 $Y2=0.995
r180 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.265
+ $Y=1.16 $X2=10.265 $Y2=1.16
r181 45 47 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.265 $Y=1.495
+ $X2=10.265 $Y2=1.16
r182 44 64 3.62176 $w=2.1e-07 $l=1.18e-07 $layer=LI1_cond $X=9.655 $Y=1.6
+ $X2=9.537 $Y2=1.6
r183 43 45 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=10.18 $Y=1.6
+ $X2=10.265 $Y2=1.495
r184 43 44 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=10.18 $Y=1.6
+ $X2=9.655 $Y2=1.6
r185 41 64 3.22275 $w=2.35e-07 $l=1.05e-07 $layer=LI1_cond $X=9.537 $Y=1.705
+ $X2=9.537 $Y2=1.6
r186 41 42 28.9337 $w=2.33e-07 $l=5.9e-07 $layer=LI1_cond $X=9.537 $Y=1.705
+ $X2=9.537 $Y2=2.295
r187 38 40 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.96 $Y=2.38
+ $X2=9.39 $Y2=2.38
r188 37 42 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=9.42 $Y=2.38
+ $X2=9.537 $Y2=2.295
r189 37 40 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=9.42 $Y=2.38 $X2=9.39
+ $Y2=2.38
r190 36 55 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.96 $Y=0.34
+ $X2=7.832 $Y2=0.34
r191 35 61 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=9.567 $Y=0.34
+ $X2=9.567 $Y2=0.43
r192 35 36 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.4 $Y=0.34
+ $X2=7.96 $Y2=0.34
r193 30 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.845 $Y=2.295
+ $X2=7.96 $Y2=2.38
r194 30 32 31.0659 $w=2.28e-07 $l=6.2e-07 $layer=LI1_cond $X=7.845 $Y=2.295
+ $X2=7.845 $Y2=1.675
r195 29 57 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.845 $Y=1.625
+ $X2=7.845 $Y2=1.51
r196 29 32 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=7.845 $Y=1.625
+ $X2=7.845 $Y2=1.675
r197 26 56 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=7.832 $Y=0.698
+ $X2=7.832 $Y2=0.825
r198 26 28 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=7.832 $Y=0.698
+ $X2=7.832 $Y2=0.66
r199 25 55 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.832 $Y=0.425
+ $X2=7.832 $Y2=0.34
r200 25 28 10.6206 $w=2.53e-07 $l=2.35e-07 $layer=LI1_cond $X=7.832 $Y=0.425
+ $X2=7.832 $Y2=0.66
r201 24 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=0.34
+ $X2=6.435 $Y2=0.34
r202 23 55 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.705 $Y=0.34
+ $X2=7.832 $Y2=0.34
r203 23 24 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=7.705 $Y=0.34
+ $X2=6.6 $Y2=0.34
r204 21 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.215 $Y=1.985
+ $X2=10.215 $Y2=1.325
r205 18 66 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.2 $Y=0.565
+ $X2=10.2 $Y2=0.995
r206 5 64 600 $w=1.7e-07 $l=5.77062e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.575 $X2=9.585 $Y2=1.62
r207 5 40 600 $w=1.7e-07 $l=9.68414e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.575 $X2=9.39 $Y2=2.38
r208 4 32 600 $w=1.7e-07 $l=8.24545e-07 $layer=licon1_PDIFF $count=1 $X=7.08
+ $Y=1.485 $X2=7.815 $Y2=1.675
r209 3 61 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.435
+ $Y=0.245 $X2=9.57 $Y2=0.43
r210 2 28 182 $w=1.7e-07 $l=4.73392e-07 $layer=licon1_NDIFF $count=1 $X=7.675
+ $Y=0.245 $X2=7.8 $Y2=0.66
r211 1 53 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.245 $X2=6.435 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_1332_297# 1 2 9 12 14 15 18 22 23 26 29 33
+ 34 35
c113 22 0 2.20923e-19 $X=11.16 $Y=1.19
c114 18 0 1.67718e-19 $X=6.795 $Y=1.62
r115 33 36 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.325 $Y=1.16
+ $X2=11.325 $Y2=1.325
r116 33 35 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.325 $Y=1.16
+ $X2=11.325 $Y2=0.995
r117 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.295
+ $Y=1.16 $X2=11.295 $Y2=1.16
r118 29 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.305 $Y=1.19
+ $X2=11.305 $Y2=1.19
r119 26 41 5.20126 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=1.19
+ $X2=6.745 $Y2=1.275
r120 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.695 $Y=1.19
+ $X2=6.695 $Y2=1.19
r121 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.84 $Y=1.19
+ $X2=6.695 $Y2=1.19
r122 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.16 $Y=1.19
+ $X2=11.305 $Y2=1.19
r123 22 23 5.34652 $w=1.4e-07 $l=4.32e-06 $layer=MET1_cond $X=11.16 $Y=1.19
+ $X2=6.84 $Y2=1.19
r124 18 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.795 $Y=1.62
+ $X2=6.795 $Y2=1.275
r125 15 26 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=6.745 $Y=1.14
+ $X2=6.745 $Y2=1.19
r126 14 21 7.52707 $w=2.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=6.745 $Y=0.925
+ $X2=6.775 $Y2=0.76
r127 14 15 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.745 $Y=0.925
+ $X2=6.745 $Y2=1.14
r128 12 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.435 $Y=1.985
+ $X2=11.435 $Y2=1.325
r129 9 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.435 $Y=0.56
+ $X2=11.435 $Y2=0.995
r130 2 18 600 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=6.66
+ $Y=1.485 $X2=6.795 $Y2=1.62
r131 1 21 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.245 $X2=6.855 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_1617_49# 1 2 7 9 12 15 17 20 21 22 28 32 33
+ 36
c119 32 0 1.52424e-19 $X=11.855 $Y=1.16
r120 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.855
+ $Y=1.16 $X2=11.855 $Y2=1.16
r121 29 33 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=11.785 $Y=1.53
+ $X2=11.785 $Y2=1.16
r122 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.765 $Y=1.53
+ $X2=11.765 $Y2=1.53
r123 25 36 6.77908 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=8.545 $Y=1.615
+ $X2=8.745 $Y2=1.615
r124 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.545 $Y=1.53
+ $X2=8.545 $Y2=1.53
r125 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.69 $Y=1.53
+ $X2=8.545 $Y2=1.53
r126 21 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.62 $Y=1.53
+ $X2=11.765 $Y2=1.53
r127 21 22 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.62 $Y=1.53
+ $X2=8.69 $Y2=1.53
r128 20 25 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=8.405 $Y=1.615
+ $X2=8.545 $Y2=1.615
r129 17 19 8.52828 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=0.76
+ $X2=8.28 $Y2=0.925
r130 15 20 7.6914 $w=3.4e-07 $l=2.10238e-07 $layer=LI1_cond $X=8.315 $Y=1.445
+ $X2=8.405 $Y2=1.615
r131 15 19 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=8.315 $Y=1.445
+ $X2=8.315 $Y2=0.925
r132 10 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.855 $Y=1.325
+ $X2=11.855 $Y2=1.16
r133 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.855 $Y=1.325
+ $X2=11.855 $Y2=1.985
r134 7 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=11.855 $Y=0.995
+ $X2=11.855 $Y2=1.16
r135 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.855 $Y=0.995
+ $X2=11.855 $Y2=0.56
r136 2 36 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=8.61
+ $Y=1.575 $X2=8.745 $Y2=1.7
r137 1 17 182 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_NDIFF $count=1 $X=8.085
+ $Y=0.245 $X2=8.24 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_27_47# 1 2 3 4 5 6 21 26 29 31 34 35 36 40
+ 42 44 45 46 47 49 50 51 54 58
c168 47 0 4.97626e-20 $X=0.255 $Y=0.805
c169 40 0 1.516e-19 $X=4.79 $Y=2.295
c170 36 0 6.77358e-20 $X=2.805 $Y=2.38
c171 31 0 1.46513e-19 $X=2.635 $Y=1.98
r172 58 61 4.60977 $w=3.48e-07 $l=1.4e-07 $layer=LI1_cond $X=5.925 $Y=0.34
+ $X2=5.925 $Y2=0.48
r173 54 55 17.5519 $w=2.12e-07 $l=3.05e-07 $layer=LI1_cond $X=4.79 $Y=0.785
+ $X2=5.095 $Y2=0.785
r174 53 54 31.9387 $w=2.12e-07 $l=5.55e-07 $layer=LI1_cond $X=4.235 $Y=0.785
+ $X2=4.79 $Y2=0.785
r175 49 50 7.07047 $w=3.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.265 $Y=1.62
+ $X2=0.265 $Y2=1.5
r176 47 50 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.17 $Y=0.805
+ $X2=0.17 $Y2=1.5
r177 45 58 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.925 $Y2=0.34
r178 45 46 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.18 $Y2=0.34
r179 44 55 2.03271 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.095 $Y=0.655
+ $X2=5.095 $Y2=0.785
r180 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.095 $Y=0.425
+ $X2=5.18 $Y2=0.34
r181 43 44 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.095 $Y=0.425
+ $X2=5.095 $Y2=0.655
r182 40 57 3.40825 $w=1.7e-07 $l=1.01833e-07 $layer=LI1_cond $X=4.79 $Y=2.295
+ $X2=4.827 $Y2=2.38
r183 40 42 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.79 $Y=2.295
+ $X2=4.79 $Y2=1.62
r184 39 54 2.03271 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.79 $Y=0.925
+ $X2=4.79 $Y2=0.785
r185 39 42 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.79 $Y=0.925
+ $X2=4.79 $Y2=1.62
r186 36 38 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.805 $Y=2.38
+ $X2=3.23 $Y2=2.38
r187 35 57 3.40825 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=4.827 $Y2=2.38
r188 35 38 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=4.705 $Y=2.38
+ $X2=3.23 $Y2=2.38
r189 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=2.295
+ $X2=2.805 $Y2=2.38
r190 33 34 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.72 $Y=2.065
+ $X2=2.72 $Y2=2.295
r191 32 51 3.86674 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=1.98
+ $X2=0.265 $Y2=1.98
r192 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.635 $Y=1.98
+ $X2=2.72 $Y2=2.065
r193 31 32 142.877 $w=1.68e-07 $l=2.19e-06 $layer=LI1_cond $X=2.635 $Y=1.98
+ $X2=0.445 $Y2=1.98
r194 27 51 2.84813 $w=3.35e-07 $l=9.66954e-08 $layer=LI1_cond $X=0.24 $Y=2.065
+ $X2=0.265 $Y2=1.98
r195 27 29 8.73626 $w=3.08e-07 $l=2.35e-07 $layer=LI1_cond $X=0.24 $Y=2.065
+ $X2=0.24 $Y2=2.3
r196 26 51 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.895
+ $X2=0.265 $Y2=1.98
r197 25 49 1.92074 $w=3.58e-07 $l=6e-08 $layer=LI1_cond $X=0.265 $Y=1.68
+ $X2=0.265 $Y2=1.62
r198 25 26 6.88265 $w=3.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.265 $Y=1.68
+ $X2=0.265 $Y2=1.895
r199 19 47 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.635
+ $X2=0.255 $Y2=0.805
r200 19 21 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=0.255 $Y=0.635
+ $X2=0.255 $Y2=0.38
r201 6 57 600 $w=1.7e-07 $l=9.55458e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.485 $X2=4.725 $Y2=2.38
r202 6 42 600 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.485 $X2=4.79 $Y2=1.62
r203 5 38 600 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=1.485 $X2=3.23 $Y2=2.38
r204 4 49 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r205 4 29 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r206 3 61 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.245 $X2=5.915 $Y2=0.48
r207 2 53 182 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.235 $Y2=0.73
r208 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%VPWR 1 2 3 4 15 19 23 27 29 31 36 41 46 56 57
+ 60 63 66 69
c115 27 0 1.52424e-19 $X=11.645 $Y=1.95
r116 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r117 66 67 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r118 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r119 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 57 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r121 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r122 54 69 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=11.687 $Y2=2.72
r123 54 56 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=12.19 $Y2=2.72
r124 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r125 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r126 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r127 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=9.89 $Y2=2.72
r128 49 52 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r129 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r130 47 66 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=10.175 $Y=2.72
+ $X2=10.007 $Y2=2.72
r131 47 49 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.175 $Y=2.72
+ $X2=10.35 $Y2=2.72
r132 46 69 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.56 $Y=2.72
+ $X2=11.687 $Y2=2.72
r133 46 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.56 $Y=2.72
+ $X2=11.27 $Y2=2.72
r134 45 67 2.09423 $w=4.8e-07 $l=7.36e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=9.89 $Y2=2.72
r135 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 44 45 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r137 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.23 $Y2=2.72
r138 42 44 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 41 66 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=9.84 $Y=2.72
+ $X2=10.007 $Y2=2.72
r140 41 44 476.909 $w=1.68e-07 $l=7.31e-06 $layer=LI1_cond $X=9.84 $Y=2.72
+ $X2=2.53 $Y2=2.72
r141 40 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r142 40 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r143 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r144 37 60 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.747 $Y2=2.72
r145 37 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.15 $Y2=2.72
r146 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.23 $Y2=2.72
r147 36 39 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 31 60 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.747 $Y2=2.72
r149 31 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r150 29 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 25 69 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.687 $Y=2.635
+ $X2=11.687 $Y2=2.72
r153 25 27 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=11.687 $Y=2.635
+ $X2=11.687 $Y2=1.95
r154 21 66 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=10.007 $Y=2.635
+ $X2=10.007 $Y2=2.72
r155 21 23 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=10.007 $Y=2.635
+ $X2=10.007 $Y2=2.36
r156 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.635
+ $X2=2.23 $Y2=2.72
r157 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.23 $Y=2.635
+ $X2=2.23 $Y2=2.32
r158 13 60 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=2.635
+ $X2=0.747 $Y2=2.72
r159 13 15 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.747 $Y=2.635
+ $X2=0.747 $Y2=2.345
r160 4 27 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=11.51
+ $Y=1.485 $X2=11.645 $Y2=1.95
r161 3 23 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=9.87
+ $Y=1.485 $X2=10.005 $Y2=2.36
r162 2 19 600 $w=1.7e-07 $l=9.54018e-07 $layer=licon1_PDIFF $count=1 $X=1.975
+ $Y=1.485 $X2=2.23 $Y2=2.32
r163 1 15 600 $w=1.7e-07 $l=9.38882e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.485 $X2=0.73 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_310_49# 1 2 3 4 5 6 21 24 25 28 29 30 32 33
+ 37 38 41 42 43 48 49 52 55 56
c173 52 0 9.12361e-20 $X=4.07 $Y=1.87
c174 41 0 8.40151e-20 $X=1.5 $Y=0.715
c175 21 0 1.95994e-19 $X=1.675 $Y=0.39
r176 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.655 $Y=1.87
+ $X2=5.655 $Y2=1.87
r177 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=1.87
+ $X2=4.07 $Y2=1.87
r178 49 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.215 $Y=1.87
+ $X2=4.07 $Y2=1.87
r179 48 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.51 $Y=1.87
+ $X2=5.655 $Y2=1.87
r180 48 49 1.60272 $w=1.4e-07 $l=1.295e-06 $layer=MET1_cond $X=5.51 $Y=1.87
+ $X2=4.215 $Y2=1.87
r181 43 46 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=4.745 $Y=0.36
+ $X2=4.745 $Y2=0.42
r182 37 52 5.84822 $w=3.33e-07 $l=1.7e-07 $layer=LI1_cond $X=4.152 $Y=2.04
+ $X2=4.152 $Y2=1.87
r183 37 38 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.985 $Y=2.04
+ $X2=3.2 $Y2=2.04
r184 34 42 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=0.36
+ $X2=3.115 $Y2=0.36
r185 34 36 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=3.2 $Y=0.36
+ $X2=3.31 $Y2=0.36
r186 33 43 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=4.65 $Y=0.36
+ $X2=4.745 $Y2=0.36
r187 33 36 70.7706 $w=2.08e-07 $l=1.34e-06 $layer=LI1_cond $X=4.65 $Y=0.36
+ $X2=3.31 $Y2=0.36
r188 32 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=1.955
+ $X2=3.2 $Y2=2.04
r189 31 42 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.115 $Y=0.465
+ $X2=3.115 $Y2=0.36
r190 31 32 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=3.115 $Y=0.465
+ $X2=3.115 $Y2=1.955
r191 29 42 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.03 $Y=0.34
+ $X2=3.115 $Y2=0.36
r192 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.03 $Y=0.34
+ $X2=2.52 $Y2=0.34
r193 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.52 $Y2=0.34
r194 27 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.435 $Y2=0.715
r195 26 41 3.08518 $w=1.7e-07 $l=3.80132e-07 $layer=LI1_cond $X=1.84 $Y=0.8
+ $X2=1.5 $Y2=0.715
r196 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.35 $Y=0.8
+ $X2=2.435 $Y2=0.715
r197 25 26 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.35 $Y=0.8
+ $X2=1.84 $Y2=0.8
r198 24 40 8.8853 $w=3.46e-07 $l=2.19465e-07 $layer=LI1_cond $X=1.717 $Y=1.445
+ $X2=1.665 $Y2=1.64
r199 23 41 3.43356 $w=2.72e-07 $l=2.97185e-07 $layer=LI1_cond $X=1.717 $Y=0.905
+ $X2=1.5 $Y2=0.715
r200 23 24 29.2151 $w=2.03e-07 $l=5.4e-07 $layer=LI1_cond $X=1.717 $Y=0.905
+ $X2=1.717 $Y2=1.445
r201 19 41 3.43356 $w=2.72e-07 $l=1.7e-07 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.5 $Y2=0.715
r202 19 21 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.39
r203 6 56 600 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.61 $X2=5.695 $Y2=1.865
r204 5 37 600 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.485 $X2=4.155 $Y2=2.04
r205 4 40 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.675 $Y2=1.64
r206 3 46 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.235 $X2=4.755 $Y2=0.42
r207 2 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.235 $X2=3.31 $Y2=0.38
r208 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.245 $X2=1.675 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%A_1640_380# 1 2 3 4 13 19 21 22 23 30 35 36 39
+ 42 43
c116 39 0 1.69007e-19 $X=9.165 $Y=1.87
c117 4 0 4.26682e-20 $X=10.29 $Y=1.485
r118 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.605 $Y=1.87
+ $X2=10.605 $Y2=1.87
r119 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.165 $Y=1.87
+ $X2=9.165 $Y2=1.87
r120 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.31 $Y=1.87
+ $X2=9.165 $Y2=1.87
r121 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.46 $Y=1.87
+ $X2=10.605 $Y2=1.87
r122 35 36 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=10.46 $Y=1.87
+ $X2=9.31 $Y2=1.87
r123 34 43 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=10.605 $Y=1.875
+ $X2=10.605 $Y2=1.87
r124 32 43 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=10.605 $Y=0.825
+ $X2=10.605 $Y2=1.87
r125 30 32 15.5946 $w=4.43e-07 $l=4.25e-07 $layer=LI1_cond $X=10.467 $Y=0.4
+ $X2=10.467 $Y2=0.825
r126 27 39 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=1.955
+ $X2=9.165 $Y2=1.87
r127 26 39 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=9.165 $Y=1.275
+ $X2=9.165 $Y2=1.87
r128 23 34 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=10.517 $Y=2.047
+ $X2=10.517 $Y2=1.875
r129 23 25 0.813333 $w=3.45e-07 $l=2.3e-08 $layer=LI1_cond $X=10.517 $Y=2.047
+ $X2=10.517 $Y2=2.07
r130 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.08 $Y=1.19
+ $X2=9.165 $Y2=1.275
r131 21 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.08 $Y=1.19
+ $X2=8.745 $Y2=1.19
r132 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.66 $Y=1.105
+ $X2=8.745 $Y2=1.19
r133 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.66 $Y=1.105
+ $X2=8.66 $Y2=0.76
r134 13 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.08 $Y=2.04
+ $X2=9.165 $Y2=1.955
r135 13 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=9.08 $Y=2.04
+ $X2=8.325 $Y2=2.04
r136 4 25 600 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=1 $X=10.29
+ $Y=1.485 $X2=10.43 $Y2=2.07
r137 3 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.2
+ $Y=1.9 $X2=8.325 $Y2=2.04
r138 2 30 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.275
+ $Y=0.245 $X2=10.41 $Y2=0.4
r139 1 19 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=8.525
+ $Y=0.245 $X2=8.66 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%COUT 1 2 12 16 17 18 19
r39 19 26 2.41516 $w=5.18e-07 $l=1.05e-07 $layer=LI1_cond $X=11.13 $Y=2.21
+ $X2=11.13 $Y2=2.315
r40 18 19 7.82051 $w=5.18e-07 $l=3.4e-07 $layer=LI1_cond $X=11.13 $Y=1.87
+ $X2=11.13 $Y2=2.21
r41 16 17 9.06626 $w=5.18e-07 $l=1.4e-07 $layer=LI1_cond $X=11.13 $Y=1.635
+ $X2=11.13 $Y2=1.495
r42 14 18 2.64517 $w=5.18e-07 $l=1.15e-07 $layer=LI1_cond $X=11.13 $Y=1.755
+ $X2=11.13 $Y2=1.87
r43 14 16 2.76018 $w=5.18e-07 $l=1.2e-07 $layer=LI1_cond $X=11.13 $Y=1.755
+ $X2=11.13 $Y2=1.635
r44 9 12 5.81876 $w=5.53e-07 $l=2.7e-07 $layer=LI1_cond $X=10.955 $Y=0.547
+ $X2=11.225 $Y2=0.547
r45 7 9 7.81693 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=10.955 $Y=0.825
+ $X2=10.955 $Y2=0.547
r46 7 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.955 $Y=0.825
+ $X2=10.955 $Y2=1.495
r47 2 26 400 $w=1.7e-07 $l=8.90309e-07 $layer=licon1_PDIFF $count=1 $X=11.1
+ $Y=1.485 $X2=11.225 $Y2=2.315
r48 2 16 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=11.1
+ $Y=1.485 $X2=11.225 $Y2=1.635
r49 1 12 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=11.09
+ $Y=0.235 $X2=11.225 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%SUM 1 2 7 8 9 10 11 12 23
r16 12 35 8.23174 $w=3.48e-07 $l=2.5e-07 $layer=LI1_cond $X=12.16 $Y=2.21
+ $X2=12.16 $Y2=1.96
r17 11 35 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=12.16 $Y=1.87
+ $X2=12.16 $Y2=1.96
r18 10 11 9.55671 $w=3.93e-07 $l=2.55e-07 $layer=LI1_cond $X=12.222 $Y=1.53
+ $X2=12.222 $Y2=1.785
r19 9 10 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=12.222 $Y=1.19
+ $X2=12.222 $Y2=1.53
r20 8 39 2.51278 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=12.157 $Y=0.795
+ $X2=12.157 $Y2=0.825
r21 8 21 4.77209 $w=3.53e-07 $l=1.47e-07 $layer=LI1_cond $X=12.157 $Y=0.795
+ $X2=12.157 $Y2=0.648
r22 8 9 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=12.222 $Y=0.88
+ $X2=12.222 $Y2=1.19
r23 8 39 2.81708 $w=2.23e-07 $l=5.5e-08 $layer=LI1_cond $X=12.222 $Y=0.88
+ $X2=12.222 $Y2=0.825
r24 7 21 4.47992 $w=3.53e-07 $l=1.38e-07 $layer=LI1_cond $X=12.157 $Y=0.51
+ $X2=12.157 $Y2=0.648
r25 7 23 3.89558 $w=3.53e-07 $l=1.2e-07 $layer=LI1_cond $X=12.157 $Y=0.51
+ $X2=12.157 $Y2=0.39
r26 2 35 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=11.93
+ $Y=1.485 $X2=12.07 $Y2=1.96
r27 1 23 91 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=2 $X=11.93
+ $Y=0.235 $X2=12.145 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__FAH_1%VGND 1 2 3 4 15 17 21 25 29 32 33 35 36 37 39
+ 58 59 62 65
r135 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r136 63 66 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r137 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r138 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r139 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r140 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r141 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r142 52 55 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r143 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r144 50 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r145 49 50 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r146 47 50 2.09423 $w=4.8e-07 $l=7.36e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=9.89
+ $Y2=0
r147 47 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r148 46 49 480.171 $w=1.68e-07 $l=7.36e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=9.89
+ $Y2=0
r149 46 47 1.09412 $w=1.7e-07 $l=1.445e-06 $layer=mcon $count=8 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r150 44 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.095
+ $Y2=0
r151 44 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.53
+ $Y2=0
r152 39 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.68
+ $Y2=0
r153 39 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r154 37 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r155 37 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r156 35 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.48 $Y=0
+ $X2=11.27 $Y2=0
r157 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=0
+ $X2=11.645 $Y2=0
r158 34 58 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.81 $Y=0
+ $X2=12.19 $Y2=0
r159 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.81 $Y=0
+ $X2=11.645 $Y2=0
r160 32 49 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=9.905 $Y=0 $X2=9.89
+ $Y2=0
r161 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.905 $Y=0 $X2=9.99
+ $Y2=0
r162 31 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.075 $Y=0
+ $X2=10.35 $Y2=0
r163 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.075 $Y=0 $X2=9.99
+ $Y2=0
r164 27 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.645 $Y=0.085
+ $X2=11.645 $Y2=0
r165 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=11.645 $Y=0.085
+ $X2=11.645 $Y2=0.39
r166 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.99 $Y=0.085
+ $X2=9.99 $Y2=0
r167 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.99 $Y=0.085
+ $X2=9.99 $Y2=0.4
r168 19 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r169 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.38
r170 18 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.68
+ $Y2=0
r171 17 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.095
+ $Y2=0
r172 17 18 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=2.01 $Y=0
+ $X2=0.765 $Y2=0
r173 13 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r174 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r175 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=11.51
+ $Y=0.235 $X2=11.645 $Y2=0.39
r176 3 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.855
+ $Y=0.245 $X2=9.99 $Y2=0.4
r177 2 21 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.245 $X2=2.095 $Y2=0.38
r178 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


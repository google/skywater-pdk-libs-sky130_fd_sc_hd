# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.56000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 0.995000 ;
        RECT 0.085000 0.995000 0.665000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.450000 1.075000 15.650000 1.285000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.925000 0.255000  3.255000 0.725000 ;
        RECT  2.925000 0.725000 16.475000 0.905000 ;
        RECT  3.765000 0.255000  4.095000 0.725000 ;
        RECT  4.605000 0.255000  4.935000 0.725000 ;
        RECT  5.445000 0.255000  5.775000 0.725000 ;
        RECT  6.285000 0.255000  6.615000 0.725000 ;
        RECT  7.125000 0.255000  7.455000 0.725000 ;
        RECT  7.965000 0.255000  8.295000 0.725000 ;
        RECT  8.805000 0.255000  9.135000 0.725000 ;
        RECT  9.645000 0.255000  9.975000 0.725000 ;
        RECT  9.685000 1.455000 16.475000 1.625000 ;
        RECT  9.685000 1.625000  9.935000 2.125000 ;
        RECT 10.485000 0.255000 10.815000 0.725000 ;
        RECT 10.525000 1.625000 10.775000 2.125000 ;
        RECT 11.325000 0.255000 11.655000 0.725000 ;
        RECT 11.365000 1.625000 11.615000 2.125000 ;
        RECT 12.165000 0.255000 12.495000 0.725000 ;
        RECT 12.205000 1.625000 12.455000 2.125000 ;
        RECT 13.005000 0.255000 13.335000 0.725000 ;
        RECT 13.045000 1.625000 13.295000 2.125000 ;
        RECT 13.845000 0.255000 14.175000 0.725000 ;
        RECT 13.885000 1.625000 14.135000 2.125000 ;
        RECT 14.685000 0.255000 15.015000 0.725000 ;
        RECT 14.725000 1.625000 14.975000 2.125000 ;
        RECT 15.525000 0.255000 15.855000 0.725000 ;
        RECT 15.565000 1.625000 15.815000 2.125000 ;
        RECT 15.820000 0.905000 16.475000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.560000 0.085000 ;
        RECT  0.485000  0.085000  0.815000 0.825000 ;
        RECT  1.365000  0.085000  1.615000 0.895000 ;
        RECT  2.205000  0.085000  2.755000 0.905000 ;
        RECT  3.425000  0.085000  3.595000 0.555000 ;
        RECT  4.265000  0.085000  4.435000 0.555000 ;
        RECT  5.105000  0.085000  5.275000 0.555000 ;
        RECT  5.945000  0.085000  6.115000 0.555000 ;
        RECT  6.785000  0.085000  6.955000 0.555000 ;
        RECT  7.625000  0.085000  7.795000 0.555000 ;
        RECT  8.465000  0.085000  8.635000 0.555000 ;
        RECT  9.305000  0.085000  9.475000 0.555000 ;
        RECT 10.145000  0.085000 10.315000 0.555000 ;
        RECT 10.985000  0.085000 11.155000 0.555000 ;
        RECT 11.825000  0.085000 11.995000 0.555000 ;
        RECT 12.665000  0.085000 12.835000 0.555000 ;
        RECT 13.505000  0.085000 13.675000 0.555000 ;
        RECT 14.345000  0.085000 14.515000 0.555000 ;
        RECT 15.185000  0.085000 15.355000 0.555000 ;
        RECT 16.025000  0.085000 16.295000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 16.560000 2.805000 ;
        RECT 0.300000 1.495000  0.515000 2.635000 ;
        RECT 1.185000 1.455000  1.355000 2.635000 ;
        RECT 2.025000 1.455000  2.270000 2.635000 ;
        RECT 2.965000 1.835000  3.215000 2.635000 ;
        RECT 3.805000 1.835000  4.055000 2.635000 ;
        RECT 4.645000 1.835000  4.895000 2.635000 ;
        RECT 5.485000 1.835000  5.735000 2.635000 ;
        RECT 6.325000 1.835000  6.575000 2.635000 ;
        RECT 7.165000 1.835000  7.415000 2.635000 ;
        RECT 8.005000 1.835000  8.255000 2.635000 ;
        RECT 8.845000 1.835000  9.095000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.685000 1.495000  1.015000 2.465000 ;
      RECT  0.835000 1.065000  2.035000 1.075000 ;
      RECT  0.835000 1.075000  9.280000 1.285000 ;
      RECT  0.835000 1.285000  1.015000 1.495000 ;
      RECT  0.985000 0.255000  1.195000 1.065000 ;
      RECT  1.525000 1.285000  1.855000 2.465000 ;
      RECT  1.785000 0.255000  2.035000 1.065000 ;
      RECT  2.475000 1.455000  9.515000 1.665000 ;
      RECT  2.475000 1.665000  2.795000 2.465000 ;
      RECT  3.385000 1.665000  3.635000 2.465000 ;
      RECT  4.225000 1.665000  4.475000 2.465000 ;
      RECT  5.065000 1.665000  5.315000 2.465000 ;
      RECT  5.905000 1.665000  6.155000 2.465000 ;
      RECT  6.745000 1.665000  6.995000 2.465000 ;
      RECT  7.585000 1.665000  7.835000 2.465000 ;
      RECT  8.425000 1.665000  8.675000 2.465000 ;
      RECT  9.265000 1.665000  9.515000 2.295000 ;
      RECT  9.265000 2.295000 16.235000 2.465000 ;
      RECT 10.105000 1.795000 10.355000 2.295000 ;
      RECT 10.945000 1.795000 11.195000 2.295000 ;
      RECT 11.785000 1.795000 12.035000 2.295000 ;
      RECT 12.625000 1.795000 12.875000 2.295000 ;
      RECT 13.465000 1.795000 13.715000 2.295000 ;
      RECT 14.305000 1.795000 14.555000 2.295000 ;
      RECT 15.145000 1.795000 15.395000 2.295000 ;
      RECT 15.985000 1.795000 16.235000 2.295000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__xnor3_2 A B C VGND VNB VPB VPWR X
M1000 VPWR a_87_21# X VPB phighvt w=1e+06u l=150000u
+  ad=1.18455e+12p pd=1.043e+07u as=2.7e+11p ps=2.54e+06u
M1001 a_827_297# B VPWR VPB phighvt w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1002 a_87_21# C a_447_49# VNB nshort w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=4.5445e+11p ps=4.02e+06u
M1003 a_827_297# B VGND VNB nshort w=650000u l=150000u
+  ad=1.6515e+11p pd=1.82e+06u as=7.893e+11p ps=7.67e+06u
M1004 X a_87_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1005 a_1198_49# a_933_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=0p ps=0u
M1006 VGND A a_933_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.8275e+11p ps=3.78e+06u
M1007 X a_87_21# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_933_297# a_827_297# a_423_325# VPB phighvt w=840000u l=150000u
+  ad=6.958e+11p pd=5.23e+06u as=5.646e+11p ps=4.74e+06u
M1009 a_1198_49# a_933_297# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=7.77e+11p pd=5.62e+06u as=0p ps=0u
M1010 a_933_297# a_827_297# a_447_49# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_423_325# B a_1198_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_423_325# B a_933_297# VNB nshort w=640000u l=150000u
+  ad=5.881e+11p pd=4.47e+06u as=0p ps=0u
M1013 a_87_21# C a_423_325# VPB phighvt w=840000u l=150000u
+  ad=3.059e+11p pd=2.63e+06u as=0p ps=0u
M1014 VPWR A a_933_297# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_447_49# B a_933_297# VPB phighvt w=840000u l=150000u
+  ad=8.0855e+11p pd=5.34e+06u as=0p ps=0u
M1016 a_1198_49# a_827_297# a_447_49# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_308_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=0p ps=0u
M1018 a_423_325# a_308_93# a_87_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_447_49# a_308_93# a_87_21# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_87_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1198_49# a_827_297# a_423_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_447_49# B a_1198_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_308_93# C VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
.ends

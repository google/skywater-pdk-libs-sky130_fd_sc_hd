# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.440000 1.355000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.255000 1.315000 0.830000 ;
        RECT 1.060000 1.560000 1.315000 2.465000 ;
        RECT 1.145000 0.830000 1.315000 1.560000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.840000 0.085000 ;
      RECT 0.000000  2.635000 1.840000 2.805000 ;
      RECT 0.175000  0.255000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.890000 0.805000 ;
      RECT 0.175000  1.535000 0.890000 1.705000 ;
      RECT 0.175000  1.705000 0.345000 2.465000 ;
      RECT 0.560000  0.085000 0.890000 0.465000 ;
      RECT 0.560000  1.875000 0.890000 2.635000 ;
      RECT 0.720000  0.805000 0.890000 0.995000 ;
      RECT 0.720000  0.995000 0.975000 1.325000 ;
      RECT 0.720000  1.325000 0.890000 1.535000 ;
      RECT 1.490000  0.085000 1.750000 0.925000 ;
      RECT 1.490000  1.485000 1.750000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
  END
END sky130_fd_sc_hd__buf_2

* File: sky130_fd_sc_hd__dlclkp_2.pex.spice
* Created: Tue Sep  1 19:04:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%CLK 4 5 7 8 10 13 17 21 25 27 29 30 33 36
+ 37 40 42 45
c134 37 0 1.03964e-19 $X=5.295 $Y=1.19
c135 33 0 6.03778e-20 $X=0.235 $Y=1.19
c136 21 0 9.76047e-20 $X=0.47 $Y=0.805
r137 45 48 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.27
+ $X2=5.375 $Y2=1.435
r138 45 47 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.27
+ $X2=5.375 $Y2=1.105
r139 40 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r140 40 42 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r141 37 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.32
+ $Y=1.27 $X2=5.32 $Y2=1.27
r142 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.295 $Y=1.19
+ $X2=5.295 $Y2=1.19
r143 33 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r144 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.235 $Y=1.19
+ $X2=0.235 $Y2=1.19
r145 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.38 $Y=1.19
+ $X2=0.235 $Y2=1.19
r146 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.15 $Y=1.19
+ $X2=5.295 $Y2=1.19
r147 29 30 5.90345 $w=1.4e-07 $l=4.77e-06 $layer=MET1_cond $X=5.15 $Y=1.19
+ $X2=0.38 $Y2=1.19
r148 27 33 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.21 $Y=1.53
+ $X2=0.21 $Y2=1.19
r149 23 25 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r150 19 21 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r151 17 48 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.49 $Y=2.165
+ $X2=5.49 $Y2=1.435
r152 13 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.49 $Y=0.445
+ $X2=5.49 $Y2=1.105
r153 8 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=1.665
r154 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r155 5 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.47 $Y2=0.805
r156 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r157 4 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r158 4 43 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r159 1 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r160 1 42 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%GATE 1 3 5 7 10 11 17
r44 16 17 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.77 $Y=1.56
+ $X2=1.985 $Y2=1.56
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.52 $X2=1.77 $Y2=1.52
r46 11 17 3.27362 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=2.1 $Y=1.56
+ $X2=1.985 $Y2=1.56
r47 10 16 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.615 $Y=1.56
+ $X2=1.77 $Y2=1.56
r48 5 15 94.1973 $w=2.36e-07 $l=4.77389e-07 $layer=POLY_cond $X=1.91 $Y=1.09
+ $X2=1.81 $Y2=1.52
r49 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.91 $Y=1.09 $X2=1.91
+ $Y2=0.805
r50 1 15 40.0744 $w=2.36e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.83 $Y=1.685
+ $X2=1.81 $Y2=1.52
r51 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.83 $Y=1.685 $X2=1.83
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%A_193_47# 1 2 9 13 17 21 26 27 28 30 34 41
c94 30 0 2.0302e-19 $X=3.06 $Y=0.9
c95 21 0 4.39096e-20 $X=2.395 $Y=1.94
c96 17 0 7.04924e-20 $X=1.1 $Y=0.425
r97 31 41 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=3.06 $Y=0.9
+ $X2=3.185 $Y2=0.9
r98 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=0.9 $X2=3.06 $Y2=0.9
r99 28 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.645 $Y=0.9
+ $X2=3.06 $Y2=0.9
r100 27 35 37.7695 $w=2.7e-07 $l=1.7e-07 $layer=POLY_cond $X=2.48 $Y=1.74
+ $X2=2.31 $Y2=1.74
r101 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.74 $X2=2.48 $Y2=1.74
r102 24 26 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.52 $Y=1.855
+ $X2=2.52 $Y2=1.74
r103 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.52 $Y=0.985
+ $X2=2.645 $Y2=0.9
r104 23 26 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=2.52 $Y=0.985
+ $X2=2.52 $Y2=1.74
r105 22 34 2.68609 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.28 $Y=1.94
+ $X2=1.147 $Y2=1.94
r106 21 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.395 $Y=1.94
+ $X2=2.52 $Y2=1.855
r107 21 22 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.395 $Y=1.94
+ $X2=1.28 $Y2=1.94
r108 15 34 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.147 $Y=1.855
+ $X2=1.147 $Y2=1.94
r109 15 17 62.1884 $w=2.63e-07 $l=1.43e-06 $layer=LI1_cond $X=1.147 $Y=1.855
+ $X2=1.147 $Y2=0.425
r110 11 41 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.185 $Y=0.765
+ $X2=3.185 $Y2=0.9
r111 11 13 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.185 $Y=0.765
+ $X2=3.185 $Y2=0.43
r112 7 35 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.31 $Y=1.875
+ $X2=2.31 $Y2=1.74
r113 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.31 $Y=1.875 $X2=2.31
+ $Y2=2.275
r114 2 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r115 1 17 182 $w=1.7e-07 $l=2.48495e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%A_27_47# 1 2 7 9 11 14 16 19 20 21 25 26 27
+ 30 32 35 39 40 41 46 48 50 52 56
c134 27 0 4.39096e-20 $X=2.535 $Y=1.32
c135 14 0 2.69707e-20 $X=0.89 $Y=2.135
c136 11 0 3.34071e-20 $X=0.89 $Y=1.09
r137 51 56 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.225
+ $X2=0.89 $Y2=1.225
r138 50 53 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.225
+ $X2=0.725 $Y2=1.39
r139 50 52 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.225
+ $X2=0.725 $Y2=1.06
r140 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.225 $X2=0.755 $Y2=1.225
r141 46 53 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.39
r142 43 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.695 $Y=0.785
+ $X2=0.695 $Y2=1.06
r143 42 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r144 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r145 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r146 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.7
+ $X2=0.695 $Y2=0.785
r147 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.7
+ $X2=0.345 $Y2=0.7
r148 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.345 $Y2=0.7
r149 33 35 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.425
r150 28 30 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.93 $Y=1.395
+ $X2=2.93 $Y2=2.275
r151 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.855 $Y=1.32
+ $X2=2.93 $Y2=1.395
r152 26 27 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.855 $Y=1.32
+ $X2=2.535 $Y2=1.32
r153 23 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.46 $Y=1.245
+ $X2=2.535 $Y2=1.32
r154 23 25 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.46 $Y=1.245
+ $X2=2.46 $Y2=0.54
r155 22 25 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.46 $Y=0.255
+ $X2=2.46 $Y2=0.54
r156 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.385 $Y=0.18
+ $X2=2.46 $Y2=0.255
r157 20 21 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=2.385 $Y=0.18
+ $X2=1.45 $Y2=0.18
r158 18 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.375 $Y=0.255
+ $X2=1.45 $Y2=0.18
r159 18 19 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.375 $Y=0.255
+ $X2=1.375 $Y2=0.73
r160 17 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=0.805
+ $X2=0.89 $Y2=0.805
r161 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.3 $Y=0.805
+ $X2=1.375 $Y2=0.73
r162 16 17 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.3 $Y=0.805
+ $X2=0.965 $Y2=0.805
r163 12 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.36
+ $X2=0.89 $Y2=1.225
r164 12 14 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=0.89 $Y=1.36
+ $X2=0.89 $Y2=2.135
r165 11 56 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.09
+ $X2=0.89 $Y2=1.225
r166 10 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.88
+ $X2=0.89 $Y2=0.805
r167 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=0.88
+ $X2=0.89 $Y2=1.09
r168 7 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.73
+ $X2=0.89 $Y2=0.805
r169 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.89 $Y=0.73 $X2=0.89
+ $Y2=0.445
r170 2 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r171 1 35 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%A_643_307# 1 2 9 13 15 17 19 21 23 24 31 36
+ 39 42 46 48 52
c111 52 0 7.10306e-21 $X=3.66 $Y=1.7
c112 13 0 1.95917e-19 $X=3.66 $Y=0.445
r113 47 54 79.2176 $w=2.16e-07 $l=3.55e-07 $layer=POLY_cond $X=4.65 $Y=1.16
+ $X2=4.65 $Y2=0.805
r114 46 48 6.67615 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.542 $Y=1.16
+ $X2=4.542 $Y2=0.995
r115 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=1.16 $X2=4.65 $Y2=1.16
r116 44 48 18.6352 $w=2.33e-07 $l=3.8e-07 $layer=LI1_cond $X=4.467 $Y=0.615
+ $X2=4.467 $Y2=0.995
r117 42 44 7.26708 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.45 $Y=0.45
+ $X2=4.45 $Y2=0.615
r118 38 39 0.196141 $w=3.11e-07 $l=5e-09 $layer=LI1_cond $X=4.02 $Y=1.7
+ $X2=4.025 $Y2=1.7
r119 36 39 20.281 $w=3.11e-07 $l=5.17e-07 $layer=LI1_cond $X=4.542 $Y=1.7
+ $X2=4.025 $Y2=1.7
r120 35 46 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=4.542 $Y=1.187
+ $X2=4.542 $Y2=1.16
r121 35 36 10.4169 $w=3.83e-07 $l=3.48e-07 $layer=LI1_cond $X=4.542 $Y=1.187
+ $X2=4.542 $Y2=1.535
r122 29 39 2.76503 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=1.865
+ $X2=4.025 $Y2=1.7
r123 29 31 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.025 $Y=1.865
+ $X2=4.025 $Y2=2.27
r124 27 52 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.52 $Y=1.7
+ $X2=3.66 $Y2=1.7
r125 27 49 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.52 $Y=1.7
+ $X2=3.29 $Y2=1.7
r126 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.52
+ $Y=1.7 $X2=3.52 $Y2=1.7
r127 24 38 3.93671 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=3.915 $Y=1.7
+ $X2=4.02 $Y2=1.7
r128 24 26 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.915 $Y=1.7
+ $X2=3.52 $Y2=1.7
r129 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.13 $Y=0.73
+ $X2=5.13 $Y2=0.445
r130 20 54 11.3495 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.785 $Y=0.805
+ $X2=4.65 $Y2=0.805
r131 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.055 $Y=0.805
+ $X2=5.13 $Y2=0.73
r132 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.055 $Y=0.805
+ $X2=4.785 $Y2=0.805
r133 15 47 41.3672 $w=2.16e-07 $l=1.92678e-07 $layer=POLY_cond $X=4.71 $Y=1.325
+ $X2=4.65 $Y2=1.16
r134 15 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.71 $Y=1.325
+ $X2=4.71 $Y2=2.165
r135 11 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.535
+ $X2=3.66 $Y2=1.7
r136 11 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.66 $Y=1.535
+ $X2=3.66 $Y2=0.445
r137 7 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.29 $Y=1.865
+ $X2=3.29 $Y2=1.7
r138 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.29 $Y=1.865
+ $X2=3.29 $Y2=2.275
r139 2 38 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.02 $Y2=1.755
r140 2 31 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.02 $Y2=2.27
r141 1 42 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.235 $X2=4.4 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%A_477_413# 1 2 9 12 14 18 23 24 25 27 30 31
+ 33 35
r90 31 36 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.132 $Y=1.16
+ $X2=4.132 $Y2=1.325
r91 31 35 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=4.132 $Y=1.16
+ $X2=4.132 $Y2=0.995
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.16 $X2=4.095 $Y2=1.16
r93 28 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=1.16
+ $X2=3.64 $Y2=1.16
r94 28 30 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.725 $Y=1.16
+ $X2=4.095 $Y2=1.16
r95 27 33 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=1.16
r96 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.64 $Y=0.56
+ $X2=3.64 $Y2=0.995
r97 24 33 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.555 $Y=1.24
+ $X2=3.64 $Y2=1.16
r98 24 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.555 $Y=1.24
+ $X2=3.23 $Y2=1.24
r99 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.145 $Y=1.325
+ $X2=3.23 $Y2=1.24
r100 22 23 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.145 $Y=1.325
+ $X2=3.145 $Y2=2.255
r101 18 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.555 $Y=0.475
+ $X2=3.64 $Y2=0.56
r102 18 20 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.555 $Y=0.475
+ $X2=2.96 $Y2=0.475
r103 14 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=2.34
+ $X2=3.145 $Y2=2.255
r104 14 16 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.06 $Y=2.34
+ $X2=2.645 $Y2=2.34
r105 12 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.23 $Y=1.985
+ $X2=4.23 $Y2=1.325
r106 9 35 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.19 $Y=0.56
+ $X2=4.19 $Y2=0.995
r107 2 16 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=2.065 $X2=2.645 $Y2=2.34
r108 1 20 182 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.33 $X2=2.96 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%A_957_369# 1 2 7 9 12 14 16 19 22 25 27 28
+ 29 30 34 37 39 42 46
c93 42 0 1.42073e-19 $X=5.875 $Y=1.325
c94 12 0 1.03964e-19 $X=5.97 $Y=1.985
r95 45 46 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.97 $Y=1.16
+ $X2=6.39 $Y2=1.16
r96 39 41 7.09737 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.992 $Y=0.455
+ $X2=4.992 $Y2=0.62
r97 37 42 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.84 $Y=1.725 $X2=5.84
+ $Y2=1.325
r98 35 45 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.91 $Y=1.16 $X2=5.97
+ $Y2=1.16
r99 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.91
+ $Y=1.16 $X2=5.91 $Y2=1.16
r100 32 42 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=5.875 $Y=1.205
+ $X2=5.875 $Y2=1.325
r101 32 34 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=5.875 $Y=1.205
+ $X2=5.875 $Y2=1.16
r102 31 34 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=5.875 $Y=0.935
+ $X2=5.875 $Y2=1.16
r103 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.755 $Y=1.81
+ $X2=5.84 $Y2=1.725
r104 29 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.755 $Y=1.81
+ $X2=5.34 $Y2=1.81
r105 27 31 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=5.755 $Y=0.85
+ $X2=5.875 $Y2=0.935
r106 27 28 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.755 $Y=0.85
+ $X2=5.15 $Y2=0.85
r107 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.175 $Y=1.895
+ $X2=5.34 $Y2=1.81
r108 23 25 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.175 $Y=1.895
+ $X2=5.175 $Y2=2
r109 22 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.04 $Y=0.765
+ $X2=5.15 $Y2=0.85
r110 22 41 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=5.04 $Y=0.765
+ $X2=5.04 $Y2=0.62
r111 17 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.39 $Y=1.325
+ $X2=6.39 $Y2=1.16
r112 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.39 $Y=1.325
+ $X2=6.39 $Y2=1.985
r113 14 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.39 $Y=0.995
+ $X2=6.39 $Y2=1.16
r114 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.39 $Y=0.995
+ $X2=6.39 $Y2=0.56
r115 10 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.16
r116 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.325
+ $X2=5.97 $Y2=1.985
r117 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=1.16
r118 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=0.56
r119 2 25 300 $w=1.7e-07 $l=4.61031e-07 $layer=licon1_PDIFF $count=2 $X=4.785
+ $Y=1.845 $X2=5.175 $Y2=2
r120 1 39 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=4.795
+ $Y=0.235 $X2=4.92 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 41 43 47
+ 49 54 59 64 69 75 78 81 84 87 91
r100 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r101 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r105 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r106 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 73 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r108 73 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r110 70 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r111 70 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=6.21 $Y2=2.72
r112 69 90 4.32257 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.53 $Y=2.72
+ $X2=6.715 $Y2=2.72
r113 69 72 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.53 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 68 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 68 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r116 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 65 84 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.6 $Y=2.72
+ $X2=4.457 $Y2=2.72
r118 65 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.6 $Y=2.72 $X2=5.29
+ $Y2=2.72
r119 64 87 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.575 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 64 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.575 $Y=2.72
+ $X2=5.29 $Y2=2.72
r121 63 82 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r122 63 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 60 78 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.82 $Y=2.72
+ $X2=1.637 $Y2=2.72
r125 60 62 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.82 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 59 81 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.4 $Y=2.72 $X2=3.55
+ $Y2=2.72
r127 59 62 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.4 $Y=2.72
+ $X2=2.07 $Y2=2.72
r128 58 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r129 58 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r130 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 55 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r132 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 54 78 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.637 $Y2=2.72
r134 54 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r135 49 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r136 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r137 47 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r139 43 46 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.67 $Y=1.66
+ $X2=6.67 $Y2=2.34
r140 41 90 3.03748 $w=2.8e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.67 $Y=2.635
+ $X2=6.715 $Y2=2.72
r141 41 46 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=6.67 $Y=2.635
+ $X2=6.67 $Y2=2.34
r142 37 87 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.75 $Y=2.635
+ $X2=5.75 $Y2=2.72
r143 37 39 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.75 $Y=2.635
+ $X2=5.75 $Y2=2.295
r144 33 84 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.457 $Y=2.635
+ $X2=4.457 $Y2=2.72
r145 33 35 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.457 $Y=2.635
+ $X2=4.457 $Y2=2.27
r146 32 81 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.55
+ $Y2=2.72
r147 31 84 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.315 $Y=2.72
+ $X2=4.457 $Y2=2.72
r148 31 32 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.315 $Y=2.72
+ $X2=3.7 $Y2=2.72
r149 27 81 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r150 27 29 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.3
r151 23 78 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.637 $Y=2.635
+ $X2=1.637 $Y2=2.72
r152 23 25 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.637 $Y=2.635
+ $X2=1.637 $Y2=2.34
r153 19 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r154 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r155 6 46 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=1.485 $X2=6.63 $Y2=2.34
r156 6 43 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=1.485 $X2=6.63 $Y2=1.66
r157 5 39 600 $w=1.7e-07 $l=5.38749e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.845 $X2=5.76 $Y2=2.295
r158 4 35 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.485 $X2=4.44 $Y2=2.27
r159 3 29 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.065 $X2=3.5 $Y2=2.3
r160 2 25 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=2.34
r161 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%GCLK 1 2 8 9 10 11 12 18 31
r24 11 12 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=6.227 $Y=1.87
+ $X2=6.227 $Y2=2.21
r25 11 18 9.13257 $w=2.63e-07 $l=2.1e-07 $layer=LI1_cond $X=6.227 $Y=1.87
+ $X2=6.227 $Y2=1.66
r26 10 31 1.59308 $w=3.38e-07 $l=4.7e-08 $layer=LI1_cond $X=6.215 $Y=0.425
+ $X2=6.262 $Y2=0.425
r27 10 31 4.00821 $w=1.95e-07 $l=1.7e-07 $layer=LI1_cond $X=6.262 $Y=0.595
+ $X2=6.262 $Y2=0.425
r28 10 27 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=6.215 $Y=0.425
+ $X2=6.18 $Y2=0.425
r29 9 10 32.6659 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=6.262 $Y=1.495
+ $X2=6.262 $Y2=0.595
r30 8 18 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=6.227 $Y=1.627
+ $X2=6.227 $Y2=1.66
r31 8 9 6.56726 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=6.227 $Y=1.627
+ $X2=6.227 $Y2=1.495
r32 2 18 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.485 $X2=6.18 $Y2=1.66
r33 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__DLCLKP_2%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43
+ 48 53 58 64 67 70 73 77
c105 77 0 2.71124e-20 $X=6.67 $Y=0
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r107 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r108 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r109 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r110 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r111 62 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r112 62 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r113 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r114 59 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.76
+ $Y2=0
r115 59 61 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=6.21 $Y2=0
r116 58 76 4.32257 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.53 $Y=0 $X2=6.715
+ $Y2=0
r117 58 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.53 $Y=0 $X2=6.21
+ $Y2=0
r118 57 74 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r119 57 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r120 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r121 54 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.02
+ $Y2=0
r122 54 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=4.37 $Y2=0
r123 53 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=0 $X2=5.76
+ $Y2=0
r124 53 56 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=5.675 $Y=0
+ $X2=4.37 $Y2=0
r125 52 71 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.91 $Y2=0
r126 52 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r127 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r128 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.65
+ $Y2=0
r129 49 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.815 $Y=0
+ $X2=2.07 $Y2=0
r130 48 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.02
+ $Y2=0
r131 48 51 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=2.07 $Y2=0
r132 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r133 47 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r134 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r135 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r136 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r137 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.65
+ $Y2=0
r138 43 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.485 $Y=0
+ $X2=1.15 $Y2=0
r139 38 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r140 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r141 36 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r142 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r143 32 76 3.03748 $w=2.8e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.67 $Y=0.085
+ $X2=6.715 $Y2=0
r144 32 34 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=6.67 $Y=0.085
+ $X2=6.67 $Y2=0.38
r145 28 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=0.085
+ $X2=5.76 $Y2=0
r146 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.76 $Y=0.085
+ $X2=5.76 $Y2=0.38
r147 24 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r148 24 26 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.445
r149 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0
r150 20 22 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0.74
r151 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r152 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.36
r153 5 34 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=6.465
+ $Y=0.235 $X2=6.63 $Y2=0.38
r154 4 30 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=5.565
+ $Y=0.235 $X2=5.76 $Y2=0.38
r155 3 26 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.235 $X2=3.98 $Y2=0.445
r156 2 22 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.525
+ $Y=0.595 $X2=1.65 $Y2=0.74
r157 1 18 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends


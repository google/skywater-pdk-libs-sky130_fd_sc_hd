* File: sky130_fd_sc_hd__dfstp_4.pex.spice
* Created: Thu Aug 27 14:15:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DFSTP_4%CLK 4 5 7 8 10 13 17 19 20 24 26
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r46 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r47 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_27_47# 1 2 9 13 15 17 20 24 28 31 35 36 37
+ 40 42 46 47 50 51 52 54 55 59 61 62 63 64 73 78 85 86 92 93 96
c273 92 0 3.16068e-19 $X=5.155 $Y=1.74
c274 86 0 3.30612e-20 $X=2.765 $Y=1.74
c275 85 0 2.53448e-20 $X=2.765 $Y=1.74
c276 73 0 1.73859e-19 $X=5.29 $Y=1.87
c277 63 0 1.39518e-19 $X=5.145 $Y=1.87
c278 61 0 1.01003e-19 $X=2.385 $Y=1.87
c279 52 0 3.12358e-20 $X=5.05 $Y=0.81
c280 51 0 1.753e-19 $X=5.82 $Y=0.81
c281 47 0 9.52104e-20 $X=2.435 $Y=0.87
c282 46 0 1.76471e-19 $X=2.435 $Y=0.87
c283 40 0 1.81794e-19 $X=0.725 $Y=1.795
c284 37 0 3.29888e-20 $X=0.61 $Y=1.88
c285 24 0 7.39505e-20 $X=5.065 $Y=2.275
r286 93 104 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.155 $Y=1.81
+ $X2=4.965 $Y2=1.81
r287 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.155
+ $Y=1.74 $X2=5.155 $Y2=1.74
r288 89 92 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.065 $Y=1.74
+ $X2=5.155 $Y2=1.74
r289 85 88 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.765 $Y=1.74
+ $X2=2.765 $Y2=1.875
r290 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.74 $X2=2.765 $Y2=1.74
r291 73 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r292 71 86 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.765 $Y2=1.765
r293 71 99 2.12292 $w=3.78e-07 $l=7e-08 $layer=LI1_cond $X=2.53 $Y=1.765
+ $X2=2.46 $Y2=1.765
r294 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r295 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.7 $Y=1.87 $X2=0.7
+ $Y2=1.87
r296 64 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.675 $Y=1.87
+ $X2=2.53 $Y2=1.87
r297 63 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r298 63 64 3.05692 $w=1.4e-07 $l=2.47e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=2.675 $Y2=1.87
r299 62 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.845 $Y=1.87
+ $X2=0.7 $Y2=1.87
r300 61 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r301 61 62 1.90594 $w=1.4e-07 $l=1.54e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=0.845 $Y2=1.87
r302 59 96 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.985 $Y=0.93
+ $X2=5.985 $Y2=0.765
r303 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=0.93 $X2=5.985 $Y2=0.93
r304 55 58 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.985 $Y=0.81
+ $X2=5.985 $Y2=0.93
r305 51 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.985 $Y2=0.81
r306 51 52 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.82 $Y=0.81
+ $X2=5.05 $Y2=0.81
r307 50 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.965 $Y=1.655
+ $X2=4.965 $Y2=1.81
r308 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.965 $Y=0.895
+ $X2=5.05 $Y2=0.81
r309 49 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.965 $Y=0.895
+ $X2=4.965 $Y2=1.655
r310 47 80 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.435 $Y=0.87
+ $X2=2.305 $Y2=0.87
r311 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=0.87 $X2=2.435 $Y2=0.87
r312 44 99 3.93508 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=1.765
r313 44 46 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=2.46 $Y=1.575
+ $X2=2.46 $Y2=0.87
r314 43 78 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r315 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r316 40 67 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.88
r317 40 42 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.725 $Y=1.795
+ $X2=0.725 $Y2=1.235
r318 39 42 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=0.805
+ $X2=0.725 $Y2=1.235
r319 38 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r320 37 67 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.725 $Y2=1.88
r321 37 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r322 35 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.725 $Y2=0.805
r323 35 36 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r324 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r325 29 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r326 28 96 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.045 $Y=0.445
+ $X2=6.045 $Y2=0.765
r327 22 89 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=1.74
r328 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.065 $Y=1.875
+ $X2=5.065 $Y2=2.275
r329 20 88 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.735 $Y=2.275
+ $X2=2.735 $Y2=1.875
r330 15 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.87
r331 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.305 $Y=0.705
+ $X2=2.305 $Y2=0.415
r332 11 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r333 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r334 7 78 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r335 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r336 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r337 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%D 3 7 9 10 14 15
c39 14 0 1.34441e-19 $X=1.855 $Y=1.17
c40 7 0 1.76471e-19 $X=1.83 $Y=2.065
r41 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.335
r42 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.17
+ $X2=1.855 $Y2=1.005
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.855
+ $Y=1.17 $X2=1.855 $Y2=1.17
r44 9 10 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.53
r45 9 15 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=1.975 $Y=1.19
+ $X2=1.975 $Y2=1.17
r46 7 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.83 $Y=2.065
+ $X2=1.83 $Y2=1.335
r47 3 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.83 $Y=0.555
+ $X2=1.83 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_193_47# 1 2 9 11 12 15 18 21 23 25 28 29
+ 30 32 33 34 41 42 45 46 53 58
c195 46 0 4.49643e-20 $X=5.31 $Y=1.19
c196 45 0 2.56901e-19 $X=5.31 $Y=1.19
c197 41 0 3.30612e-20 $X=2.99 $Y=0.85
c198 34 0 2.53448e-20 $X=3.135 $Y=1.19
c199 33 0 1.51904e-19 $X=5.165 $Y=1.19
c200 32 0 9.52104e-20 $X=3.027 $Y=1.12
c201 25 0 1.80017e-19 $X=5.605 $Y=2.275
c202 23 0 1.753e-19 $X=5.605 $Y=1.455
c203 9 0 4.43992e-20 $X=2.315 $Y=2.275
r204 53 56 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=1.095
r205 53 55 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=0.93
+ $X2=2.915 $Y2=0.765
r206 46 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.26 $X2=5.315 $Y2=1.26
r207 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.31 $Y=1.19
+ $X2=5.31 $Y2=1.19
r208 42 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=0.93 $X2=2.915 $Y2=0.93
r209 41 43 0.0661242 $w=2.9e-07 $l=1.15e-07 $layer=MET1_cond $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.965
r210 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0.85
+ $X2=2.99 $Y2=0.85
r211 37 62 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=1.96
r212 37 58 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.127 $Y=0.85
+ $X2=1.127 $Y2=0.51
r213 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0.85
+ $X2=1.15 $Y2=0.85
r214 33 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.165 $Y=1.19
+ $X2=5.31 $Y2=1.19
r215 33 34 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=5.165 $Y=1.19
+ $X2=3.135 $Y2=1.19
r216 32 34 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.135 $Y2=1.19
r217 32 43 0.110669 $w=2.15e-07 $l=1.55e-07 $layer=MET1_cond $X=3.027 $Y=1.12
+ $X2=3.027 $Y2=0.965
r218 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=0.85
+ $X2=1.15 $Y2=0.85
r219 29 41 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=2.99 $Y2=0.85
r220 29 30 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=2.845 $Y=0.85
+ $X2=1.295 $Y2=0.85
r221 28 49 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.47 $Y=1.26
+ $X2=5.315 $Y2=1.26
r222 23 28 52.102 $w=1.88e-07 $l=2.09464e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.575 $Y2=1.26
r223 23 25 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.605 $Y=1.455
+ $X2=5.605 $Y2=2.275
r224 19 28 36.719 $w=1.88e-07 $l=1.39911e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.575 $Y2=1.26
r225 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.565 $Y=1.125
+ $X2=5.565 $Y2=0.445
r226 18 56 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=1.245
+ $X2=2.855 $Y2=1.095
r227 15 55 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.855 $Y=0.415
+ $X2=2.855 $Y2=0.765
r228 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.855 $Y2=1.245
r229 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.78 $Y=1.32
+ $X2=2.39 $Y2=1.32
r230 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.39 $Y2=1.32
r231 7 9 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.315 $Y=1.395
+ $X2=2.315 $Y2=2.275
r232 2 62 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r233 1 58 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_652_21# 1 2 9 13 15 19 21 25 28 30 31 35
+ 38
c115 38 0 1.30404e-19 $X=4.625 $Y=0.895
c116 35 0 2.11834e-19 $X=4.075 $Y=1.96
c117 28 0 3.15264e-19 $X=4.625 $Y=1.835
c118 21 0 1.75093e-19 $X=4.54 $Y=1.96
r119 36 38 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.435 $Y=0.895
+ $X2=4.625 $Y2=0.895
r120 31 42 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.905
r121 31 41 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.74
+ $X2=3.42 $Y2=1.575
r122 30 33 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=3.485 $Y=1.74
+ $X2=3.485 $Y2=1.96
r123 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.74 $X2=3.445 $Y2=1.74
r124 27 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=0.895
r125 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.625 $Y=1.065
+ $X2=4.625 $Y2=1.835
r126 23 36 2.53954 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.895
r127 23 25 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.435 $Y=0.725
+ $X2=4.435 $Y2=0.46
r128 22 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.96
+ $X2=4.075 $Y2=1.96
r129 21 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.625 $Y2=1.835
r130 21 22 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.54 $Y=1.96
+ $X2=4.16 $Y2=1.96
r131 17 35 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=1.96
r132 17 19 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=2.085
+ $X2=4.075 $Y2=2.21
r133 16 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=1.96
+ $X2=3.485 $Y2=1.96
r134 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=4.075 $Y2=1.96
r135 15 16 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=3.99 $Y=1.96
+ $X2=3.61 $Y2=1.96
r136 13 42 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.335 $Y=2.275
+ $X2=3.335 $Y2=1.905
r137 9 41 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.335 $Y=0.445
+ $X2=3.335 $Y2=1.575
r138 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=2.065 $X2=4.075 $Y2=2.21
r139 1 25 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.235 $X2=4.475 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%SET_B 1 3 7 11 17 19 20 24 26 27 29 30 36 37
c134 37 0 1.72331e-19 $X=7.13 $Y=0.85
c135 29 0 2.95874e-19 $X=6.985 $Y=0.85
c136 26 0 1.49785e-19 $X=6.99 $Y=0.9
c137 19 0 1.13317e-19 $X=6.895 $Y=1.535
c138 1 0 9.39349e-20 $X=3.865 $Y=1.145
r139 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0.85
+ $X2=7.13 $Y2=0.85
r140 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.055 $Y=0.85
+ $X2=3.91 $Y2=0.85
r141 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=7.13 $Y2=0.85
r142 29 30 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=6.985 $Y=0.85
+ $X2=4.055 $Y2=0.85
r143 27 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=0.98 $X2=3.775 $Y2=0.98
r144 27 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0.85
+ $X2=3.91 $Y2=0.85
r145 26 37 5.97563 $w=2.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.99 $Y=0.87
+ $X2=7.13 $Y2=0.87
r146 24 44 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=1.145
r147 24 43 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=0.98
+ $X2=6.825 $Y2=0.815
r148 23 26 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0.9
+ $X2=6.99 $Y2=0.9
r149 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.825
+ $Y=0.98 $X2=6.825 $Y2=0.98
r150 19 20 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=6.895 $Y=1.535
+ $X2=6.895 $Y2=1.685
r151 19 44 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.885 $Y=1.535
+ $X2=6.885 $Y2=1.145
r152 17 20 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.905 $Y=2.275
+ $X2=6.905 $Y2=1.685
r153 11 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.765 $Y=0.445
+ $X2=6.765 $Y2=0.815
r154 5 40 38.5432 $w=3.18e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.81 $Y2=0.98
r155 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.905 $Y=0.815
+ $X2=3.905 $Y2=0.445
r156 1 40 38.5432 $w=3.18e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.81 $Y2=0.98
r157 1 3 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.865 $Y=1.145
+ $X2=3.865 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_476_47# 1 2 7 9 11 14 16 20 22 24 25 26 30
+ 35 37 38 43 44 53
c157 53 0 1.95729e-19 $X=4.705 $Y=1.4
c158 43 0 4.43992e-20 $X=3.44 $Y=1.3
c159 26 0 1.01003e-19 $X=3.02 $Y=2.335
c160 22 0 3.64688e-20 $X=5.205 $Y=0.735
c161 16 0 1.15925e-19 $X=5.13 $Y=0.825
c162 7 0 3.12358e-20 $X=4.265 $Y=0.735
r163 48 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.705 $Y2=1.4
r164 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.285 $Y=1.4
+ $X2=4.265 $Y2=1.4
r165 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.4 $X2=4.285 $Y2=1.4
r166 44 47 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.245 $Y=1.32
+ $X2=4.245 $Y2=1.4
r167 42 43 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=1.3
+ $X2=3.44 $Y2=1.3
r168 40 42 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=3.105 $Y=1.3
+ $X2=3.355 $Y2=1.3
r169 38 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=4.245 $Y2=1.32
r170 38 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.12 $Y=1.32
+ $X2=3.44 $Y2=1.32
r171 37 42 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.355 $Y=1.195
+ $X2=3.355 $Y2=1.3
r172 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.355 $Y=0.465
+ $X2=3.355 $Y2=1.195
r173 34 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=1.3
r174 34 35 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.105 $Y=1.405
+ $X2=3.105 $Y2=2.25
r175 30 36 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=3.355 $Y2=0.465
r176 30 32 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.27 $Y=0.365
+ $X2=2.59 $Y2=0.365
r177 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.105 $Y2=2.25
r178 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=2.525 $Y2=2.335
r179 22 24 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.205 $Y=0.735
+ $X2=5.205 $Y2=0.445
r180 18 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=1.4
r181 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.705 $Y=1.565
+ $X2=4.705 $Y2=2.275
r182 17 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.34 $Y=0.825
+ $X2=4.265 $Y2=0.825
r183 16 22 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=5.205 $Y2=0.735
r184 16 17 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=5.13 $Y=0.825
+ $X2=4.34 $Y2=0.825
r185 12 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=1.4
r186 12 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.285 $Y=1.565
+ $X2=4.285 $Y2=2.275
r187 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.235
+ $X2=4.265 $Y2=1.4
r188 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=0.825
r189 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.265 $Y=0.915
+ $X2=4.265 $Y2=1.235
r190 7 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.825
r191 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.265 $Y=0.735
+ $X2=4.265 $Y2=0.445
r192 2 28 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.065 $X2=2.525 $Y2=2.335
r193 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_1178_261# 1 2 9 13 18 21 25 29 32 36 39 40
c80 39 0 1.80017e-19 $X=7.51 $Y=1.67
c81 32 0 1.13317e-19 $X=7.745 $Y=1.575
c82 18 0 6.36338e-20 $X=6.405 $Y=1.38
r83 38 40 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.745 $Y2=1.67
r84 38 39 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=1.67
+ $X2=7.51 $Y2=1.67
r85 34 36 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=7.595 $Y=0.515
+ $X2=7.745 $Y2=0.515
r86 32 40 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=7.745 $Y=1.575
+ $X2=7.745 $Y2=1.67
r87 31 36 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0.68
+ $X2=7.745 $Y2=0.515
r88 31 32 47.2684 $w=2.08e-07 $l=8.95e-07 $layer=LI1_cond $X=7.745 $Y=0.68
+ $X2=7.745 $Y2=1.575
r89 27 38 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.67
r90 27 29 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.595 $Y=1.765
+ $X2=7.595 $Y2=1.87
r91 24 39 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=6.075 $Y=1.66
+ $X2=7.51 $Y2=1.66
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.075
+ $Y=1.66 $X2=6.075 $Y2=1.66
r93 20 25 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=6.05 $Y=1.665
+ $X2=6.05 $Y2=1.66
r94 20 21 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=6.05 $Y=1.665
+ $X2=6.05 $Y2=1.825
r95 16 25 36.9668 $w=3.2e-07 $l=2.05e-07 $layer=POLY_cond $X=6.05 $Y=1.455
+ $X2=6.05 $Y2=1.66
r96 16 18 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.05 $Y=1.38
+ $X2=6.405 $Y2=1.38
r97 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=1.38
r98 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.405 $Y2=0.445
r99 9 21 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=5.965 $Y=2.275
+ $X2=5.965 $Y2=1.825
r100 2 29 300 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=2 $X=7.46
+ $Y=1.645 $X2=7.595 $Y2=1.87
r101 1 34 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_1028_413# 1 2 3 12 16 18 22 26 28 29 34 35
+ 39 40 41 44 49 51 54 56 57 58
c162 54 0 9.39049e-20 $X=6.405 $Y=1.32
c163 34 0 7.39505e-20 $X=5.655 $Y=1.915
c164 29 0 1.39518e-19 $X=5.57 $Y=2.29
r165 56 58 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=1.29
+ $X2=7.14 $Y2=1.29
r166 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.305
+ $Y=1.26 $X2=7.305 $Y2=1.26
r167 47 49 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=2.085
+ $X2=6.66 $Y2=2.21
r168 46 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=6.405 $Y2=1.32
r169 46 58 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.49 $Y=1.32
+ $X2=7.14 $Y2=1.32
r170 44 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.235
+ $X2=6.405 $Y2=1.32
r171 43 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.405 $Y=0.475
+ $X2=6.405 $Y2=1.235
r172 42 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.74 $Y=2 $X2=5.655
+ $Y2=2
r173 41 47 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=6.54 $Y=2
+ $X2=6.66 $Y2=2.085
r174 41 42 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=6.54 $Y=2 $X2=5.74
+ $Y2=2
r175 39 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=6.405 $Y2=1.32
r176 39 40 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=6.32 $Y=1.32
+ $X2=5.74 $Y2=1.32
r177 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=6.405 $Y2=0.475
r178 35 37 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.32 $Y=0.39
+ $X2=5.805 $Y2=0.39
r179 34 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=1.915
+ $X2=5.655 $Y2=2
r180 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.655 $Y=1.405
+ $X2=5.74 $Y2=1.32
r181 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.655 $Y=1.405
+ $X2=5.655 $Y2=1.915
r182 29 51 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.655 $Y=2.29
+ $X2=5.655 $Y2=2
r183 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.57 $Y=2.29
+ $X2=5.275 $Y2=2.29
r184 24 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=1.425
+ $X2=8.325 $Y2=1.26
r185 24 26 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.325 $Y=1.425
+ $X2=8.325 $Y2=2.165
r186 20 28 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=1.095
+ $X2=8.325 $Y2=1.26
r187 20 22 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=8.325 $Y=1.095
+ $X2=8.325 $Y2=0.445
r188 19 57 5.03009 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.46 $Y=1.26
+ $X2=7.315 $Y2=1.26
r189 18 28 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.25 $Y=1.26
+ $X2=8.325 $Y2=1.26
r190 18 19 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=8.25 $Y=1.26
+ $X2=7.46 $Y2=1.26
r191 14 57 37.0704 $w=1.5e-07 $l=1.96914e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.315 $Y2=1.26
r192 14 16 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.385 $Y=1.425
+ $X2=7.385 $Y2=2.065
r193 10 57 37.0704 $w=1.5e-07 $l=1.96914e-07 $layer=POLY_cond $X=7.385 $Y=1.095
+ $X2=7.315 $Y2=1.26
r194 10 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.385 $Y=1.095
+ $X2=7.385 $Y2=0.505
r195 3 49 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.065 $X2=6.695 $Y2=2.21
r196 2 31 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=2.065 $X2=5.275 $Y2=2.33
r197 1 37 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=5.64
+ $Y=0.235 $X2=5.805 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_1598_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 51 60 64 65 66 74
r126 71 72 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.64 $Y=1.16
+ $X2=10.06 $Y2=1.16
r127 70 71 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=9.22 $Y=1.16
+ $X2=9.64 $Y2=1.16
r128 64 65 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=2
+ $X2=8.115 $Y2=1.915
r129 61 74 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=10.25 $Y=1.16
+ $X2=10.48 $Y2=1.16
r130 61 72 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=10.25 $Y=1.16
+ $X2=10.06 $Y2=1.16
r131 60 61 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.25
+ $Y=1.16 $X2=10.25 $Y2=1.16
r132 58 70 73.3173 $w=2.7e-07 $l=3.3e-07 $layer=POLY_cond $X=8.89 $Y=1.16
+ $X2=9.22 $Y2=1.16
r133 58 67 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=8.89 $Y=1.16 $X2=8.8
+ $Y2=1.16
r134 57 60 71.2419 $w=2.18e-07 $l=1.36e-06 $layer=LI1_cond $X=8.89 $Y=1.165
+ $X2=10.25 $Y2=1.165
r135 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.89
+ $Y=1.16 $X2=8.89 $Y2=1.16
r136 55 66 1.80668 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.28 $Y=1.165
+ $X2=8.155 $Y2=1.165
r137 55 57 31.9541 $w=2.18e-07 $l=6.1e-07 $layer=LI1_cond $X=8.28 $Y=1.165
+ $X2=8.89 $Y2=1.165
r138 53 66 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.155 $Y=1.275
+ $X2=8.155 $Y2=1.165
r139 53 65 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=8.155 $Y=1.275
+ $X2=8.155 $Y2=1.915
r140 49 66 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.155 $Y=1.055
+ $X2=8.155 $Y2=1.165
r141 49 51 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=8.155 $Y=1.055
+ $X2=8.155 $Y2=0.51
r142 43 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.48 $Y=1.295
+ $X2=10.48 $Y2=1.16
r143 43 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.48 $Y=1.295
+ $X2=10.48 $Y2=1.985
r144 39 74 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.48 $Y=1.025
+ $X2=10.48 $Y2=1.16
r145 39 41 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.48 $Y=1.025
+ $X2=10.48 $Y2=0.56
r146 35 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=1.295
+ $X2=10.06 $Y2=1.16
r147 35 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=10.06 $Y=1.295
+ $X2=10.06 $Y2=1.985
r148 31 72 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=1.025
+ $X2=10.06 $Y2=1.16
r149 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.06 $Y=1.025
+ $X2=10.06 $Y2=0.56
r150 27 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.64 $Y=1.295
+ $X2=9.64 $Y2=1.16
r151 27 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.64 $Y=1.295
+ $X2=9.64 $Y2=1.985
r152 23 71 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.64 $Y=1.025
+ $X2=9.64 $Y2=1.16
r153 23 25 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.64 $Y=1.025
+ $X2=9.64 $Y2=0.56
r154 19 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.22 $Y=1.295
+ $X2=9.22 $Y2=1.16
r155 19 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.22 $Y=1.295
+ $X2=9.22 $Y2=1.985
r156 15 70 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.22 $Y=1.025
+ $X2=9.22 $Y2=1.16
r157 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.22 $Y=1.025
+ $X2=9.22 $Y2=0.56
r158 11 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.8 $Y=1.295
+ $X2=8.8 $Y2=1.16
r159 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.8 $Y=1.295
+ $X2=8.8 $Y2=1.985
r160 7 67 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=8.8 $Y=1.025
+ $X2=8.8 $Y2=1.16
r161 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.8 $Y=1.025 $X2=8.8
+ $Y2=0.56
r162 2 64 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=7.99
+ $Y=1.845 $X2=8.115 $Y2=2
r163 1 51 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=7.99
+ $Y=0.235 $X2=8.115 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 36 40 44 48 52
+ 56 58 60 62 68 73 78 86 91 96 101 108 109 112 115 118 125 128 135 138 141 144
c195 109 0 1.81794e-19 $X=10.81 $Y=2.72
c196 1 0 3.29888e-20 $X=0.545 $Y=1.815
r197 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r198 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r199 138 139 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r200 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r201 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r202 128 131 10.4269 $w=4.18e-07 $l=3.8e-07 $layer=LI1_cond $X=6.13 $Y=2.34
+ $X2=6.13 $Y2=2.72
r203 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r204 122 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r205 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r206 118 121 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.62 $Y=2.34
+ $X2=3.62 $Y2=2.72
r207 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r208 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r209 109 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r210 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r211 106 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.435 $Y=2.72
+ $X2=10.27 $Y2=2.72
r212 106 108 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.435 $Y=2.72
+ $X2=10.81 $Y2=2.72
r213 105 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r214 105 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r215 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r216 102 141 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.595 $Y=2.72
+ $X2=9.467 $Y2=2.72
r217 102 104 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.595 $Y=2.72
+ $X2=9.89 $Y2=2.72
r218 101 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.105 $Y=2.72
+ $X2=10.27 $Y2=2.72
r219 101 104 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.105 $Y=2.72
+ $X2=9.89 $Y2=2.72
r220 100 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r221 100 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r222 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r223 97 138 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.745 $Y=2.72
+ $X2=8.602 $Y2=2.72
r224 97 99 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.745 $Y=2.72
+ $X2=8.97 $Y2=2.72
r225 96 141 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.34 $Y=2.72
+ $X2=9.467 $Y2=2.72
r226 96 99 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.34 $Y=2.72
+ $X2=8.97 $Y2=2.72
r227 95 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r228 95 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r229 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r230 92 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.175 $Y2=2.72
r231 92 94 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.34 $Y=2.72
+ $X2=7.59 $Y2=2.72
r232 91 138 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.46 $Y=2.72
+ $X2=8.602 $Y2=2.72
r233 91 94 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.46 $Y=2.72
+ $X2=7.59 $Y2=2.72
r234 90 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r235 90 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=6.21 $Y2=2.72
r236 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r237 87 131 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.13 $Y2=2.72
r238 87 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.34 $Y=2.72
+ $X2=6.67 $Y2=2.72
r239 86 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.175 $Y2=2.72
r240 86 89 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r241 85 132 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r242 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r243 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r244 82 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r245 81 84 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r246 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r247 79 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.495 $Y2=2.72
r248 79 81 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.66 $Y=2.72
+ $X2=4.83 $Y2=2.72
r249 78 131 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.13 $Y2=2.72
r250 78 84 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.75 $Y2=2.72
r251 77 122 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r252 77 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r253 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r254 74 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.62 $Y2=2.72
r255 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=2.07 $Y2=2.72
r256 73 121 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=3.62 $Y2=2.72
r257 73 76 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.43 $Y=2.72
+ $X2=2.07 $Y2=2.72
r258 72 116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r259 72 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r260 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r261 69 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r262 69 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r263 68 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.62 $Y2=2.72
r264 68 71 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r265 62 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r266 60 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r267 58 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r268 58 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r269 54 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.27 $Y=2.635
+ $X2=10.27 $Y2=2.72
r270 54 56 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=10.27 $Y=2.635
+ $X2=10.27 $Y2=2.02
r271 50 141 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.467 $Y=2.635
+ $X2=9.467 $Y2=2.72
r272 50 52 21.4671 $w=2.53e-07 $l=4.75e-07 $layer=LI1_cond $X=9.467 $Y=2.635
+ $X2=9.467 $Y2=2.16
r273 46 138 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.602 $Y=2.635
+ $X2=8.602 $Y2=2.72
r274 46 48 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=8.602 $Y=2.635
+ $X2=8.602 $Y2=2
r275 42 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.72
r276 42 44 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.175 $Y=2.635
+ $X2=7.175 $Y2=2.21
r277 38 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.72
r278 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.495 $Y=2.635
+ $X2=4.495 $Y2=2.34
r279 37 121 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.62 $Y2=2.72
r280 36 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=4.495 $Y2=2.72
r281 36 37 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.81 $Y2=2.72
r282 32 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.72
r283 32 34 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.62 $Y=2.635
+ $X2=1.62 $Y2=2.22
r284 28 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r285 28 30 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r286 9 56 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=10.135
+ $Y=1.485 $X2=10.27 $Y2=2.02
r287 8 52 600 $w=1.7e-07 $l=7.39425e-07 $layer=licon1_PDIFF $count=1 $X=9.295
+ $Y=1.485 $X2=9.43 $Y2=2.16
r288 7 48 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=8.4
+ $Y=1.845 $X2=8.59 $Y2=2
r289 6 44 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=6.98
+ $Y=2.065 $X2=7.175 $Y2=2.21
r290 5 128 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.04
+ $Y=2.065 $X2=6.175 $Y2=2.34
r291 4 40 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.065 $X2=4.495 $Y2=2.34
r292 3 118 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.065 $X2=3.595 $Y2=2.34
r293 2 34 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.645 $X2=1.62 $Y2=2.22
r294 1 30 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%A_381_47# 1 2 8 9 10 11 12 15 20
c59 20 0 1.34441e-19 $X=2.04 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0.635
+ $X2=2.04 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=2.04 $Y2=1.88
r62 11 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=1.88
+ $X2=1.6 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=2.04 $Y2=0.635
r64 9 10 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=1.955 $Y=0.73
+ $X2=1.6 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.515 $Y=1.795
+ $X2=1.6 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.6 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.515 $Y=0.825
+ $X2=1.515 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.645 $X2=2.04 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%Q 1 2 3 4 5 6 19 20 21 22 23 28 30 32 36 37
+ 38 39 40 41 42 43 44 45 46 83
r78 81 83 5.92685 $w=3.48e-07 $l=1.8e-07 $layer=LI1_cond $X=10.78 $Y=1.64
+ $X2=10.78 $Y2=1.82
r79 69 74 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=0.715
+ $X2=10.78 $Y2=0.63
r80 45 46 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=10.78 $Y=1.87
+ $X2=10.78 $Y2=2.21
r81 45 83 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=10.78 $Y=1.87
+ $X2=10.78 $Y2=1.82
r82 44 76 3.24686 $w=2.9e-07 $l=1.11018e-07 $layer=LI1_cond $X=10.78 $Y=1.555
+ $X2=10.84 $Y2=1.47
r83 44 81 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=1.555
+ $X2=10.78 $Y2=1.64
r84 44 76 0.651381 $w=2.28e-07 $l=1.3e-08 $layer=LI1_cond $X=10.84 $Y=1.457
+ $X2=10.84 $Y2=1.47
r85 43 44 13.3784 $w=2.28e-07 $l=2.67e-07 $layer=LI1_cond $X=10.84 $Y=1.19
+ $X2=10.84 $Y2=1.457
r86 42 69 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.78 $Y=0.8
+ $X2=10.78 $Y2=0.715
r87 42 75 3.24686 $w=2.9e-07 $l=1.11018e-07 $layer=LI1_cond $X=10.78 $Y=0.8
+ $X2=10.84 $Y2=0.885
r88 42 43 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=10.84 $Y=0.91
+ $X2=10.84 $Y2=1.19
r89 42 75 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=10.84 $Y=0.91
+ $X2=10.84 $Y2=0.885
r90 41 74 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=10.78 $Y=0.51
+ $X2=10.78 $Y2=0.63
r91 39 40 18.345 $w=2.43e-07 $l=3.9e-07 $layer=LI1_cond $X=9.047 $Y=1.82
+ $X2=9.047 $Y2=2.21
r92 38 62 5.64462 $w=2.43e-07 $l=1.2e-07 $layer=LI1_cond $X=9.047 $Y=0.51
+ $X2=9.047 $Y2=0.63
r93 35 39 8.46693 $w=2.43e-07 $l=1.8e-07 $layer=LI1_cond $X=9.047 $Y=1.64
+ $X2=9.047 $Y2=1.82
r94 34 62 3.99827 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=9.047 $Y=0.715
+ $X2=9.047 $Y2=0.63
r95 33 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=1.555
+ $X2=9.85 $Y2=1.555
r96 32 44 3.3199 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=10.605 $Y=1.555
+ $X2=10.78 $Y2=1.555
r97 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.605 $Y=1.555
+ $X2=9.935 $Y2=1.555
r98 31 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.935 $Y=0.8 $X2=9.85
+ $Y2=0.8
r99 30 42 3.3199 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=10.605 $Y=0.8
+ $X2=10.78 $Y2=0.8
r100 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.605 $Y=0.8
+ $X2=9.935 $Y2=0.8
r101 26 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.85 $Y=1.64
+ $X2=9.85 $Y2=1.555
r102 26 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.85 $Y=1.64
+ $X2=9.85 $Y2=1.82
r103 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.85 $Y=0.715
+ $X2=9.85 $Y2=0.8
r104 23 25 6.1 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.85 $Y=0.715 $X2=9.85
+ $Y2=0.63
r105 22 35 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=9.17 $Y=1.555
+ $X2=9.047 $Y2=1.64
r106 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.765 $Y=1.555
+ $X2=9.85 $Y2=1.555
r107 21 22 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=9.765 $Y=1.555
+ $X2=9.17 $Y2=1.555
r108 20 34 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=9.17 $Y=0.8
+ $X2=9.047 $Y2=0.715
r109 19 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.765 $Y=0.8
+ $X2=9.85 $Y2=0.8
r110 19 20 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=9.765 $Y=0.8
+ $X2=9.17 $Y2=0.8
r111 6 83 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=10.555
+ $Y=1.485 $X2=10.69 $Y2=1.82
r112 5 28 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=9.715
+ $Y=1.485 $X2=9.85 $Y2=1.82
r113 4 39 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=8.875
+ $Y=1.485 $X2=9.01 $Y2=1.82
r114 3 74 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=10.555
+ $Y=0.235 $X2=10.69 $Y2=0.63
r115 2 25 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=0.235 $X2=9.85 $Y2=0.63
r116 1 62 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=0.235 $X2=9.01 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HD__DFSTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53
+ 55 57 63 68 76 86 91 96 103 104 107 110 113 116 121 127 129 132 135
c183 121 0 1.49785e-19 $X=6.67 $Y=0.24
c184 104 0 1.99443e-19 $X=10.81 $Y=0
r185 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r186 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r187 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r188 125 127 11.126 $w=6.48e-07 $l=2e-07 $layer=LI1_cond $X=7.13 $Y=0.24
+ $X2=7.33 $Y2=0.24
r189 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r190 123 125 1.01207 $w=6.48e-07 $l=5.5e-08 $layer=LI1_cond $X=7.075 $Y=0.24
+ $X2=7.13 $Y2=0.24
r191 120 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r192 119 123 7.45249 $w=6.48e-07 $l=4.05e-07 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=7.075 $Y2=0.24
r193 119 121 7.44573 $w=6.48e-07 $l=4.45988e-08 $layer=LI1_cond $X=6.67 $Y=0.24
+ $X2=6.67 $Y2=0.24
r194 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r195 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r196 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r197 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r198 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r199 104 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=10.35 $Y2=0
r200 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r201 101 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.435 $Y=0
+ $X2=10.27 $Y2=0
r202 101 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.435 $Y=0
+ $X2=10.81 $Y2=0
r203 100 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r204 100 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=9.43 $Y2=0
r205 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r206 97 132 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.595 $Y=0
+ $X2=9.467 $Y2=0
r207 97 99 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.595 $Y=0 $X2=9.89
+ $Y2=0
r208 96 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.105 $Y=0
+ $X2=10.27 $Y2=0
r209 96 99 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.105 $Y=0
+ $X2=9.89 $Y2=0
r210 95 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r211 95 130 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.51 $Y2=0
r212 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r213 92 129 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.745 $Y=0
+ $X2=8.602 $Y2=0
r214 92 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.745 $Y=0
+ $X2=8.97 $Y2=0
r215 91 132 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.34 $Y=0
+ $X2=9.467 $Y2=0
r216 91 94 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.34 $Y=0 $X2=8.97
+ $Y2=0
r217 90 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r218 90 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r219 89 127 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.59 $Y=0 $X2=7.33
+ $Y2=0
r220 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r221 86 129 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.46 $Y=0
+ $X2=8.602 $Y2=0
r222 86 89 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.46 $Y=0 $X2=7.59
+ $Y2=0
r223 85 120 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r224 85 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=4.83 $Y2=0
r225 84 121 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=6.67 $Y2=0
r226 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r227 82 116 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.91
+ $Y2=0
r228 82 84 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.29
+ $Y2=0
r229 80 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r230 80 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=3.91 $Y2=0
r231 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r232 77 113 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0
+ $X2=3.815 $Y2=0
r233 77 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.37
+ $Y2=0
r234 76 116 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.91
+ $Y2=0
r235 76 79 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.37
+ $Y2=0
r236 75 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=3.91 $Y2=0
r237 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r238 72 75 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r239 72 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r240 71 74 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r241 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r242 69 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.62 $Y2=0
r243 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.07 $Y2=0
r244 68 113 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.61 $Y=0
+ $X2=3.815 $Y2=0
r245 68 74 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.45
+ $Y2=0
r246 67 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r247 67 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r248 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r249 64 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.68 $Y2=0
r250 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.15 $Y2=0
r251 63 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.62 $Y2=0
r252 63 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r253 57 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.68 $Y2=0
r254 55 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r255 53 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r256 53 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r257 49 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.27 $Y=0.085
+ $X2=10.27 $Y2=0
r258 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.27 $Y=0.085
+ $X2=10.27 $Y2=0.38
r259 45 132 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.467 $Y=0.085
+ $X2=9.467 $Y2=0
r260 45 47 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=9.467 $Y=0.085
+ $X2=9.467 $Y2=0.38
r261 41 129 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.602 $Y=0.085
+ $X2=8.602 $Y2=0
r262 41 43 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=8.602 $Y=0.085
+ $X2=8.602 $Y2=0.38
r263 37 116 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0
r264 37 39 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=4.91 $Y=0.085
+ $X2=4.91 $Y2=0.38
r265 33 113 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r266 33 35 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.36
r267 29 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r268 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.38
r269 25 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r270 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r271 8 51 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=0.235 $X2=10.27 $Y2=0.38
r272 7 47 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.235 $X2=9.43 $Y2=0.38
r273 6 43 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=8.4
+ $Y=0.235 $X2=8.59 $Y2=0.38
r274 5 123 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.235 $X2=7.075 $Y2=0.48
r275 4 39 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=4.995 $Y2=0.38
r276 3 35 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.235 $X2=3.695 $Y2=0.36
r277 2 31 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.38
r278 1 27 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o21ba_2.pex.spice
* Created: Tue Sep  1 19:21:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21BA_2%B1_N 3 6 8 9 13 15
c36 13 0 1.51906e-19 $X=0.51 $Y=1.16
r37 17 22 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=1.325
+ $X2=0.685 $Y2=1.16
r38 14 22 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.51 $Y=1.16
+ $X2=0.685 $Y2=1.16
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.16
+ $X2=0.51 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r42 9 17 12.6313 $w=1.78e-07 $l=2.05e-07 $layer=LI1_cond $X=0.685 $Y=1.53
+ $X2=0.685 $Y2=1.325
r43 8 22 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.685
+ $Y2=1.16
r44 6 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.695
+ $X2=0.47 $Y2=1.325
r45 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.675
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%A_174_21# 1 2 7 9 12 14 16 19 21 25 28 31 35
+ 38 40 48
c101 48 0 1.5767e-19 $X=1.375 $Y=1.16
c102 35 0 6.65026e-20 $X=2.107 $Y=0.74
c103 31 0 7.75504e-20 $X=1.44 $Y=0.74
r104 45 46 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.955 $Y=1.16
+ $X2=1.365 $Y2=1.16
r105 43 45 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.945 $Y=1.16
+ $X2=0.955 $Y2=1.16
r106 38 40 0.474307 $w=5.78e-07 $l=2.3e-08 $layer=LI1_cond $X=2.562 $Y=1.745
+ $X2=2.585 $Y2=1.745
r107 36 38 7.6714 $w=5.78e-07 $l=3.72e-07 $layer=LI1_cond $X=2.19 $Y=1.745
+ $X2=2.562 $Y2=1.745
r108 34 48 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.375 $Y2=1.16
r109 34 46 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.37 $Y=1.16
+ $X2=1.365 $Y2=1.16
r110 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r111 31 33 24.9951 $w=2.05e-07 $l=4.2e-07 $layer=LI1_cond $X=1.44 $Y=0.74
+ $X2=1.44 $Y2=1.16
r112 28 36 8.09873 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=2.19 $Y=1.455
+ $X2=2.19 $Y2=1.745
r113 27 35 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=2.19 $Y=0.825
+ $X2=2.107 $Y2=0.74
r114 27 28 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.19 $Y=0.825
+ $X2=2.19 $Y2=1.455
r115 23 35 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=0.655
+ $X2=2.107 $Y2=0.74
r116 23 25 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=2.107 $Y=0.655
+ $X2=2.107 $Y2=0.38
r117 22 31 1.83547 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.595 $Y=0.74
+ $X2=1.44 $Y2=0.74
r118 21 35 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.94 $Y=0.74
+ $X2=2.107 $Y2=0.74
r119 21 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.94 $Y=0.74
+ $X2=1.595 $Y2=0.74
r120 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.16
r121 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.375 $Y=1.325
+ $X2=1.375 $Y2=1.985
r122 14 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r123 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.56
r124 10 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.16
r125 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=1.325
+ $X2=0.955 $Y2=1.985
r126 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=1.16
r127 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.945 $Y=0.995
+ $X2=0.945 $Y2=0.56
r128 2 40 300 $w=1.7e-07 $l=5.64137e-07 $layer=licon1_PDIFF $count=2 $X=2.39
+ $Y=1.485 $X2=2.585 $Y2=1.96
r129 2 40 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.485 $X2=2.585 $Y2=1.62
r130 1 25 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.235 $X2=2.105 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%A_27_93# 1 2 7 9 12 14 15 18 21 22 23 26 32
+ 34
c76 22 0 1.51906e-19 $X=1.765 $Y=1.95
r77 29 32 2.62582 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.627 $X2=0.26
+ $Y2=0.627
r78 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.16 $X2=1.85 $Y2=1.16
r79 24 26 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.85 $Y=1.865
+ $X2=1.85 $Y2=1.16
r80 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.765 $Y=1.95
+ $X2=1.85 $Y2=1.865
r81 22 23 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.765 $Y=1.95
+ $X2=0.395 $Y2=1.95
r82 19 23 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.24 $Y=1.865
+ $X2=0.395 $Y2=1.95
r83 19 21 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=1.865
+ $X2=0.24 $Y2=1.66
r84 18 34 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=1.65
+ $X2=0.24 $Y2=1.495
r85 18 21 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=1.65 $X2=0.24
+ $Y2=1.66
r86 16 29 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.627
r87 16 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.495
r88 14 27 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=2.24 $Y=1.16
+ $X2=1.85 $Y2=1.16
r89 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.24 $Y=1.16
+ $X2=2.315 $Y2=1.16
r90 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.16
r91 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.315 $Y=1.325
+ $X2=2.315 $Y2=1.985
r92 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=1.16
r93 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=0.56
r94 2 21 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r95 1 32 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%A2 3 6 8 11 12 13
c37 13 0 6.65026e-20 $X=2.735 $Y=0.995
c38 11 0 1.44727e-19 $X=2.735 $Y=1.16
r39 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.735 $Y2=1.325
r40 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.16
+ $X2=2.735 $Y2=0.995
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r42 8 12 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=2.53 $Y=1.18
+ $X2=2.735 $Y2=1.18
r43 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.795 $Y=1.985
+ $X2=2.795 $Y2=1.325
r44 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.79 $Y=0.56 $X2=2.79
+ $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%A1 3 7 8 9 13 14 15
r29 13 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=3.255 $Y2=1.325
r30 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=3.255 $Y2=0.995
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.16 $X2=3.265 $Y2=1.16
r32 8 9 8.21549 $w=4.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.347 $Y=1.19
+ $X2=3.347 $Y2=1.53
r33 8 14 0.724896 $w=4.93e-07 $l=3e-08 $layer=LI1_cond $X=3.347 $Y=1.19
+ $X2=3.347 $Y2=1.16
r34 7 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.21 $Y=0.56 $X2=3.21
+ $Y2=0.995
r35 3 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.155 $Y=1.985
+ $X2=3.155 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%VPWR 1 2 3 12 14 16 18 20 30 36 40 44 47
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 42 44 10.0564 $w=5.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.07 $Y=2.505
+ $X2=2.23 $Y2=2.505
r57 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 39 42 0.0996732 $w=5.98e-07 $l=5e-09 $layer=LI1_cond $X=2.065 $Y=2.505
+ $X2=2.07 $Y2=2.505
r59 39 40 19.8244 $w=5.98e-07 $l=6.5e-07 $layer=LI1_cond $X=2.065 $Y=2.505
+ $X2=1.415 $Y2=2.505
r60 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r61 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 34 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 33 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.23 $Y2=2.72
r64 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 30 46 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.2 $Y=2.72 $X2=3.44
+ $Y2=2.72
r66 30 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.2 $Y=2.72 $X2=2.99
+ $Y2=2.72
r67 29 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r68 29 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 28 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.415 $Y2=2.72
r70 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 26 36 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=0.715 $Y2=2.72
r72 26 28 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.91 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 20 36 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.715 $Y2=2.72
r74 20 22 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r75 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r77 14 46 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.365 $Y=2.635
+ $X2=3.44 $Y2=2.72
r78 14 16 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.365 $Y=2.635
+ $X2=3.365 $Y2=1.96
r79 10 36 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r80 10 12 10.1947 $w=3.88e-07 $l=3.45e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.29
r81 3 16 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=3.23
+ $Y=1.485 $X2=3.365 $Y2=1.96
r82 2 39 300 $w=1.7e-07 $l=1.06916e-06 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=1.485 $X2=2.065 $Y2=2.29
r83 1 12 600 $w=1.7e-07 $l=8.99458e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.745 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%X 1 2 8 11 13 23
r29 13 23 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=0.425
+ $X2=1.155 $Y2=0.425
r30 13 18 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.15 $Y=0.425
+ $X2=1.03 $Y2=0.425
r31 13 18 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.03 $Y=0.595
+ $X2=1.03 $Y2=0.425
r32 8 13 47.7707 $w=2.18e-07 $l=9e-07 $layer=LI1_cond $X=1.03 $Y=1.495 $X2=1.03
+ $Y2=0.595
r33 7 11 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=1.03 $Y=1.595
+ $X2=1.165 $Y2=1.595
r34 7 8 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.03 $Y=1.595 $X2=1.03
+ $Y2=1.495
r35 2 11 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.485 $X2=1.165 $Y2=1.61
r36 1 23 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
c62 16 0 1.5767e-19 $X=1.575 $Y=0.38
r63 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r64 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r65 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r66 42 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r67 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r68 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0 $X2=3
+ $Y2=0
r69 39 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.45
+ $Y2=0
r70 38 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r71 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r72 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 35 48 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.59
+ $Y2=0
r74 35 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.07
+ $Y2=0
r75 34 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0 $X2=3
+ $Y2=0
r76 34 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.07
+ $Y2=0
r77 33 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r78 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r79 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r80 30 45 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.685
+ $Y2=0
r81 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=1.15
+ $Y2=0
r82 29 48 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.59
+ $Y2=0
r83 29 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r84 24 45 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.685
+ $Y2=0
r85 24 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r86 22 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r87 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r88 18 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0
r89 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0.39
r90 14 48 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r91 14 16 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.38
r92 10 45 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.085
+ $X2=0.685 $Y2=0
r93 10 12 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.685 $Y=0.085
+ $X2=0.685 $Y2=0.66
r94 3 20 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3 $Y2=0.39
r95 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.38
r96 1 12 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.68 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HD__O21BA_2%A_478_47# 1 2 9 11 12 15
c28 11 0 1.44727e-19 $X=3.255 $Y=0.82
r29 13 15 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.422 $Y=0.735
+ $X2=3.422 $Y2=0.39
r30 11 13 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.255 $Y=0.82
+ $X2=3.422 $Y2=0.735
r31 11 12 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.255 $Y=0.82
+ $X2=2.745 $Y2=0.82
r32 7 12 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.595 $Y=0.735
+ $X2=2.745 $Y2=0.82
r33 7 9 5.95429 $w=2.98e-07 $l=1.55e-07 $layer=LI1_cond $X=2.595 $Y=0.735
+ $X2=2.595 $Y2=0.58
r34 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.235 $X2=3.42 $Y2=0.39
r35 1 9 182 $w=1.7e-07 $l=4.29622e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.58 $Y2=0.58
.ends


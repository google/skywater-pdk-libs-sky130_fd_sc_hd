# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__a2111oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 0.995000 2.725000 1.400000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.350000 3.090000 1.020000 ;
        RECT 2.905000 1.020000 3.540000 1.290000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.050000 2.270000 1.400000 ;
        RECT 1.940000 1.400000 2.215000 2.455000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.050000 1.770000 2.455000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785000 1.050000 1.235000 2.455000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.388750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.700000 1.375000 0.705000 ;
        RECT 0.145000 0.705000 2.420000 0.815000 ;
        RECT 0.145000 0.815000 2.300000 0.880000 ;
        RECT 0.145000 0.880000 0.530000 2.460000 ;
        RECT 1.045000 0.260000 1.375000 0.700000 ;
        RECT 2.090000 0.305000 2.420000 0.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.315000  0.085000 0.630000 0.525000 ;
        RECT 1.550000  0.085000 1.880000 0.535000 ;
        RECT 3.270000  0.085000 3.510000 0.760000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 2.800000 1.920000 3.130000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.395000 1.580000 3.505000 1.750000 ;
      RECT 2.395000 1.750000 2.625000 2.460000 ;
      RECT 3.310000 1.750000 3.505000 2.460000 ;
  END
END sky130_fd_sc_hd__a2111oi_1

* File: sky130_fd_sc_hd__edfxbp_1.spice
* Created: Tue Sep  1 19:07:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__edfxbp_1.pex.spice"
.subckt sky130_fd_sc_hd__edfxbp_1  VNB VPB CLK D DE VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* DE	DE
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_193_47#_M1015_d N_A_27_47#_M1015_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_381_47# N_D_M1002_g N_A_299_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_DE_M1004_g A_381_47# VNB NSHORT L=0.15 W=0.42 AD=0.1092
+ AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_DE_M1031_g N_A_423_343#_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1092 PD=0.71 PS=1.36 NRD=1.428 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1016 A_729_47# N_A_423_343#_M1016_g N_VGND_M1031_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0609 PD=0.78 PS=0.71 NRD=35.712 NRS=1.428 M=1 R=2.8 SA=75000.6
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1034 N_A_299_47#_M1034_d N_A_791_264#_M1034_g A_729_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.155723 AS=0.0756 PD=1.27077 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8
+ SA=75001.1 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_986_413#_M1005_d N_A_27_47#_M1005_g N_A_299_47#_M1034_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0522 AS=0.133477 PD=0.65 PS=1.08923 NRD=0 NRS=161.664 M=1
+ R=2.4 SA=75002 SB=75001.8 A=0.054 P=1.02 MULT=1
MM1030 A_1101_47# N_A_193_47#_M1030_g N_A_986_413#_M1005_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0700615 AS=0.0522 PD=0.738462 PS=0.65 NRD=46.536 NRS=4.992 M=1
+ R=2.4 SA=75002.5 SB=75001.3 A=0.054 P=1.02 MULT=1
MM1035 N_VGND_M1035_d N_A_1150_159#_M1035_g A_1101_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0958472 AS=0.0817385 PD=0.859811 PS=0.861538 NRD=0 NRS=39.888 M=1 R=2.8
+ SA=75002.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1022 N_A_1150_159#_M1022_d N_A_986_413#_M1022_g N_VGND_M1035_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.146053 PD=1.8 PS=1.31019 NRD=0 NRS=30.936 M=1
+ R=4.26667 SA=75002.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 A_1514_47# N_A_1150_159#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0730154 AS=0.1092 PD=0.813077 PS=1.36 NRD=33.948 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_1591_413#_M1003_d N_A_193_47#_M1003_g A_1514_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0684 AS=0.0625846 PD=0.74 PS=0.696923 NRD=3.324 NRS=39.612 M=1
+ R=2.4 SA=75000.7 SB=75001.7 A=0.054 P=1.02 MULT=1
MM1006 A_1717_47# N_A_27_47#_M1006_g N_A_1591_413#_M1003_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0684 PD=0.687692 PS=0.74 NRD=38.076 NRS=30 M=1 R=2.4
+ SA=75001.2 SB=75001.1 A=0.054 P=1.02 MULT=1
MM1019 N_VGND_M1019_d N_A_791_264#_M1019_g A_1717_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.0710769 PD=0.773271 PS=0.802308 NRD=17.136 NRS=32.628 M=1
+ R=2.8 SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_Q_N_M1023_d N_A_791_264#_M1023_g N_VGND_M1019_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.121799 PD=1.82 PS=1.19673 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A_1591_413#_M1020_g N_A_791_264#_M1020_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0787009 AS=0.1092 PD=0.773271 PS=1.36 NRD=17.136 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1024 N_Q_M1024_d N_A_1591_413#_M1024_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.121799 PD=1.86 PS=1.19673 NRD=0.912 NRS=0 M=1 R=4.33333
+ SA=75000.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_VPWR_M1013_d N_CLK_M1013_g N_A_27_47#_M1013_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_193_47#_M1000_d N_A_27_47#_M1000_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 A_381_369# N_D_M1021_g N_A_299_47#_M1021_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1664 PD=0.85 PS=1.8 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.5 A=0.096 P=1.58 MULT=1
MM1027 N_VPWR_M1027_d N_A_423_343#_M1027_g A_381_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1664 AS=0.0672 PD=1.8 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_DE_M1011_g N_A_423_343#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0928 AS=0.1664 PD=0.93 PS=1.8 NRD=1.5366 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1014 A_729_369# N_DE_M1014_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.0928 PD=1 PS=0.93 NRD=38.4741 NRS=1.5366 M=1 R=4.26667
+ SA=75000.6 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1029 N_A_299_47#_M1029_d N_A_791_264#_M1029_g A_729_369# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.193026 AS=0.1152 PD=1.52755 PS=1 NRD=0 NRS=38.4741 M=1 R=4.26667
+ SA=75001.1 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_986_413#_M1008_d N_A_193_47#_M1008_g N_A_299_47#_M1029_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.06405 AS=0.126674 PD=0.725 PS=1.00245 NRD=4.6886
+ NRS=165.322 M=1 R=2.8 SA=75001.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 A_1077_413# N_A_27_47#_M1009_g N_A_986_413#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.07665 AS=0.06405 PD=0.785 PS=0.725 NRD=59.7895 NRS=7.0329 M=1
+ R=2.8 SA=75002.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_1150_159#_M1001_g A_1077_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.128423 AS=0.07665 PD=0.904615 PS=0.785 NRD=97.318 NRS=59.7895 M=1
+ R=2.8 SA=75002.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1012 N_A_1150_159#_M1012_d N_A_986_413#_M1012_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.15 W=0.75 AD=0.195 AS=0.229327 PD=2.02 PS=1.61538 NRD=0 NRS=6.5601 M=1 R=5
+ SA=75002.1 SB=75000.2 A=0.1125 P=1.8 MULT=1
MM1025 A_1500_413# N_A_1150_159#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06405 AS=0.1092 PD=0.725 PS=1.36 NRD=45.7237 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1032 N_A_1591_413#_M1032_d N_A_27_47#_M1032_g A_1500_413# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0567 AS=0.06405 PD=0.69 PS=0.725 NRD=0 NRS=45.7237 M=1 R=2.8
+ SA=75000.6 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1026 A_1675_413# N_A_193_47#_M1026_g N_A_1591_413#_M1032_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0882 AS=0.0567 PD=0.84 PS=0.69 NRD=72.693 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_A_791_264#_M1018_g A_1675_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0862183 AS=0.0882 PD=0.789718 PS=0.84 NRD=29.3136 NRS=72.693 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_Q_N_M1007_d N_A_791_264#_M1007_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.205282 PD=2.52 PS=1.88028 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1028 N_VPWR_M1028_d N_A_1591_413#_M1028_g N_A_791_264#_M1028_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.120195 AS=0.1728 PD=1.04195 PS=1.82 NRD=18.4589 NRS=1.5366
+ M=1 R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1017 N_Q_M1017_d N_A_1591_413#_M1017_g N_VPWR_M1028_d VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.187805 PD=2.56 PS=1.62805 NRD=0.9653 NRS=0 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.8057 P=27.89
c_227 VPB 0 1.40584e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__edfxbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__lpflow_isobufsrc_8.pex.spice
* Created: Tue Sep  1 19:12:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A 3 5 7 10 12 14 17 27 31
r43 29 31 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=0.265 $Y=1.175
+ $X2=0.27 $Y2=1.175
r44 26 27 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.96 $Y=1.16 $X2=1.2
+ $Y2=1.16
r45 25 26 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.78 $Y=1.16 $X2=0.96
+ $Y2=1.16
r46 24 25 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.54 $Y=1.16
+ $X2=0.78 $Y2=1.16
r47 21 24 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.36 $Y=1.16 $X2=0.54
+ $Y2=1.16
r48 17 29 3.10749 $w=2.2e-07 $l=9e-08 $layer=LI1_cond $X=0.175 $Y=1.175
+ $X2=0.265 $Y2=1.175
r49 17 31 2.09535 $w=2.18e-07 $l=4e-08 $layer=LI1_cond $X=0.31 $Y=1.175 $X2=0.27
+ $Y2=1.175
r50 17 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r51 12 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=0.995
+ $X2=1.2 $Y2=1.16
r52 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.2 $Y=0.995 $X2=1.2
+ $Y2=0.56
r53 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.325
+ $X2=0.96 $Y2=1.16
r54 8 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.96 $Y=1.325
+ $X2=0.96 $Y2=1.985
r55 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=0.995
+ $X2=0.78 $Y2=1.16
r56 5 7 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.78 $Y=0.995 $X2=0.78
+ $Y2=0.56
r57 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.325
+ $X2=0.54 $Y2=1.16
r58 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.54 $Y=1.325 $X2=0.54
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_123_297# 1 2 7 9 12 14 16 19 21
+ 23 26 28 30 33 35 37 40 42 44 47 49 51 54 56 58 61 65 67 73 80 83 84 95
r176 92 93 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=4.06 $Y=1.16
+ $X2=4.48 $Y2=1.16
r177 91 92 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.64 $Y=1.16
+ $X2=4.06 $Y2=1.16
r178 90 91 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=3.22 $Y=1.16
+ $X2=3.64 $Y2=1.16
r179 89 90 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.8 $Y=1.16
+ $X2=3.22 $Y2=1.16
r180 88 89 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.38 $Y=1.16
+ $X2=2.8 $Y2=1.16
r181 81 95 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=4.9 $Y2=1.16
r182 81 93 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=4.79 $Y=1.16
+ $X2=4.48 $Y2=1.16
r183 80 81 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=4.79
+ $Y=1.16 $X2=4.79 $Y2=1.16
r184 78 88 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=2.07 $Y=1.16
+ $X2=2.38 $Y2=1.16
r185 78 85 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=2.07 $Y=1.16
+ $X2=1.96 $Y2=1.16
r186 77 80 143.654 $w=2.08e-07 $l=2.72e-06 $layer=LI1_cond $X=2.07 $Y=1.18
+ $X2=4.79 $Y2=1.18
r187 77 78 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r188 75 84 1.9773 $w=2.1e-07 $l=2.07485e-07 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=0.95 $Y2=1.175
r189 75 77 48.3247 $w=2.08e-07 $l=9.15e-07 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=2.07 $Y2=1.18
r190 71 84 4.45781 $w=2.5e-07 $l=1.28452e-07 $layer=LI1_cond $X=0.99 $Y=1.065
+ $X2=0.95 $Y2=1.175
r191 71 73 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.99 $Y=1.065
+ $X2=0.99 $Y2=0.39
r192 69 84 4.45781 $w=2.5e-07 $l=1.66132e-07 $layer=LI1_cond $X=0.83 $Y=1.285
+ $X2=0.95 $Y2=1.175
r193 69 83 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.83 $Y=1.285
+ $X2=0.83 $Y2=1.455
r194 65 83 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.62
+ $X2=0.75 $Y2=1.455
r195 65 67 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.75 $Y=1.62
+ $X2=0.75 $Y2=2.3
r196 59 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.325
+ $X2=4.9 $Y2=1.16
r197 59 61 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.9 $Y=1.325
+ $X2=4.9 $Y2=1.985
r198 56 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=1.16
r199 56 58 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=0.56
r200 52 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=1.325
+ $X2=4.48 $Y2=1.16
r201 52 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.48 $Y=1.325
+ $X2=4.48 $Y2=1.985
r202 49 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.48 $Y=0.995
+ $X2=4.48 $Y2=1.16
r203 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.48 $Y=0.995
+ $X2=4.48 $Y2=0.56
r204 45 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=1.325
+ $X2=4.06 $Y2=1.16
r205 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.06 $Y=1.325
+ $X2=4.06 $Y2=1.985
r206 42 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=1.16
r207 42 44 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.06 $Y=0.995
+ $X2=4.06 $Y2=0.56
r208 38 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.325
+ $X2=3.64 $Y2=1.16
r209 38 40 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.64 $Y=1.325
+ $X2=3.64 $Y2=1.985
r210 35 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=1.16
r211 35 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.64 $Y=0.995
+ $X2=3.64 $Y2=0.56
r212 31 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.325
+ $X2=3.22 $Y2=1.16
r213 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.22 $Y=1.325
+ $X2=3.22 $Y2=1.985
r214 28 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.22 $Y2=1.16
r215 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.22 $Y=0.995
+ $X2=3.22 $Y2=0.56
r216 24 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.325
+ $X2=2.8 $Y2=1.16
r217 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.8 $Y=1.325
+ $X2=2.8 $Y2=1.985
r218 21 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.995
+ $X2=2.8 $Y2=1.16
r219 21 23 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.8 $Y=0.995
+ $X2=2.8 $Y2=0.56
r220 17 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.325
+ $X2=2.38 $Y2=1.16
r221 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.38 $Y=1.325
+ $X2=2.38 $Y2=1.985
r222 14 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=0.995
+ $X2=2.38 $Y2=1.16
r223 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.38 $Y=0.995
+ $X2=2.38 $Y2=0.56
r224 10 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.325
+ $X2=1.96 $Y2=1.16
r225 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.96 $Y=1.325
+ $X2=1.96 $Y2=1.985
r226 7 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=0.995
+ $X2=1.96 $Y2=1.16
r227 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.96 $Y=0.995
+ $X2=1.96 $Y2=0.56
r228 2 67 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.485 $X2=0.75 $Y2=2.3
r229 2 65 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.485 $X2=0.75 $Y2=1.62
r230 1 73 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.855
+ $Y=0.235 $X2=0.99 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%SLEEP 1 3 6 8 10 13 15 17 20 22
+ 24 27 29 31 34 36 38 41 43 45 48 50 52 55 57 71 73
r143 72 73 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7.84 $Y=1.16
+ $X2=8.26 $Y2=1.16
r144 70 72 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.825 $Y=1.16
+ $X2=7.84 $Y2=1.16
r145 70 71 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=7.825
+ $Y=1.16 $X2=7.825 $Y2=1.16
r146 68 70 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=7.42 $Y=1.16
+ $X2=7.825 $Y2=1.16
r147 67 68 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=7 $Y=1.16 $X2=7.42
+ $Y2=1.16
r148 66 67 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.58 $Y=1.16 $X2=7
+ $Y2=1.16
r149 65 66 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.16 $Y=1.16
+ $X2=6.58 $Y2=1.16
r150 64 65 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.74 $Y=1.16
+ $X2=6.16 $Y2=1.16
r151 62 64 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.445 $Y=1.16
+ $X2=5.74 $Y2=1.16
r152 62 63 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=5.445
+ $Y=1.16 $X2=5.445 $Y2=1.16
r153 59 62 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.32 $Y=1.16
+ $X2=5.445 $Y2=1.16
r154 57 71 115.068 $w=1.98e-07 $l=2.075e-06 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=7.825 $Y2=1.175
r155 57 63 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.445 $Y2=1.175
r156 53 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=1.325
+ $X2=8.26 $Y2=1.16
r157 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.26 $Y=1.325
+ $X2=8.26 $Y2=1.985
r158 50 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=0.995
+ $X2=8.26 $Y2=1.16
r159 50 52 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.26 $Y=0.995
+ $X2=8.26 $Y2=0.56
r160 46 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.84 $Y=1.325
+ $X2=7.84 $Y2=1.16
r161 46 48 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.84 $Y=1.325
+ $X2=7.84 $Y2=1.985
r162 43 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.84 $Y=0.995
+ $X2=7.84 $Y2=1.16
r163 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.84 $Y=0.995
+ $X2=7.84 $Y2=0.56
r164 39 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.42 $Y=1.325
+ $X2=7.42 $Y2=1.16
r165 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.42 $Y=1.325
+ $X2=7.42 $Y2=1.985
r166 36 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.42 $Y=0.995
+ $X2=7.42 $Y2=1.16
r167 36 38 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.42 $Y=0.995
+ $X2=7.42 $Y2=0.56
r168 32 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.325 $X2=7
+ $Y2=1.16
r169 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7 $Y=1.325 $X2=7
+ $Y2=1.985
r170 29 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=0.995 $X2=7
+ $Y2=1.16
r171 29 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7 $Y=0.995 $X2=7
+ $Y2=0.56
r172 25 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.58 $Y=1.325
+ $X2=6.58 $Y2=1.16
r173 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.58 $Y=1.325
+ $X2=6.58 $Y2=1.985
r174 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=1.16
r175 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=0.56
r176 18 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.325
+ $X2=6.16 $Y2=1.16
r177 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.16 $Y=1.325
+ $X2=6.16 $Y2=1.985
r178 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.16
r179 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r180 11 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.325
+ $X2=5.74 $Y2=1.16
r181 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.74 $Y=1.325
+ $X2=5.74 $Y2=1.985
r182 8 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.16
r183 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r184 4 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.325
+ $X2=5.32 $Y2=1.16
r185 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.32 $Y=1.325
+ $X2=5.32 $Y2=1.985
r186 1 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.16
r187 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VPWR 1 2 3 4 5 6 19 21 25 29 33
+ 37 41 45 49 52 53 55 56 57 59 75 76 82 85 88
r124 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r125 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r128 75 76 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r129 73 76 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=8.51 $Y2=2.72
r130 72 75 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=8.51 $Y2=2.72
r131 72 73 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r132 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r133 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r134 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 67 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r136 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r137 64 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.01 $Y2=2.72
r138 64 66 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.135 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 63 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r140 63 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r142 60 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.17 $Y2=2.72
r143 60 62 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.295 $Y=2.72
+ $X2=2.53 $Y2=2.72
r144 59 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.885 $Y=2.72
+ $X2=3.01 $Y2=2.72
r145 59 62 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.885 $Y=2.72
+ $X2=2.53 $Y2=2.72
r146 57 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r147 57 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r148 55 69 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.37 $Y2=2.72
r149 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.69 $Y2=2.72
r150 54 72 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.83 $Y2=2.72
r151 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.815 $Y=2.72
+ $X2=4.69 $Y2=2.72
r152 52 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.45 $Y2=2.72
r153 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=2.72
+ $X2=3.85 $Y2=2.72
r154 51 69 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=4.37 $Y2=2.72
r155 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.975 $Y=2.72
+ $X2=3.85 $Y2=2.72
r156 47 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=2.635
+ $X2=4.69 $Y2=2.72
r157 47 49 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.69 $Y=2.635
+ $X2=4.69 $Y2=2
r158 43 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2.72
r159 43 45 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.85 $Y=2.635
+ $X2=3.85 $Y2=2
r160 39 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=2.635
+ $X2=3.01 $Y2=2.72
r161 39 41 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.01 $Y=2.635
+ $X2=3.01 $Y2=2
r162 35 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.72
r163 35 37 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2
r164 34 82 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.33 $Y=2.72
+ $X2=1.207 $Y2=2.72
r165 33 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=2.72
+ $X2=2.17 $Y2=2.72
r166 33 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.045 $Y=2.72
+ $X2=1.33 $Y2=2.72
r167 29 32 32.9269 $w=2.43e-07 $l=7e-07 $layer=LI1_cond $X=1.207 $Y=1.64
+ $X2=1.207 $Y2=2.34
r168 27 82 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.207 $Y=2.635
+ $X2=1.207 $Y2=2.72
r169 27 32 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.207 $Y=2.635
+ $X2=1.207 $Y2=2.34
r170 26 79 3.70423 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.207 $Y2=2.72
r171 25 82 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=1.207 $Y2=2.72
r172 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.085 $Y=2.72
+ $X2=0.415 $Y2=2.72
r173 21 24 36.6686 $w=2.18e-07 $l=7e-07 $layer=LI1_cond $X=0.305 $Y=1.64
+ $X2=0.305 $Y2=2.34
r174 19 79 3.25901 $w=2.2e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.207 $Y2=2.72
r175 19 24 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.305 $Y=2.635
+ $X2=0.305 $Y2=2.34
r176 6 49 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.555
+ $Y=1.485 $X2=4.69 $Y2=2
r177 5 45 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=3.715
+ $Y=1.485 $X2=3.85 $Y2=2
r178 4 41 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.875
+ $Y=1.485 $X2=3.01 $Y2=2
r179 3 37 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.035
+ $Y=1.485 $X2=2.17 $Y2=2
r180 2 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.485 $X2=1.17 $Y2=2.34
r181 2 29 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.485 $X2=1.17 $Y2=1.64
r182 1 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.485 $X2=0.33 $Y2=2.34
r183 1 21 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.485 $X2=0.33 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%A_321_297# 1 2 3 4 5 6 7 8 9 28
+ 30 32 36 38 42 44 48 50 52 53 54 58 60 64 66 70 72 76 81 83 85 90 91 92
r104 74 76 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.47 $Y=2.295
+ $X2=8.47 $Y2=1.96
r105 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.755 $Y=2.38
+ $X2=7.63 $Y2=2.38
r106 72 74 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.345 $Y=2.38
+ $X2=8.47 $Y2=2.295
r107 72 73 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.345 $Y=2.38
+ $X2=7.755 $Y2=2.38
r108 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=2.295
+ $X2=7.63 $Y2=2.38
r109 68 70 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.63 $Y=2.295
+ $X2=7.63 $Y2=1.96
r110 67 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.915 $Y=2.38
+ $X2=6.79 $Y2=2.38
r111 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.505 $Y=2.38
+ $X2=7.63 $Y2=2.38
r112 66 67 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.505 $Y=2.38
+ $X2=6.915 $Y2=2.38
r113 62 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.79 $Y=2.295
+ $X2=6.79 $Y2=2.38
r114 62 64 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.79 $Y=2.295
+ $X2=6.79 $Y2=1.96
r115 61 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.075 $Y=2.38
+ $X2=5.95 $Y2=2.38
r116 60 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.665 $Y=2.38
+ $X2=6.79 $Y2=2.38
r117 60 61 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.665 $Y=2.38
+ $X2=6.075 $Y2=2.38
r118 56 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.295
+ $X2=5.95 $Y2=2.38
r119 56 58 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.95 $Y=2.295
+ $X2=5.95 $Y2=1.96
r120 55 89 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.235 $Y=2.38
+ $X2=5.11 $Y2=2.38
r121 54 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=2.38
+ $X2=5.95 $Y2=2.38
r122 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.825 $Y=2.38
+ $X2=5.235 $Y2=2.38
r123 53 89 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=2.295
+ $X2=5.11 $Y2=2.38
r124 52 87 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.11 $Y=1.665
+ $X2=5.11 $Y2=1.56
r125 52 53 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=5.11 $Y=1.665
+ $X2=5.11 $Y2=2.295
r126 51 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.395 $Y=1.56
+ $X2=4.27 $Y2=1.56
r127 50 87 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.985 $Y=1.56
+ $X2=5.11 $Y2=1.56
r128 50 51 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.985 $Y=1.56
+ $X2=4.395 $Y2=1.56
r129 46 85 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.27 $Y=1.665
+ $X2=4.27 $Y2=1.56
r130 46 48 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.27 $Y=1.665
+ $X2=4.27 $Y2=2.3
r131 45 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.555 $Y=1.56
+ $X2=3.43 $Y2=1.56
r132 44 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.145 $Y=1.56
+ $X2=4.27 $Y2=1.56
r133 44 45 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.145 $Y=1.56
+ $X2=3.555 $Y2=1.56
r134 40 83 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.43 $Y=1.665
+ $X2=3.43 $Y2=1.56
r135 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.43 $Y=1.665
+ $X2=3.43 $Y2=2.3
r136 39 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.715 $Y=1.56
+ $X2=2.59 $Y2=1.56
r137 38 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.305 $Y=1.56
+ $X2=3.43 $Y2=1.56
r138 38 39 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=3.305 $Y=1.56
+ $X2=2.715 $Y2=1.56
r139 34 81 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.59 $Y=1.665
+ $X2=2.59 $Y2=1.56
r140 34 36 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.59 $Y=1.665
+ $X2=2.59 $Y2=2.3
r141 33 79 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=1.875 $Y=1.56
+ $X2=1.715 $Y2=1.56
r142 32 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.465 $Y=1.56
+ $X2=2.59 $Y2=1.56
r143 32 33 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=2.465 $Y=1.56
+ $X2=1.875 $Y2=1.56
r144 28 79 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=1.665
+ $X2=1.715 $Y2=1.56
r145 28 30 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=1.715 $Y=1.665
+ $X2=1.715 $Y2=2.3
r146 9 76 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=8.335
+ $Y=1.485 $X2=8.47 $Y2=1.96
r147 8 70 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=1.485 $X2=7.63 $Y2=1.96
r148 7 64 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.655
+ $Y=1.485 $X2=6.79 $Y2=1.96
r149 6 58 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.815
+ $Y=1.485 $X2=5.95 $Y2=1.96
r150 5 89 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.485 $X2=5.11 $Y2=2.3
r151 5 87 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.485 $X2=5.11 $Y2=1.62
r152 4 85 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.27 $Y2=1.62
r153 4 48 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.27 $Y2=2.3
r154 3 83 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.485 $X2=3.43 $Y2=1.62
r155 3 42 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.485 $X2=3.43 $Y2=2.3
r156 2 81 400 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.485 $X2=2.59 $Y2=1.62
r157 2 36 400 $w=1.7e-07 $l=8.79915e-07 $layer=licon1_PDIFF $count=1 $X=2.455
+ $Y=1.485 $X2=2.59 $Y2=2.3
r158 1 79 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.485 $X2=1.75 $Y2=1.62
r159 1 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.485 $X2=1.75 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%X 1 2 3 4 5 6 7 8 9 10 11 12 39
+ 41 42 45 47 51 53 57 59 63 67 69 70 71 75 79 81 83 87 91 93 95 99 103 105 106
+ 107 108 109 110 111 112 114 115
r224 113 115 10.4916 $w=6.43e-07 $l=5.4e-07 $layer=LI1_cond $X=8.417 $Y=0.905
+ $X2=8.417 $Y2=1.445
r225 113 114 2.53538 $w=4.02e-07 $l=1.86652e-07 $layer=LI1_cond $X=8.417
+ $Y=0.905 $X2=8.27 $Y2=0.815
r226 101 115 2.64909 $w=3.62e-07 $l=2.79285e-07 $layer=LI1_cond $X=8.05 $Y=1.615
+ $X2=8.29 $Y2=1.53
r227 101 103 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.05 $Y=1.615
+ $X2=8.05 $Y2=1.62
r228 97 114 2.53538 $w=4.02e-07 $l=2.61151e-07 $layer=LI1_cond $X=8.05 $Y=0.725
+ $X2=8.27 $Y2=0.815
r229 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.05 $Y=0.725
+ $X2=8.05 $Y2=0.39
r230 96 111 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=0.815
+ $X2=7.21 $Y2=0.815
r231 95 114 4.34862 $w=1.8e-07 $l=3.85e-07 $layer=LI1_cond $X=7.885 $Y=0.815
+ $X2=8.27 $Y2=0.815
r232 95 96 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.885 $Y=0.815
+ $X2=7.375 $Y2=0.815
r233 94 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=1.53
+ $X2=7.21 $Y2=1.53
r234 93 115 4.16724 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=7.925 $Y=1.53
+ $X2=8.29 $Y2=1.53
r235 93 94 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.925 $Y=1.53
+ $X2=7.335 $Y2=1.53
r236 89 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.21 $Y=1.615
+ $X2=7.21 $Y2=1.53
r237 89 91 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=7.21 $Y=1.615
+ $X2=7.21 $Y2=1.62
r238 85 111 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.21 $Y=0.725
+ $X2=7.21 $Y2=0.815
r239 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.21 $Y=0.725
+ $X2=7.21 $Y2=0.39
r240 84 109 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=0.815
+ $X2=6.37 $Y2=0.815
r241 83 111 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.045 $Y=0.815
+ $X2=7.21 $Y2=0.815
r242 83 84 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=7.045 $Y=0.815
+ $X2=6.535 $Y2=0.815
r243 82 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.495 $Y=1.53
+ $X2=6.37 $Y2=1.53
r244 81 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.085 $Y=1.53
+ $X2=7.21 $Y2=1.53
r245 81 82 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.085 $Y=1.53
+ $X2=6.495 $Y2=1.53
r246 77 110 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.37 $Y=1.615
+ $X2=6.37 $Y2=1.53
r247 77 79 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.37 $Y=1.615
+ $X2=6.37 $Y2=1.62
r248 73 109 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.37 $Y=0.725
+ $X2=6.37 $Y2=0.815
r249 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.37 $Y=0.725
+ $X2=6.37 $Y2=0.39
r250 72 108 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=0.815
+ $X2=5.53 $Y2=0.815
r251 71 109 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0.815
+ $X2=6.37 $Y2=0.815
r252 71 72 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=6.205 $Y=0.815
+ $X2=5.695 $Y2=0.815
r253 69 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.245 $Y=1.53
+ $X2=6.37 $Y2=1.53
r254 69 70 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.245 $Y=1.53
+ $X2=5.655 $Y2=1.53
r255 65 70 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.53 $Y=1.615
+ $X2=5.655 $Y2=1.53
r256 65 67 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.53 $Y=1.615
+ $X2=5.53 $Y2=1.62
r257 61 108 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.53 $Y=0.725
+ $X2=5.53 $Y2=0.815
r258 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.53 $Y=0.725
+ $X2=5.53 $Y2=0.39
r259 60 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=0.815
+ $X2=4.69 $Y2=0.815
r260 59 108 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=0.815
+ $X2=5.53 $Y2=0.815
r261 59 60 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=5.365 $Y=0.815
+ $X2=4.855 $Y2=0.815
r262 55 107 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.69 $Y=0.725
+ $X2=4.69 $Y2=0.815
r263 55 57 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.69 $Y=0.725
+ $X2=4.69 $Y2=0.39
r264 54 106 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0.815
+ $X2=3.85 $Y2=0.815
r265 53 107 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=0.815
+ $X2=4.69 $Y2=0.815
r266 53 54 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=4.525 $Y=0.815
+ $X2=4.015 $Y2=0.815
r267 49 106 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.85 $Y=0.725
+ $X2=3.85 $Y2=0.815
r268 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.85 $Y=0.725
+ $X2=3.85 $Y2=0.39
r269 48 105 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0.815
+ $X2=3.01 $Y2=0.815
r270 47 106 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0.815
+ $X2=3.85 $Y2=0.815
r271 47 48 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.685 $Y=0.815
+ $X2=3.175 $Y2=0.815
r272 43 105 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.01 $Y=0.725
+ $X2=3.01 $Y2=0.815
r273 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.01 $Y=0.725
+ $X2=3.01 $Y2=0.39
r274 41 105 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=0.815
+ $X2=3.01 $Y2=0.815
r275 41 42 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.845 $Y=0.815
+ $X2=2.335 $Y2=0.815
r276 37 42 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.17 $Y=0.725
+ $X2=2.335 $Y2=0.815
r277 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.17 $Y=0.725
+ $X2=2.17 $Y2=0.39
r278 12 103 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=7.915
+ $Y=1.485 $X2=8.05 $Y2=1.62
r279 11 91 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=7.075
+ $Y=1.485 $X2=7.21 $Y2=1.62
r280 10 79 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=6.235
+ $Y=1.485 $X2=6.37 $Y2=1.62
r281 9 67 300 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.485 $X2=5.53 $Y2=1.62
r282 8 99 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.915
+ $Y=0.235 $X2=8.05 $Y2=0.39
r283 7 87 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.075
+ $Y=0.235 $X2=7.21 $Y2=0.39
r284 6 75 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.235
+ $Y=0.235 $X2=6.37 $Y2=0.39
r285 5 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.39
r286 4 57 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.555
+ $Y=0.235 $X2=4.69 $Y2=0.39
r287 3 51 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.715
+ $Y=0.235 $X2=3.85 $Y2=0.39
r288 2 45 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.875
+ $Y=0.235 $X2=3.01 $Y2=0.39
r289 1 39 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.035
+ $Y=0.235 $X2=2.17 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HD__LPFLOW_ISOBUFSRC_8%VGND 1 2 3 4 5 6 7 8 9 10 33 37
+ 39 43 47 51 55 59 63 65 69 71 73 76 77 79 80 82 83 85 86 88 89 90 91 92 98 118
+ 124 127 130 134
r160 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r161 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r162 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r163 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=2.53 $Y2=0
r164 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r165 122 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r166 122 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r167 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r168 119 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.63 $Y2=0
r169 119 121 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=8.05 $Y2=0
r170 118 133 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=8.385 $Y=0
+ $X2=8.562 $Y2=0
r171 118 121 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.385 $Y=0
+ $X2=8.05 $Y2=0
r172 117 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r173 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r174 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r175 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r176 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r177 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r178 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r179 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r180 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r181 105 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.53 $Y2=0
r182 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r183 102 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0
+ $X2=2.59 $Y2=0
r184 102 104 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.675 $Y=0
+ $X2=2.99 $Y2=0
r185 101 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r186 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r187 98 124 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.58 $Y2=0
r188 98 100 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.15 $Y2=0
r189 92 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r190 92 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r191 90 116 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.67 $Y2=0
r192 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.705 $Y=0 $X2=6.79
+ $Y2=0
r193 88 113 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.865 $Y=0
+ $X2=5.75 $Y2=0
r194 88 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.95
+ $Y2=0
r195 87 116 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.035 $Y=0
+ $X2=6.67 $Y2=0
r196 87 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.035 $Y=0 $X2=5.95
+ $Y2=0
r197 85 110 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=4.83 $Y2=0
r198 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=0 $X2=5.11
+ $Y2=0
r199 84 113 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.195 $Y=0
+ $X2=5.75 $Y2=0
r200 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.11
+ $Y2=0
r201 82 107 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=3.91 $Y2=0
r202 82 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.27
+ $Y2=0
r203 81 110 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=4.83 $Y2=0
r204 81 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.27
+ $Y2=0
r205 79 104 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=2.99 $Y2=0
r206 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=0 $X2=3.43
+ $Y2=0
r207 78 107 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.515 $Y=0
+ $X2=3.91 $Y2=0
r208 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.43
+ $Y2=0
r209 76 95 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.23 $Y2=0
r210 76 77 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.545
+ $Y2=0
r211 75 100 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=0.655 $Y=0
+ $X2=1.15 $Y2=0
r212 75 77 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.655 $Y=0 $X2=0.545
+ $Y2=0
r213 71 133 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=8.52 $Y=0.085
+ $X2=8.562 $Y2=0
r214 71 73 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.52 $Y=0.085
+ $X2=8.52 $Y2=0.39
r215 67 130 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=0.085
+ $X2=7.63 $Y2=0
r216 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.63 $Y=0.085
+ $X2=7.63 $Y2=0.39
r217 66 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=0 $X2=6.79
+ $Y2=0
r218 65 130 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=0 $X2=7.63
+ $Y2=0
r219 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=6.875 $Y2=0
r220 61 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.79 $Y=0.085
+ $X2=6.79 $Y2=0
r221 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.79 $Y=0.085
+ $X2=6.79 $Y2=0.39
r222 57 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0
r223 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0.39
r224 53 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0
r225 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0.39
r226 49 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r227 49 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.39
r228 45 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0
r229 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.43 $Y=0.085
+ $X2=3.43 $Y2=0.39
r230 41 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r231 41 43 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.39
r232 40 124 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=1.58 $Y2=0
r233 39 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.59
+ $Y2=0
r234 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.505 $Y=0
+ $X2=1.835 $Y2=0
r235 35 124 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r236 35 37 7.15302 $w=5.08e-07 $l=3.05e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.39
r237 31 77 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=0.085
+ $X2=0.545 $Y2=0
r238 31 33 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0.085
+ $X2=0.545 $Y2=0.39
r239 10 73 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.335
+ $Y=0.235 $X2=8.47 $Y2=0.39
r240 9 69 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.495
+ $Y=0.235 $X2=7.63 $Y2=0.39
r241 8 63 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.79 $Y2=0.39
r242 7 59 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.39
r243 6 55 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.235 $X2=5.11 $Y2=0.39
r244 5 51 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.135
+ $Y=0.235 $X2=4.27 $Y2=0.39
r245 4 47 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.235 $X2=3.43 $Y2=0.39
r246 3 43 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.455
+ $Y=0.235 $X2=2.59 $Y2=0.39
r247 2 37 45.5 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_NDIFF $count=4 $X=1.275
+ $Y=0.235 $X2=1.75 $Y2=0.39
r248 1 33 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.445
+ $Y=0.235 $X2=0.57 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__o22a_4.spice
* Created: Thu Aug 27 14:37:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o22a_4.spice.pex"
.subckt sky130_fd_sc_hd__o22a_4  VNB VPB B1 B2 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_X_M1000_d N_A_96_21#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1004 N_X_M1000_d N_A_96_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_96_21#_M1005_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1017 N_X_M1005_d N_A_96_21#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1022 N_A_96_21#_M1022_d N_B1_M1022_g N_A_484_47#_M1022_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_96_21#_M1022_d N_B2_M1001_g N_A_484_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.8 A=0.0975 P=1.6 MULT=1
MM1018 N_A_96_21#_M1018_d N_B2_M1018_g N_A_484_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1023 N_A_96_21#_M1018_d N_B1_M1023_g N_A_484_47#_M1023_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.11375 PD=0.92 PS=1 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75001.4 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1012 N_A_484_47#_M1023_s N_A1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.08775 PD=1 PS=0.92 NRD=5.532 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1014 N_A_484_47#_M1014_d N_A2_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1015 N_A_484_47#_M1014_d N_A2_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1016 N_A_484_47#_M1016_d N_A1_M1016_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_96_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.4 A=0.15 P=2.3 MULT=1
MM1006 N_VPWR_M1006_d N_A_96_21#_M1006_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75005 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1006_d N_A_96_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.6 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A_96_21#_M1019_g N_X_M1007_s VPB PHIGHVT L=0.15 W=1
+ AD=0.395 AS=0.135 PD=1.79 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75004.2 A=0.15 P=2.3 MULT=1
MM1013 N_A_566_297#_M1013_d N_B1_M1013_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.395 PD=1.27 PS=1.79 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1009 N_A_566_297#_M1013_d N_B2_M1009_g N_A_96_21#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1010 N_A_566_297#_M1010_d N_B2_M1010_g N_A_96_21#_M1009_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1021 N_A_566_297#_M1010_d N_B1_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.7
+ SB=75002 A=0.15 P=2.3 MULT=1
MM1002 N_A_918_297#_M1002_d N_A1_M1002_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.175 PD=1.27 PS=1.35 NRD=0 NRS=14.7553 M=1 R=6.66667 SA=75004.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1011 N_A_918_297#_M1002_d N_A2_M1011_g N_A_96_21#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75004.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1020 N_A_918_297#_M1020_d N_A2_M1020_g N_A_96_21#_M1011_s VPB PHIGHVT L=0.15
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75005
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_918_297#_M1020_d N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.285 PD=1.27 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.4
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hd__o22a_4.spice.SKY130_FD_SC_HD__O22A_4.pxi"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 Y B1 VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=3.927e+11p ps=4.39e+06u
M1001 a_313_369# B1 a_241_369# VPB phighvt w=640000u l=150000u
+  ad=3.744e+11p pd=3.73e+06u as=1.344e+11p ps=1.7e+06u
M1002 VGND C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_427_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VGND A2 a_427_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_313_369# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1006 a_241_369# C1 a_169_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1007 a_169_369# D1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.888e+11p ps=1.87e+06u
M1008 Y D1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_313_369# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

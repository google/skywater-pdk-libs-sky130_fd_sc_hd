* File: sky130_fd_sc_hd__fahcon_1.spice
* Created: Tue Sep  1 19:09:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__fahcon_1.pex.spice"
.subckt sky130_fd_sc_hd__fahcon_1  VNB VPB A B CI VPWR COUT_N SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT_N	COUT_N
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_67_199#_M1012_g N_A_28_47#_M1012_s VNB NSHORT L=0.15
+ W=0.64 AD=0.104434 AS=0.1664 PD=0.967442 PS=1.8 NRD=4.68 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1023 N_A_67_199#_M1023_d N_A_M1023_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.323715 AS=0.106066 PD=1.65775 PS=0.982558 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_434_49#_M1009_d N_B_M1009_g N_A_67_199#_M1023_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.318735 PD=0.91 PS=1.63225 NRD=0 NRS=67.02 M=1 R=4.26667
+ SA=75001.8 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_28_47#_M1002_d N_A_488_21#_M1002_g N_A_434_49#_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2176 AS=0.0864 PD=1.96 PS=0.91 NRD=14.052 NRS=0 M=1
+ R=4.26667 SA=75002.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1015 N_A_726_47#_M1015_d N_A_488_21#_M1015_g N_A_67_199#_M1015_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.165675 AS=0.1792 PD=1.165 PS=1.84 NRD=44.988 NRS=2.808 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1031 N_A_28_47#_M1031_d N_B_M1031_g N_A_726_47#_M1015_d VNB NSHORT L=0.15
+ W=0.64 AD=0.16285 AS=0.165675 PD=1.8 PS=1.165 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1027 N_VGND_M1027_d N_B_M1027_g N_A_488_21#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.110903 AS=0.16715 PD=0.997674 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1005 N_A_1144_49#_M1005_d N_B_M1005_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1664 AS=0.109197 PD=1.8 PS=0.982326 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_COUT_N_M1013_d N_A_434_49#_M1013_g N_A_1261_49#_M1013_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.088 AS=0.1664 PD=0.915 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1029 N_A_1144_49#_M1029_d N_A_726_47#_M1029_g N_COUT_N_M1013_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1952 AS=0.088 PD=1.89 PS=0.915 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_1710_49#_M1007_d N_A_726_47#_M1007_g N_A_1589_49#_M1007_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.0928 AS=0.2912 PD=0.93 PS=2.19 NRD=2.808 NRS=29.052 M=1
+ R=4.26667 SA=75000.4 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_1634_315#_M1008_d N_A_434_49#_M1008_g N_A_1710_49#_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3136 AS=0.0928 PD=1.62 PS=0.93 NRD=130.308 NRS=0 M=1
+ R=4.26667 SA=75000.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A_1589_49#_M1020_g N_A_1634_315#_M1008_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.104434 AS=0.3136 PD=0.967442 PS=1.62 NRD=4.68 NRS=0.936 M=1
+ R=4.26667 SA=75001.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_1589_49#_M1003_d N_CI_M1003_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.106066 PD=1.82 PS=0.982558 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75002.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1026_d N_CI_M1026_g N_A_1261_49#_M1026_s VNB NSHORT L=0.15 W=0.64
+ AD=0.104434 AS=0.1664 PD=0.967442 PS=1.8 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1006 N_SUM_M1006_d N_A_1710_49#_M1006_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.65 AD=0.17875 AS=0.106066 PD=1.85 PS=0.982558 NRD=1.836 NRS=9.228 M=1
+ R=4.33333 SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1018 N_VPWR_M1018_d N_A_67_199#_M1018_g N_A_28_47#_M1018_s VPB PHIGHVT L=0.15
+ W=1 AD=0.175 AS=0.26 PD=1.35 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1017 N_A_67_199#_M1017_d N_A_M1017_g N_VPWR_M1018_d VPB PHIGHVT L=0.15 W=1
+ AD=0.3184 AS=0.175 PD=2.88 PS=1.35 NRD=34.4553 NRS=14.7553 M=1 R=6.66667
+ SA=75000.7 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1028 N_A_434_49#_M1028_d N_B_M1028_g N_A_28_47#_M1028_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1134 AS=0.2629 PD=1.11 PS=2.64 NRD=0 NRS=18.7544 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_A_67_199#_M1010_d N_A_488_21#_M1010_g N_A_434_49#_M1028_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2184 AS=0.1134 PD=2.2 PS=1.11 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 N_A_726_47#_M1014_d N_A_488_21#_M1014_g N_A_28_47#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.151637 AS=0.3314 PD=1.3 PS=2.75 NRD=0 NRS=12.3125 M=1 R=5.6
+ SA=75000.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_67_199#_M1019_d N_B_M1019_g N_A_726_47#_M1014_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2352 AS=0.151637 PD=2.24 PS=1.3 NRD=0 NRS=14.0658 M=1 R=5.6
+ SA=75000.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_488_21#_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.18 AS=0.26 PD=1.36 PS=2.52 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1001 N_A_1144_49#_M1001_d N_B_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.41587 AS=0.18 PD=1.94565 PS=1.36 NRD=50.2153 NRS=0 M=1 R=6.66667
+ SA=75000.7 SB=75001.6 A=0.15 P=2.3 MULT=1
MM1025 N_COUT_N_M1025_d N_A_434_49#_M1025_g N_A_1144_49#_M1001_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1134 AS=0.34933 PD=1.11 PS=1.63435 NRD=0 NRS=59.7895 M=1
+ R=5.6 SA=75001.6 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1004 N_A_1261_49#_M1004_d N_A_726_47#_M1004_g N_COUT_N_M1025_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.4536 AS=0.1134 PD=2.76 PS=1.11 NRD=59.7895 NRS=0 M=1 R=5.6
+ SA=75002.1 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1024 N_A_1710_49#_M1024_d N_A_726_47#_M1024_g N_A_1634_315#_M1024_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1022 N_A_1589_49#_M1022_d N_A_434_49#_M1022_g N_A_1710_49#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3024 AS=0.1134 PD=2.4 PS=1.11 NRD=17.5724 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1030 N_VPWR_M1030_d N_A_1589_49#_M1030_g N_A_1634_315#_M1030_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.135 AS=0.35 PD=1.27 PS=2.7 NRD=0 NRS=7.8603 M=1 R=6.66667
+ SA=75000.3 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_1589_49#_M1016_d N_CI_M1016_g N_VPWR_M1030_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.7
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1021 N_VPWR_M1021_d N_CI_M1021_g N_A_1261_49#_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1011 N_SUM_M1011_d N_A_1710_49#_M1011_g N_VPWR_M1021_d VPB PHIGHVT L=0.15 W=1
+ AD=0.285 AS=0.135 PD=2.57 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.544 P=28.81
pX33_noxref noxref_20 B B PROBETYPE=1
c_208 VPB 0 1.11799e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__fahcon_1.pxi.spice"
*
.ends
*
*

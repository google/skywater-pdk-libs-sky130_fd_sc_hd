# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.900000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.075000 2.690000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.075000 4.300000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 0.255000 1.285000 0.725000 ;
        RECT 0.955000 0.725000 6.760000 0.905000 ;
        RECT 1.795000 0.255000 2.125000 0.725000 ;
        RECT 3.155000 0.255000 3.485000 0.725000 ;
        RECT 3.995000 0.255000 4.325000 0.725000 ;
        RECT 4.835000 0.255000 5.165000 0.725000 ;
        RECT 4.875000 1.455000 6.760000 1.625000 ;
        RECT 4.875000 1.625000 5.125000 2.125000 ;
        RECT 5.675000 0.255000 6.005000 0.725000 ;
        RECT 5.715000 1.625000 5.965000 2.125000 ;
        RECT 6.420000 0.905000 6.760000 1.455000 ;
        RECT 6.515000 0.315000 6.760000 0.725000 ;
        RECT 6.555000 1.625000 6.760000 2.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.900000 0.085000 ;
        RECT 0.615000  0.085000 0.785000 0.555000 ;
        RECT 1.455000  0.085000 1.625000 0.555000 ;
        RECT 2.295000  0.085000 2.985000 0.555000 ;
        RECT 3.655000  0.085000 3.825000 0.555000 ;
        RECT 4.495000  0.085000 4.665000 0.555000 ;
        RECT 5.335000  0.085000 5.505000 0.555000 ;
        RECT 6.175000  0.085000 6.345000 0.555000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.900000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.900000 2.805000 ;
        RECT 0.575000 1.795000 0.825000 2.635000 ;
        RECT 1.415000 2.135000 1.665000 2.635000 ;
        RECT 2.255000 2.135000 2.505000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.900000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.255000 0.445000 0.735000 ;
      RECT 0.110000 0.735000 0.785000 0.905000 ;
      RECT 0.110000 1.455000 4.705000 1.625000 ;
      RECT 0.110000 1.625000 0.405000 2.465000 ;
      RECT 0.615000 0.905000 0.785000 1.455000 ;
      RECT 0.995000 1.795000 4.285000 1.965000 ;
      RECT 0.995000 1.965000 1.245000 2.465000 ;
      RECT 1.835000 1.965000 2.085000 2.465000 ;
      RECT 2.775000 2.135000 3.025000 2.295000 ;
      RECT 2.775000 2.295000 6.385000 2.465000 ;
      RECT 3.195000 1.965000 3.445000 2.125000 ;
      RECT 3.615000 2.135000 3.865000 2.295000 ;
      RECT 4.035000 1.965000 4.285000 2.125000 ;
      RECT 4.455000 1.795000 4.705000 2.295000 ;
      RECT 4.535000 1.075000 6.125000 1.285000 ;
      RECT 4.535000 1.285000 4.705000 1.455000 ;
      RECT 5.295000 1.795000 5.545000 2.295000 ;
      RECT 6.135000 1.795000 6.385000 2.295000 ;
  END
END sky130_fd_sc_hd__nor3b_4
END LIBRARY

* File: sky130_fd_sc_hd__or3_4.spice
* Created: Tue Sep  1 19:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__or3_4.pex.spice"
.subckt sky130_fd_sc_hd__or3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_C_M1012_g N_A_27_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_B_M1004_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_27_47#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.26 AS=0.08775 PD=1.45 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1007_d N_A_27_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26 AS=0.08775 PD=1.45 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_27_47#_M1010_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1011 N_VGND_M1010_d N_A_27_47#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A_27_47#_M1013_g N_X_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.08775 PD=1.93 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 A_109_297# N_C_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=15.7403 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75003.3
+ A=0.15 P=2.3 MULT=1
MM1002 A_193_297# N_B_M1002_g A_109_297# VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=15.7403 NRS=15.7403 M=1 R=6.66667 SA=75000.6
+ SB=75002.9 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_193_297# VPB PHIGHVT L=0.15 W=1 AD=0.4
+ AS=0.135 PD=1.8 PS=1.27 NRD=11.8003 NRS=15.7403 M=1 R=6.66667 SA=75001
+ SB=75002.5 A=0.15 P=2.3 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.4 PD=1.27 PS=1.8 NRD=0 NRS=0 M=1 R=6.66667 SA=75002 SB=75001.5
+ A=0.15 P=2.3 MULT=1
MM1003 N_X_M1001_d N_A_27_47#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.4
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.7 A=0.15 P=2.3 MULT=1
MM1006 N_X_M1005_d N_A_27_47#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.36 PD=1.27 PS=2.72 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75000.3 A=0.15 P=2.3 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__or3_4.pxi.spice"
*
.ends
*
*

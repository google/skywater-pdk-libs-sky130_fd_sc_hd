* File: sky130_fd_sc_hd__a211o_4.spice
* Created: Thu Aug 27 13:59:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a211o_4.spice.pex"
.subckt sky130_fd_sc_hd__a211o_4  VNB VPB B1 C1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_79_204#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75005.3 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1003_d N_A_79_204#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1013_d N_A_79_204#_M1013_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.091 PD=0.945 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1022 N_X_M1013_d N_A_79_204#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.095875 AS=0.092625 PD=0.945 PS=0.935 NRD=2.76 NRS=0.912 M=1 R=4.33333
+ SA=75001.5 SB=75004 A=0.0975 P=1.6 MULT=1
MM1014 N_A_79_204#_M1014_d N_B1_M1014_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.092625 PD=0.97 PS=0.935 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1002 N_A_79_204#_M1014_d N_C1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.108875 PD=0.97 PS=0.985 NRD=7.38 NRS=2.76 M=1 R=4.33333
+ SA=75002.4 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1007 N_A_79_204#_M1007_d N_C1_M1007_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.108875 PD=1.04 PS=0.985 NRD=11.076 NRS=7.38 M=1 R=4.33333
+ SA=75002.9 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_79_204#_M1007_d N_B1_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12675 AS=0.13975 PD=1.04 PS=1.08 NRD=9.228 NRS=7.38 M=1 R=4.33333
+ SA=75003.4 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1017_s N_A2_M1005_g A_951_47# VNB NSHORT L=0.15 W=0.65 AD=0.13975
+ AS=0.091 PD=1.08 PS=0.93 NRD=20.304 NRS=15.684 M=1 R=4.33333 SA=75004
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1018 A_951_47# N_A1_M1018_g N_A_79_204#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1019 A_1123_47# N_A1_M1019_g N_A_79_204#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=15.684 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_1123_47# VNB NSHORT L=0.15 W=0.65 AD=0.169
+ AS=0.091 PD=1.82 PS=0.93 NRD=0 NRS=15.684 M=1 R=4.33333 SA=75005.3 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_204#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1004_d N_A_79_204#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001
+ A=0.15 P=2.3 MULT=1
MM1012 N_VPWR_M1004_d N_A_79_204#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1015 N_VPWR_M1015_d N_A_79_204#_M1015_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1023 N_A_473_297#_M1023_d N_B1_M1023_g A_555_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=16.7253 M=1 R=6.66667 SA=75000.2
+ SB=75003.5 A=0.15 P=2.3 MULT=1
MM1008 A_555_297# N_C1_M1008_g N_A_79_204#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75003 A=0.15 P=2.3 MULT=1
MM1020 A_727_297# N_C1_M1020_g N_A_79_204#_M1008_s VPB PHIGHVT L=0.15 W=1
+ AD=0.16 AS=0.14 PD=1.32 PS=1.28 NRD=20.6653 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75002.6 A=0.15 P=2.3 MULT=1
MM1010 N_A_473_297#_M1010_d N_B1_M1010_g A_727_297# VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.16 PD=1.39 PS=1.32 NRD=7.8603 NRS=20.6653 M=1 R=6.66667
+ SA=75001.5 SB=75002.1 A=0.15 P=2.3 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_473_297#_M1010_d VPB PHIGHVT L=0.15 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=0 NRS=13.7703 M=1 R=6.66667 SA=75002.1
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1016 N_A_473_297#_M1016_d N_A1_M1016_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.195 PD=1.28 PS=1.39 NRD=0 NRS=21.67 M=1 R=6.66667 SA=75002.6
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1021 N_A_473_297#_M1016_d N_A1_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003 SB=75000.6
+ A=0.15 P=2.3 MULT=1
MM1009 N_VPWR_M1021_s N_A2_M1009_g N_A_473_297#_M1009_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.26 PD=1.28 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.5
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref VNB VPB NWDIODE A=10.9461 P=16.85
c_101 VPB 0 2.77707e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hd__a211o_4.spice.SKY130_FD_SC_HD__A211O_4.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__a311oi_2.spice.pex
* Created: Thu Aug 27 14:04:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__A311OI_2%A3 1 3 6 8 10 13 15 16 24
r36 22 24 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.89 $Y2=1.16
r37 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r38 19 22 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.47 $Y=1.16
+ $X2=0.595 $Y2=1.16
r39 16 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.595 $Y2=1.16
r40 15 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.235 $Y=1.16
+ $X2=0.595 $Y2=1.16
r41 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.16
r42 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.985
r43 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r44 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r45 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r46 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.985
r47 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A2 1 3 6 8 10 13 15 16 23 25
r46 24 25 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.73 $Y=1.16 $X2=1.74
+ $Y2=1.16
r47 22 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.71 $Y=1.16 $X2=1.73
+ $Y2=1.16
r48 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.16 $X2=1.71 $Y2=1.16
r49 19 22 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=1.31 $Y=1.16 $X2=1.71
+ $Y2=1.16
r50 16 23 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=1.71 $Y2=1.16
r51 15 16 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.155 $Y=1.16
+ $X2=1.615 $Y2=1.16
r52 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.325
+ $X2=1.74 $Y2=1.16
r53 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.74 $Y=1.325
+ $X2=1.74 $Y2=1.985
r54 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r55 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.325
+ $X2=1.31 $Y2=1.16
r57 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.31 $Y=1.325 $X2=1.31
+ $Y2=1.985
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A1 3 7 9 11 12 14 15 16 17 31
r48 29 31 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.92 $Y=1.16
+ $X2=3.09 $Y2=1.16
r49 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=1.16 $X2=2.92 $Y2=1.16
r50 27 29 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.67 $Y=1.16
+ $X2=2.92 $Y2=1.16
r51 26 27 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.6 $Y=1.16 $X2=2.67
+ $Y2=1.16
r52 24 26 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.24 $Y=1.16 $X2=2.6
+ $Y2=1.16
r53 24 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r54 21 24 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.18 $Y=1.16 $X2=2.24
+ $Y2=1.16
r55 17 30 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.015 $Y=1.16
+ $X2=2.92 $Y2=1.16
r56 16 30 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.555 $Y=1.16
+ $X2=2.92 $Y2=1.16
r57 16 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.555 $Y=1.16
+ $X2=2.24 $Y2=1.16
r58 15 25 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.095 $Y=1.16
+ $X2=2.24 $Y2=1.16
r59 12 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=1.16
r60 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.09 $Y=0.995
+ $X2=3.09 $Y2=0.56
r61 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=1.16
r62 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.67 $Y=0.995
+ $X2=2.67 $Y2=0.56
r63 5 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.325 $X2=2.6
+ $Y2=1.16
r64 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.6 $Y=1.325 $X2=2.6
+ $Y2=1.985
r65 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=1.325
+ $X2=2.18 $Y2=1.16
r66 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.18 $Y=1.325 $X2=2.18
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%B1 1 3 6 8 10 13 15 16 24
r50 22 24 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.89 $Y=1.16 $X2=3.96
+ $Y2=1.16
r51 19 22 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=3.54 $Y=1.16
+ $X2=3.89 $Y2=1.16
r52 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.89
+ $Y=1.16 $X2=3.89 $Y2=1.16
r53 15 16 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.495 $Y=1.16
+ $X2=3.89 $Y2=1.16
r54 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=1.325
+ $X2=3.96 $Y2=1.16
r55 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.96 $Y=1.325
+ $X2=3.96 $Y2=1.985
r56 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.96 $Y=0.995
+ $X2=3.96 $Y2=1.16
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.96 $Y=0.995
+ $X2=3.96 $Y2=0.56
r58 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.325
+ $X2=3.54 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.54 $Y=1.325 $X2=3.54
+ $Y2=1.985
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=0.995
+ $X2=3.54 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.54 $Y=0.995 $X2=3.54
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%C1 1 3 6 8 10 13 15 16 17 22 26 30
r47 22 24 29.7437 $w=3.16e-07 $l=1.95e-07 $layer=POLY_cond $X=5.05 $Y=1.16
+ $X2=5.245 $Y2=1.16
r48 21 22 64.0633 $w=3.16e-07 $l=4.2e-07 $layer=POLY_cond $X=4.63 $Y=1.16
+ $X2=5.05 $Y2=1.16
r49 17 30 11.5244 $w=2.33e-07 $l=2.35e-07 $layer=LI1_cond $X=5.292 $Y=1.53
+ $X2=5.292 $Y2=1.295
r50 16 30 3.30782 $w=2.35e-07 $l=1.1e-07 $layer=LI1_cond $X=5.292 $Y=1.185
+ $X2=5.292 $Y2=1.295
r51 16 26 3.51831 $w=2.2e-07 $l=1.17e-07 $layer=LI1_cond $X=5.292 $Y=1.185
+ $X2=5.175 $Y2=1.185
r52 16 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.245
+ $Y=1.16 $X2=5.245 $Y2=1.16
r53 15 26 18.3343 $w=2.18e-07 $l=3.5e-07 $layer=LI1_cond $X=4.825 $Y=1.185
+ $X2=5.175 $Y2=1.185
r54 11 22 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.16
r55 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.325
+ $X2=5.05 $Y2=1.985
r56 8 22 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=1.16
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.995
+ $X2=5.05 $Y2=0.56
r58 4 21 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=1.325
+ $X2=4.63 $Y2=1.16
r59 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.63 $Y=1.325 $X2=4.63
+ $Y2=1.985
r60 1 21 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=0.995
+ $X2=4.63 $Y2=1.16
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.63 $Y=0.995 $X2=4.63
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%VPWR 1 2 3 4 13 15 21 25 29 32 33 35 36 37
+ 39 55 56 62
r77 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 53 56 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 52 55 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 50 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r84 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r85 47 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r86 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.1 $Y2=2.72
r88 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=1.61 $Y2=2.72
r89 43 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r90 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 40 59 4.03846 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r92 40 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r93 39 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=1.1 $Y2=2.72
r94 39 42 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 37 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 35 49 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.53 $Y2=2.72
r98 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=2.72
+ $X2=2.81 $Y2=2.72
r99 34 52 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.975 $Y=2.72
+ $X2=2.99 $Y2=2.72
r100 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=2.72
+ $X2=2.81 $Y2=2.72
r101 32 46 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.61 $Y2=2.72
r102 32 33 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.785 $Y=2.72
+ $X2=1.96 $Y2=2.72
r103 31 49 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 31 33 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=1.96 $Y2=2.72
r105 27 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=2.635
+ $X2=2.81 $Y2=2.72
r106 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.81 $Y=2.635
+ $X2=2.81 $Y2=2
r107 23 33 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.635
+ $X2=1.96 $Y2=2.72
r108 23 25 20.9086 $w=3.48e-07 $l=6.35e-07 $layer=LI1_cond $X=1.96 $Y=2.635
+ $X2=1.96 $Y2=2
r109 19 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.635 $X2=1.1
+ $Y2=2.72
r110 19 21 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.1 $Y=2.635
+ $X2=1.1 $Y2=2
r111 15 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.22 $Y=1.66
+ $X2=0.22 $Y2=2.34
r112 13 59 3.10471 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.22 $Y=2.635
+ $X2=0.172 $Y2=2.72
r113 13 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.22 $Y=2.635
+ $X2=0.22 $Y2=2.34
r114 4 29 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.675
+ $Y=1.485 $X2=2.81 $Y2=2
r115 3 25 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.815
+ $Y=1.485 $X2=1.95 $Y2=2
r116 2 21 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.485 $X2=1.1 $Y2=2
r117 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r118 1 15 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A_109_297# 1 2 3 4 15 17 18 21 23 27 29 33
+ 34 36
r49 30 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=1.66
+ $X2=2.39 $Y2=1.66
r50 29 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=1.66
+ $X2=3.75 $Y2=1.66
r51 29 30 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.585 $Y=1.66
+ $X2=2.475 $Y2=1.66
r52 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=1.745
+ $X2=2.39 $Y2=1.66
r53 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.39 $Y=1.745
+ $X2=2.39 $Y2=1.96
r54 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.66
+ $X2=1.52 $Y2=1.66
r55 23 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=1.66
+ $X2=2.39 $Y2=1.66
r56 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.305 $Y=1.66
+ $X2=1.605 $Y2=1.66
r57 19 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=1.745
+ $X2=1.52 $Y2=1.66
r58 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.52 $Y=1.745
+ $X2=1.52 $Y2=1.96
r59 17 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=1.52 $Y2=1.66
r60 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=1.66
+ $X2=0.765 $Y2=1.66
r61 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.765 $Y2=1.66
r62 13 15 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.68 $Y=1.745
+ $X2=0.68 $Y2=1.96
r63 4 36 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.485 $X2=3.75 $Y2=1.66
r64 3 27 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.255
+ $Y=1.485 $X2=2.39 $Y2=1.96
r65 2 21 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=1.385
+ $Y=1.485 $X2=1.52 $Y2=1.96
r66 1 15 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A_641_297# 1 2 3 10 16 18 22 25
r36 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.26 $Y=2.255
+ $X2=5.26 $Y2=1.96
r37 19 25 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=4.44 $Y=2.34
+ $X2=4.275 $Y2=2.36
r38 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.175 $Y=2.34
+ $X2=5.26 $Y2=2.255
r39 18 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.175 $Y=2.34
+ $X2=4.44 $Y2=2.34
r40 14 25 0.89609 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.275 $Y=2.255
+ $X2=4.275 $Y2=2.36
r41 14 16 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.275 $Y=2.255
+ $X2=4.275 $Y2=2
r42 10 25 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=4.11 $Y=2.34
+ $X2=4.275 $Y2=2.36
r43 10 12 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.11 $Y=2.34
+ $X2=3.33 $Y2=2.34
r44 3 22 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=1.96
r45 2 25 600 $w=1.7e-07 $l=9.67587e-07 $layer=licon1_PDIFF $count=1 $X=4.035
+ $Y=1.485 $X2=4.275 $Y2=2.34
r46 2 16 600 $w=1.7e-07 $l=6.23558e-07 $layer=licon1_PDIFF $count=1 $X=4.035
+ $Y=1.485 $X2=4.275 $Y2=2
r47 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.485 $X2=3.33 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%Y 1 2 3 4 5 16 22 24 28 30 32 36 38 39 42
+ 43 44 45 54 56 61 64
r76 61 64 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.825 $Y=1.915
+ $X2=4.825 $Y2=1.87
r77 53 56 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=4.367 $Y=0.825
+ $X2=4.367 $Y2=0.85
r78 45 61 0.707246 $w=3.45e-07 $l=2e-08 $layer=LI1_cond $X=4.825 $Y=1.935
+ $X2=4.825 $Y2=1.915
r79 45 64 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=4.825 $Y=1.85
+ $X2=4.825 $Y2=1.87
r80 44 54 3.05574 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.367 $Y=1.595
+ $X2=4.367 $Y2=1.51
r81 44 54 1.76887 $w=2.13e-07 $l=3.3e-08 $layer=LI1_cond $X=4.367 $Y=1.477
+ $X2=4.367 $Y2=1.51
r82 43 44 15.3838 $w=2.13e-07 $l=2.87e-07 $layer=LI1_cond $X=4.367 $Y=1.19
+ $X2=4.367 $Y2=1.477
r83 42 53 0.130481 $w=1.68e-07 $l=2e-09 $layer=LI1_cond $X=4.365 $Y=0.74
+ $X2=4.367 $Y2=0.74
r84 42 65 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.365 $Y=0.74
+ $X2=4.17 $Y2=0.74
r85 42 43 16.6166 $w=2.13e-07 $l=3.1e-07 $layer=LI1_cond $X=4.367 $Y=0.88
+ $X2=4.367 $Y2=1.19
r86 42 56 1.60806 $w=2.13e-07 $l=3e-08 $layer=LI1_cond $X=4.367 $Y=0.88
+ $X2=4.367 $Y2=0.85
r87 39 45 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.825 $Y=1.745
+ $X2=4.825 $Y2=1.85
r88 39 41 2.95067 $w=3.3e-07 $l=1.2145e-07 $layer=LI1_cond $X=4.825 $Y=1.745
+ $X2=4.832 $Y2=1.627
r89 34 36 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.26 $Y=0.655
+ $X2=5.26 $Y2=0.42
r90 33 44 3.88258 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=4.475 $Y=1.595
+ $X2=4.367 $Y2=1.595
r91 32 41 4.8155 $w=1.7e-07 $l=1.87318e-07 $layer=LI1_cond $X=4.66 $Y=1.595
+ $X2=4.832 $Y2=1.627
r92 32 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.66 $Y=1.595
+ $X2=4.475 $Y2=1.595
r93 31 53 7.04599 $w=1.68e-07 $l=1.08e-07 $layer=LI1_cond $X=4.475 $Y=0.74
+ $X2=4.367 $Y2=0.74
r94 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.175 $Y=0.74
+ $X2=5.26 $Y2=0.655
r95 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.175 $Y=0.74
+ $X2=4.475 $Y2=0.74
r96 26 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.655
+ $X2=4.17 $Y2=0.74
r97 26 28 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.17 $Y=0.655
+ $X2=4.17 $Y2=0.42
r98 25 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=0.74
+ $X2=3.32 $Y2=0.74
r99 24 65 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.74
+ $X2=4.17 $Y2=0.74
r100 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.085 $Y=0.74
+ $X2=3.405 $Y2=0.74
r101 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=0.655
+ $X2=3.32 $Y2=0.74
r102 20 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.32 $Y=0.655
+ $X2=3.32 $Y2=0.42
r103 16 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=0.74
+ $X2=3.32 $Y2=0.74
r104 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.235 $Y=0.74
+ $X2=2.46 $Y2=0.74
r105 5 41 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=4.705
+ $Y=1.485 $X2=4.84 $Y2=1.66
r106 4 36 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.42
r107 3 28 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.035
+ $Y=0.235 $X2=4.17 $Y2=0.42
r108 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.235 $X2=3.32 $Y2=0.42
r109 1 18 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.46 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A_27_47# 1 2 3 12 14 15 18 22 24
r31 20 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.74 $X2=1.1
+ $Y2=0.74
r32 20 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=0.74
+ $X2=1.94 $Y2=0.74
r33 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.655 $X2=1.1
+ $Y2=0.74
r34 16 18 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.1 $Y=0.655
+ $X2=1.1 $Y2=0.42
r35 14 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.74 $X2=1.1
+ $Y2=0.74
r36 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.015 $Y=0.74
+ $X2=0.345 $Y2=0.74
r37 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.655
+ $X2=0.345 $Y2=0.74
r38 10 12 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.26 $Y=0.655
+ $X2=0.26 $Y2=0.42
r39 3 22 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.74
r40 2 18 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.42
r41 1 12 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%VGND 1 2 3 12 16 20 23 24 25 27 39 45 46 49
+ 52
r82 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r83 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r84 46 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r85 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r86 43 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=4.84
+ $Y2=0
r87 43 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.29
+ $Y2=0
r88 42 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r89 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r90 39 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.84
+ $Y2=0
r91 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.675 $Y=0 $X2=4.37
+ $Y2=0
r92 38 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r93 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r94 35 38 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r95 35 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r96 34 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r97 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r98 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r99 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.15
+ $Y2=0
r100 27 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r101 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r102 25 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r103 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r104 23 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.585 $Y=0
+ $X2=3.45 $Y2=0
r105 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.75
+ $Y2=0
r106 22 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.915 $Y=0
+ $X2=4.37 $Y2=0
r107 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.75
+ $Y2=0
r108 18 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0
r109 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0.38
r110 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0
r111 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0.38
r112 10 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r113 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r114 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.705
+ $Y=0.235 $X2=4.84 $Y2=0.38
r115 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.235 $X2=3.75 $Y2=0.38
r116 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__A311OI_2%A_277_47# 1 2 11
r18 8 11 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.52 $Y=0.39
+ $X2=2.88 $Y2=0.39
r19 2 11 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.745
+ $Y=0.235 $X2=2.88 $Y2=0.39
r20 1 8 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.39
.ends


* File: sky130_fd_sc_hd__or2b_2.spice.pex
* Created: Thu Aug 27 14:43:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__OR2B_2%B_N 3 7 9 15 18
r24 12 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.26 $Y=1.16
+ $X2=0.47 $Y2=1.16
r25 9 18 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r26 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r27 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=1.325
+ $X2=0.47 $Y2=1.16
r28 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.47 $Y=1.325 $X2=0.47
+ $Y2=1.695
r29 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r30 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%A_27_53# 1 2 9 13 17 19 20 23 27 37
r44 36 37 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.365 $Y=1.16
+ $X2=1.425 $Y2=1.16
r45 28 36 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.215 $Y=1.16
+ $X2=1.365 $Y2=1.16
r46 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r47 25 33 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.717 $Y=1.16
+ $X2=0.717 $Y2=1.325
r48 25 27 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.84 $Y=1.16
+ $X2=1.215 $Y2=1.16
r49 23 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.68 $Y=1.63
+ $X2=0.68 $Y2=1.325
r50 19 25 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.717 $Y=0.82
+ $X2=0.717 $Y2=1.16
r51 19 20 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.595 $Y=0.82
+ $X2=0.42 $Y2=0.82
r52 15 20 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=0.262 $Y=0.735
+ $X2=0.42 $Y2=0.82
r53 15 17 10.6098 $w=3.13e-07 $l=2.9e-07 $layer=LI1_cond $X=0.262 $Y=0.735
+ $X2=0.262 $Y2=0.445
r54 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.325
+ $X2=1.425 $Y2=1.16
r55 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.425 $Y=1.325
+ $X2=1.425 $Y2=1.695
r56 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=1.16
r57 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.365 $Y=0.995
+ $X2=1.365 $Y2=0.475
r58 2 23 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.63
r59 1 17 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%A 1 5 8 9 15
r36 12 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=2.28
+ $X2=1.17 $Y2=2.28
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.005
+ $Y=2.28 $X2=1.005 $Y2=2.28
r38 9 13 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.15 $Y=2.25
+ $X2=1.005 $Y2=2.25
r39 5 8 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=1.785 $Y=0.475
+ $X2=1.785 $Y2=1.695
r40 3 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.785 $Y=2.265
+ $X2=1.785 $Y2=1.695
r41 1 3 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.71 $Y=2.34
+ $X2=1.785 $Y2=2.265
r42 1 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.71 $Y=2.34 $X2=1.17
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%A_218_297# 1 2 7 9 12 14 16 19 21 25 27 28 32
+ 33 39 41 46
c76 32 0 1.06604e-19 $X=2.145 $Y=1.495
r77 45 46 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.275 $Y=1.16
+ $X2=2.695 $Y2=1.16
r78 40 45 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.205 $Y=1.16
+ $X2=2.275 $Y2=1.16
r79 39 42 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.16
+ $X2=2.175 $Y2=1.325
r80 39 41 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.16
+ $X2=2.175 $Y2=0.995
r81 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.205
+ $Y=1.16 $X2=2.205 $Y2=1.16
r82 33 36 2.88111 $w=4.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.195 $Y=1.58
+ $X2=1.195 $Y2=1.685
r83 32 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.145 $Y=1.495
+ $X2=2.145 $Y2=1.325
r84 29 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.145 $Y=0.825
+ $X2=2.145 $Y2=0.995
r85 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.74
+ $X2=2.145 $Y2=0.825
r86 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.06 $Y=0.74 $X2=1.66
+ $Y2=0.74
r87 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.575 $Y=0.655
+ $X2=1.66 $Y2=0.74
r88 23 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.575 $Y=0.655
+ $X2=1.575 $Y2=0.47
r89 22 33 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.405 $Y=1.58
+ $X2=1.195 $Y2=1.58
r90 21 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=1.58
+ $X2=2.145 $Y2=1.495
r91 21 22 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.06 $Y=1.58
+ $X2=1.405 $Y2=1.58
r92 17 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.325
+ $X2=2.695 $Y2=1.16
r93 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.695 $Y=1.325
+ $X2=2.695 $Y2=1.985
r94 14 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=0.995
+ $X2=2.695 $Y2=1.16
r95 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.695 $Y=0.995
+ $X2=2.695 $Y2=0.56
r96 10 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.325
+ $X2=2.275 $Y2=1.16
r97 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.275 $Y=1.325
+ $X2=2.275 $Y2=1.985
r98 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.995
+ $X2=2.275 $Y2=0.56
r100 2 36 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.485 $X2=1.215 $Y2=1.685
r101 1 25 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.265 $X2=1.575 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%VPWR 1 2 3 10 12 16 18 20 24 26 34 43 47
c39 2 0 1.06604e-19 $X=1.86 $Y=1.485
r40 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r43 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 35 43 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.19 $Y=2.72 $X2=2.05
+ $Y2=2.72
r46 35 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.19 $Y=2.72
+ $X2=2.53 $Y2=2.72
r47 34 46 3.98735 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=2.72 $X2=3.01
+ $Y2=2.72
r48 34 37 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.8 $Y=2.72 $X2=2.53
+ $Y2=2.72
r49 33 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r51 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 29 32 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 27 40 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r55 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 26 43 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=2.05
+ $Y2=2.72
r57 26 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.91 $Y=2.72 $X2=1.61
+ $Y2=2.72
r58 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r60 20 23 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=2.927 $Y=1.65
+ $X2=2.927 $Y2=2.33
r61 18 46 3.18988 $w=2.55e-07 $l=1.19499e-07 $layer=LI1_cond $X=2.927 $Y=2.635
+ $X2=3.01 $Y2=2.72
r62 18 23 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=2.927 $Y=2.635
+ $X2=2.927 $Y2=2.33
r63 14 43 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.635
+ $X2=2.05 $Y2=2.72
r64 14 16 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.05 $Y=2.635
+ $X2=2.05 $Y2=2
r65 10 40 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r66 10 12 43.2166 $w=2.58e-07 $l=9.75e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.66
r67 3 23 400 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=2.77 $Y=1.485
+ $X2=2.905 $Y2=2.33
r68 3 20 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.485 $X2=2.905 $Y2=1.65
r69 2 16 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.485 $X2=2.06 $Y2=2
r70 1 12 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%X 1 2 10 13 14 15
r24 13 15 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=2.515 $Y=1.61
+ $X2=2.515 $Y2=1.845
r25 13 14 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.515 $Y=1.61
+ $X2=2.515 $Y2=1.495
r26 12 14 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.545 $Y=0.76
+ $X2=2.545 $Y2=1.495
r27 10 12 9.32577 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.515 $Y=0.59
+ $X2=2.515 $Y2=0.76
r28 2 15 300 $w=1.7e-07 $l=4.22137e-07 $layer=licon1_PDIFF $count=2 $X=2.35
+ $Y=1.485 $X2=2.485 $Y2=1.845
r29 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.485 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HD__OR2B_2%VGND 1 2 3 12 14 16 18 25 30 38 44 46 50
r48 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r50 43 44 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=0.24
+ $X2=1.32 $Y2=0.24
r51 40 43 0.092006 $w=6.48e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=0.24
+ $X2=1.155 $Y2=0.24
r52 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 37 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r54 36 40 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r55 36 38 9.28585 $w=6.48e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=0.24 $X2=0.59
+ $Y2=0.24
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 34 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r58 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r59 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 31 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.02
+ $Y2=0
r61 31 33 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.53
+ $Y2=0
r62 30 49 3.98735 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.01
+ $Y2=0
r63 30 33 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.53
+ $Y2=0
r64 29 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r65 29 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r66 28 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.32
+ $Y2=0
r67 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r68 25 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=2.02
+ $Y2=0
r69 25 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.61
+ $Y2=0
r70 22 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.59
+ $Y2=0
r71 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r72 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r73 14 49 3.18988 $w=2.55e-07 $l=1.19499e-07 $layer=LI1_cond $X=2.927 $Y=0.085
+ $X2=3.01 $Y2=0
r74 14 16 13.5582 $w=2.53e-07 $l=3e-07 $layer=LI1_cond $X=2.927 $Y=0.085
+ $X2=2.927 $Y2=0.385
r75 10 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r76 10 12 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.4
r77 3 16 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=2.77
+ $Y=0.235 $X2=2.905 $Y2=0.385
r78 2 12 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.265 $X2=2.045 $Y2=0.4
r79 1 43 91 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.265 $X2=1.155 $Y2=0.4
.ends


* File: sky130_fd_sc_hd__nand2_8.pxi.spice
* Created: Thu Aug 27 14:28:57 2020
* 
x_PM_SKY130_FD_SC_HD__NAND2_8%B N_B_M1012_g N_B_M1001_g N_B_M1015_g N_B_M1004_g
+ N_B_M1016_g N_B_M1008_g N_B_M1018_g N_B_M1009_g N_B_M1020_g N_B_M1019_g
+ N_B_M1025_g N_B_M1022_g N_B_M1026_g N_B_M1027_g N_B_M1029_g N_B_M1028_g B B B
+ B B B N_B_c_179_p N_B_c_141_n PM_SKY130_FD_SC_HD__NAND2_8%B
x_PM_SKY130_FD_SC_HD__NAND2_8%A N_A_M1000_g N_A_M1002_g N_A_M1005_g N_A_M1003_g
+ N_A_M1007_g N_A_M1006_g N_A_M1021_g N_A_M1010_g N_A_M1023_g N_A_M1011_g
+ N_A_M1024_g N_A_M1013_g N_A_M1030_g N_A_M1014_g N_A_M1031_g N_A_M1017_g A A A
+ A A N_A_c_310_n PM_SKY130_FD_SC_HD__NAND2_8%A
x_PM_SKY130_FD_SC_HD__NAND2_8%VPWR N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1009_s
+ N_VPWR_M1022_s N_VPWR_M1028_s N_VPWR_M1003_d N_VPWR_M1010_d N_VPWR_M1013_d
+ N_VPWR_M1017_d N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n
+ N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n
+ N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n
+ N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n
+ VPWR N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_432_n
+ PM_SKY130_FD_SC_HD__NAND2_8%VPWR
x_PM_SKY130_FD_SC_HD__NAND2_8%Y N_Y_M1000_s N_Y_M1007_s N_Y_M1023_s N_Y_M1030_s
+ N_Y_M1001_d N_Y_M1008_d N_Y_M1019_d N_Y_M1027_d N_Y_M1002_s N_Y_M1006_s
+ N_Y_M1011_s N_Y_M1014_s N_Y_c_556_n N_Y_c_576_n N_Y_c_557_n N_Y_c_583_n
+ N_Y_c_558_n N_Y_c_591_n N_Y_c_559_n N_Y_c_599_n N_Y_c_560_n N_Y_c_620_n
+ N_Y_c_552_n N_Y_c_553_n N_Y_c_606_n N_Y_c_554_n N_Y_c_562_n N_Y_c_643_n
+ N_Y_c_563_n N_Y_c_651_n N_Y_c_564_n N_Y_c_659_n N_Y_c_662_n N_Y_c_555_n
+ N_Y_c_566_n N_Y_c_567_n N_Y_c_568_n N_Y_c_569_n N_Y_c_570_n N_Y_c_571_n Y Y
+ PM_SKY130_FD_SC_HD__NAND2_8%Y
x_PM_SKY130_FD_SC_HD__NAND2_8%A_27_47# N_A_27_47#_M1012_d N_A_27_47#_M1015_d
+ N_A_27_47#_M1018_d N_A_27_47#_M1025_d N_A_27_47#_M1029_d N_A_27_47#_M1005_d
+ N_A_27_47#_M1021_d N_A_27_47#_M1024_d N_A_27_47#_M1031_d N_A_27_47#_c_741_n
+ N_A_27_47#_c_742_n N_A_27_47#_c_743_n N_A_27_47#_c_760_n N_A_27_47#_c_744_n
+ N_A_27_47#_c_768_n N_A_27_47#_c_745_n N_A_27_47#_c_776_n N_A_27_47#_c_746_n
+ N_A_27_47#_c_784_n N_A_27_47#_c_747_n N_A_27_47#_c_799_n N_A_27_47#_c_748_n
+ N_A_27_47#_c_749_n N_A_27_47#_c_750_n N_A_27_47#_c_751_n N_A_27_47#_c_752_n
+ PM_SKY130_FD_SC_HD__NAND2_8%A_27_47#
x_PM_SKY130_FD_SC_HD__NAND2_8%VGND N_VGND_M1012_s N_VGND_M1016_s N_VGND_M1020_s
+ N_VGND_M1026_s N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n
+ N_VGND_c_874_n N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n
+ N_VGND_c_879_n N_VGND_c_880_n N_VGND_c_881_n VGND N_VGND_c_882_n
+ N_VGND_c_883_n PM_SKY130_FD_SC_HD__NAND2_8%VGND
cc_1 VNB N_B_M1012_g 0.0238771f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_B_M1001_g 7.2052e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_3 VNB N_B_M1015_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_4 VNB N_B_M1004_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_5 VNB N_B_M1016_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_6 VNB N_B_M1008_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_7 VNB N_B_M1018_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_8 VNB N_B_M1009_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_9 VNB N_B_M1020_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.56
cc_10 VNB N_B_M1019_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_11 VNB N_B_M1025_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.56
cc_12 VNB N_B_M1022_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.985
cc_13 VNB N_B_M1026_g 0.0173009f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.56
cc_14 VNB N_B_M1027_g 4.50027e-19 $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.985
cc_15 VNB N_B_M1029_g 0.0175542f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.56
cc_16 VNB N_B_M1028_g 4.63459e-19 $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_17 VNB N_B_c_141_n 0.138159f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.16
cc_18 VNB N_A_M1000_g 0.0171841f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB N_A_M1002_g 3.75525e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_20 VNB N_A_M1005_g 0.0172531f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_21 VNB N_A_M1003_g 4.47565e-19 $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_22 VNB N_A_M1007_g 0.0172831f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_23 VNB N_A_M1006_g 4.49831e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_24 VNB N_A_M1021_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_25 VNB N_A_M1010_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_26 VNB N_A_M1023_g 0.0173051f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.56
cc_27 VNB N_A_M1011_g 4.50211e-19 $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_28 VNB N_A_M1024_g 0.0172829f $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=0.56
cc_29 VNB N_A_M1013_g 4.49821e-19 $X=-0.19 $Y=-0.24 $X2=2.57 $Y2=1.985
cc_30 VNB N_A_M1030_g 0.0172529f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.56
cc_31 VNB N_A_M1014_g 4.47552e-19 $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.985
cc_32 VNB N_A_M1031_g 0.023255f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.56
cc_33 VNB N_A_M1017_g 6.82813e-19 $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_34 VNB N_A_c_310_n 0.138594f $X=-0.19 $Y=-0.24 $X2=3.2 $Y2=1.16
cc_35 VNB N_VPWR_c_432_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_552_n 0.0011304f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_37 VNB N_Y_c_553_n 0.00317716f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_38 VNB N_Y_c_554_n 0.0123853f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_39 VNB N_Y_c_555_n 0.00122694f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_741_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_41 VNB N_A_27_47#_c_742_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_743_n 0.013432f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.025
cc_43 VNB N_A_27_47#_c_744_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_44 VNB N_A_27_47#_c_745_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_c_746_n 0.00218355f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.56
cc_46 VNB N_A_27_47#_c_747_n 0.00317367f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.295
cc_47 VNB N_A_27_47#_c_748_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.985
cc_48 VNB N_A_27_47#_c_749_n 0.0234171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_27_47#_c_750_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.105
cc_50 VNB N_A_27_47#_c_751_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=1.53 $Y2=1.105
cc_51 VNB N_A_27_47#_c_752_n 0.00223024f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.105
cc_52 VNB N_VGND_c_870_n 0.00410835f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_53 VNB N_VGND_c_871_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_54 VNB N_VGND_c_872_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_55 VNB N_VGND_c_873_n 0.00410284f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_56 VNB N_VGND_c_874_n 0.0171909f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_57 VNB N_VGND_c_875_n 0.00323658f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.985
cc_58 VNB N_VGND_c_876_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.025
cc_59 VNB N_VGND_c_877_n 0.00323658f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=0.56
cc_60 VNB N_VGND_c_878_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_879_n 0.00323658f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.295
cc_62 VNB N_VGND_c_880_n 0.0166933f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.985
cc_63 VNB N_VGND_c_881_n 0.00323621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_882_n 0.0942509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_883_n 0.352291f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=1.295
cc_66 VPB N_B_M1001_g 0.0275655f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_67 VPB N_B_M1004_g 0.0193519f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_68 VPB N_B_M1008_g 0.0193519f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_69 VPB N_B_M1009_g 0.0193519f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_70 VPB N_B_M1019_g 0.0193519f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_71 VPB N_B_M1022_g 0.0193519f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_72 VPB N_B_M1027_g 0.0193486f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.985
cc_73 VPB N_B_M1028_g 0.0196272f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_74 VPB N_A_M1002_g 0.0180768f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_75 VPB N_A_M1003_g 0.0193049f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_76 VPB N_A_M1006_g 0.0193281f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_77 VPB N_A_M1010_g 0.0193519f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_78 VPB N_A_M1011_g 0.0193519f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.985
cc_79 VPB N_A_M1013_g 0.0193279f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_80 VPB N_A_M1014_g 0.0193046f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.985
cc_81 VPB N_A_M1017_g 0.0268823f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_82 VPB N_VPWR_c_433_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_434_n 0.0425966f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_84 VPB N_VPWR_c_435_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_436_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_437_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_438_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_439_n 0.00358901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_440_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.985
cc_90 VPB N_VPWR_c_441_n 0.00358901f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_91 VPB N_VPWR_c_442_n 0.00410835f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_92 VPB N_VPWR_c_443_n 0.0118743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_444_n 0.0452122f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.105
cc_94 VPB N_VPWR_c_445_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_446_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_447_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_448_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_449_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_99 VPB N_VPWR_c_450_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_451_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_101 VPB N_VPWR_c_452_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_102 VPB N_VPWR_c_453_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_103 VPB N_VPWR_c_454_n 0.00323736f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_104 VPB N_VPWR_c_455_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_105 VPB N_VPWR_c_456_n 0.00323736f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.16
cc_106 VPB N_VPWR_c_457_n 0.0185821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_458_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_432_n 0.0432074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_556_n 0.00224287f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.295
cc_110 VPB N_Y_c_557_n 0.00220047f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.025
cc_111 VPB N_Y_c_558_n 0.00220047f $X=-0.19 $Y=1.305 $X2=2.57 $Y2=1.985
cc_112 VPB N_Y_c_559_n 0.00220047f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.295
cc_113 VPB N_Y_c_560_n 0.00236841f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=0.56
cc_114 VPB N_Y_c_553_n 0.00412226f $X=-0.19 $Y=1.305 $X2=3.41 $Y2=1.985
cc_115 VPB N_Y_c_562_n 0.00228354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_Y_c_563_n 0.00228354f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.16
cc_117 VPB N_Y_c_564_n 0.00228354f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_118 VPB N_Y_c_555_n 0.00151227f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_566_n 0.00224287f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.185
cc_120 VPB N_Y_c_567_n 0.00224287f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.185
cc_121 VPB N_Y_c_568_n 0.00224287f $X=-0.19 $Y=1.305 $X2=2.075 $Y2=1.185
cc_122 VPB N_Y_c_569_n 0.00232853f $X=-0.19 $Y=1.305 $X2=2.995 $Y2=1.185
cc_123 VPB N_Y_c_570_n 0.00232853f $X=-0.19 $Y=1.305 $X2=3.2 $Y2=1.185
cc_124 VPB N_Y_c_571_n 6.7693e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 N_B_M1029_g N_A_M1000_g 0.0187087f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_126 N_B_M1028_g N_A_M1002_g 0.0187087f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_127 N_B_c_141_n N_A_c_310_n 0.0187087f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B_M1001_g N_VPWR_c_434_n 0.00321527f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B_M1004_g N_VPWR_c_435_n 0.00146448f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_130 N_B_M1008_g N_VPWR_c_435_n 0.00146448f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_131 N_B_M1009_g N_VPWR_c_436_n 0.00146448f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_132 N_B_M1019_g N_VPWR_c_436_n 0.00146448f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_133 N_B_M1022_g N_VPWR_c_437_n 0.00146448f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_134 N_B_M1027_g N_VPWR_c_437_n 0.00146448f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_135 N_B_M1028_g N_VPWR_c_438_n 0.00146448f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B_M1001_g N_VPWR_c_445_n 0.00541359f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B_M1004_g N_VPWR_c_445_n 0.00541359f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B_M1008_g N_VPWR_c_447_n 0.00541359f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_139 N_B_M1009_g N_VPWR_c_447_n 0.00541359f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_140 N_B_M1019_g N_VPWR_c_449_n 0.00541359f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_141 N_B_M1022_g N_VPWR_c_449_n 0.00541359f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_142 N_B_M1027_g N_VPWR_c_451_n 0.00541359f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_143 N_B_M1028_g N_VPWR_c_451_n 0.00541359f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_144 N_B_M1001_g N_VPWR_c_432_n 0.0104557f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_145 N_B_M1004_g N_VPWR_c_432_n 0.00950154f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_146 N_B_M1008_g N_VPWR_c_432_n 0.00950154f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_147 N_B_M1009_g N_VPWR_c_432_n 0.00950154f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_148 N_B_M1019_g N_VPWR_c_432_n 0.00950154f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_149 N_B_M1022_g N_VPWR_c_432_n 0.00950154f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_150 N_B_M1027_g N_VPWR_c_432_n 0.00950154f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_151 N_B_M1028_g N_VPWR_c_432_n 0.00952874f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_152 N_B_M1001_g N_Y_c_556_n 0.00395732f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_153 N_B_M1004_g N_Y_c_556_n 0.00120279f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_154 N_B_c_179_p N_Y_c_556_n 0.0268132f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B_c_141_n N_Y_c_556_n 0.00201507f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_156 N_B_M1001_g N_Y_c_576_n 0.00902485f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_157 N_B_M1004_g N_Y_c_576_n 0.00975139f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_158 N_B_M1008_g N_Y_c_576_n 6.1949e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_159 N_B_M1004_g N_Y_c_557_n 0.0115138f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_160 N_B_M1008_g N_Y_c_557_n 0.0115138f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_161 N_B_c_179_p N_Y_c_557_n 0.0366715f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B_c_141_n N_Y_c_557_n 0.00194394f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_163 N_B_M1004_g N_Y_c_583_n 6.1949e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_164 N_B_M1008_g N_Y_c_583_n 0.00975139f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_165 N_B_M1009_g N_Y_c_583_n 0.00975139f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_166 N_B_M1019_g N_Y_c_583_n 6.1949e-19 $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_167 N_B_M1009_g N_Y_c_558_n 0.0115138f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_168 N_B_M1019_g N_Y_c_558_n 0.0115138f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_169 N_B_c_179_p N_Y_c_558_n 0.0366715f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B_c_141_n N_Y_c_558_n 0.00194394f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B_M1009_g N_Y_c_591_n 6.1949e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_172 N_B_M1019_g N_Y_c_591_n 0.00975139f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_173 N_B_M1022_g N_Y_c_591_n 0.00975139f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_174 N_B_M1027_g N_Y_c_591_n 6.1949e-19 $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_175 N_B_M1022_g N_Y_c_559_n 0.0115138f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_176 N_B_M1027_g N_Y_c_559_n 0.0115138f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_177 N_B_c_179_p N_Y_c_559_n 0.0366715f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_178 N_B_c_141_n N_Y_c_559_n 0.00194394f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B_M1022_g N_Y_c_599_n 6.1949e-19 $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_180 N_B_M1027_g N_Y_c_599_n 0.00975139f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_181 N_B_M1028_g N_Y_c_599_n 0.00975139f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_182 N_B_M1028_g N_Y_c_560_n 0.0129763f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_183 N_B_M1029_g N_Y_c_552_n 8.79518e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_184 N_B_c_179_p N_Y_c_553_n 0.0131646f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_185 N_B_c_141_n N_Y_c_553_n 0.00643298f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_186 N_B_M1028_g N_Y_c_606_n 6.1949e-19 $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_187 N_B_M1008_g N_Y_c_566_n 0.00120279f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_188 N_B_M1009_g N_Y_c_566_n 0.00120279f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_189 N_B_c_179_p N_Y_c_566_n 0.0268132f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_190 N_B_c_141_n N_Y_c_566_n 0.00201507f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_191 N_B_M1019_g N_Y_c_567_n 0.00120279f $X=2.15 $Y=1.985 $X2=0 $Y2=0
cc_192 N_B_M1022_g N_Y_c_567_n 0.00120279f $X=2.57 $Y=1.985 $X2=0 $Y2=0
cc_193 N_B_c_179_p N_Y_c_567_n 0.0268132f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_194 N_B_c_141_n N_Y_c_567_n 0.00201507f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B_M1027_g N_Y_c_568_n 0.00120279f $X=2.99 $Y=1.985 $X2=0 $Y2=0
cc_196 N_B_M1028_g N_Y_c_568_n 0.00120279f $X=3.41 $Y=1.985 $X2=0 $Y2=0
cc_197 N_B_c_179_p N_Y_c_568_n 0.0268132f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_c_141_n N_Y_c_568_n 0.00201507f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B_M1012_g N_A_27_47#_c_741_n 0.00641402f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_200 N_B_M1015_g N_A_27_47#_c_741_n 5.25091e-19 $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_201 N_B_M1012_g N_A_27_47#_c_742_n 0.0110674f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_202 N_B_M1015_g N_A_27_47#_c_742_n 0.00850187f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_203 N_B_c_179_p N_A_27_47#_c_742_n 0.0303686f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B_c_141_n N_A_27_47#_c_742_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B_M1012_g N_A_27_47#_c_743_n 0.00234776f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_206 N_B_M1012_g N_A_27_47#_c_760_n 5.25176e-19 $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_207 N_B_M1015_g N_A_27_47#_c_760_n 0.00641402f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_208 N_B_M1016_g N_A_27_47#_c_760_n 0.00641402f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_209 N_B_M1018_g N_A_27_47#_c_760_n 5.25176e-19 $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_210 N_B_M1016_g N_A_27_47#_c_744_n 0.00850187f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_211 N_B_M1018_g N_A_27_47#_c_744_n 0.00850187f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_212 N_B_c_179_p N_A_27_47#_c_744_n 0.0362126f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B_c_141_n N_A_27_47#_c_744_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B_M1016_g N_A_27_47#_c_768_n 5.25176e-19 $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B_M1018_g N_A_27_47#_c_768_n 0.00641402f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B_M1020_g N_A_27_47#_c_768_n 0.00641402f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_217 N_B_M1025_g N_A_27_47#_c_768_n 5.25176e-19 $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B_M1020_g N_A_27_47#_c_745_n 0.00850187f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_219 N_B_M1025_g N_A_27_47#_c_745_n 0.00850187f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_220 N_B_c_179_p N_A_27_47#_c_745_n 0.0362126f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_221 N_B_c_141_n N_A_27_47#_c_745_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_M1020_g N_A_27_47#_c_776_n 5.25176e-19 $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_223 N_B_M1025_g N_A_27_47#_c_776_n 0.00641402f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B_M1026_g N_A_27_47#_c_776_n 0.00641402f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B_M1029_g N_A_27_47#_c_776_n 5.25176e-19 $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_226 N_B_M1026_g N_A_27_47#_c_746_n 0.00845772f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_227 N_B_M1029_g N_A_27_47#_c_746_n 0.00962612f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_228 N_B_c_179_p N_A_27_47#_c_746_n 0.0300229f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B_c_141_n N_A_27_47#_c_746_n 0.00205431f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B_M1029_g N_A_27_47#_c_784_n 0.00265763f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B_M1026_g N_A_27_47#_c_747_n 4.58193e-19 $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_232 N_B_M1029_g N_A_27_47#_c_747_n 0.00523631f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B_M1015_g N_A_27_47#_c_750_n 0.00110555f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_234 N_B_M1016_g N_A_27_47#_c_750_n 0.00110555f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_235 N_B_c_179_p N_A_27_47#_c_750_n 0.0267108f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B_c_141_n N_A_27_47#_c_750_n 0.00213429f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_237 N_B_M1018_g N_A_27_47#_c_751_n 0.00110555f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1020_g N_A_27_47#_c_751_n 0.00110555f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_c_179_p N_A_27_47#_c_751_n 0.0267108f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B_c_141_n N_A_27_47#_c_751_n 0.00213429f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_241 N_B_M1025_g N_A_27_47#_c_752_n 0.00110555f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1026_g N_A_27_47#_c_752_n 0.00110555f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_c_179_p N_A_27_47#_c_752_n 0.0267108f $X=3.2 $Y=1.16 $X2=0 $Y2=0
cc_244 N_B_c_141_n N_A_27_47#_c_752_n 0.00213429f $X=3.41 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B_M1012_g N_VGND_c_870_n 0.00268723f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B_M1015_g N_VGND_c_870_n 0.00146448f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_247 N_B_M1016_g N_VGND_c_871_n 0.00146448f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_248 N_B_M1018_g N_VGND_c_871_n 0.00146448f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B_M1020_g N_VGND_c_872_n 0.00146448f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B_M1025_g N_VGND_c_872_n 0.00146448f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B_M1026_g N_VGND_c_873_n 0.00146448f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_252 N_B_M1029_g N_VGND_c_873_n 0.00268723f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_253 N_B_M1012_g N_VGND_c_874_n 0.00424416f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_254 N_B_M1015_g N_VGND_c_876_n 0.00424416f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_255 N_B_M1016_g N_VGND_c_876_n 0.00424416f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_256 N_B_M1018_g N_VGND_c_878_n 0.00424416f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_257 N_B_M1020_g N_VGND_c_878_n 0.00424416f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_258 N_B_M1025_g N_VGND_c_880_n 0.00424416f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_259 N_B_M1026_g N_VGND_c_880_n 0.00424416f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_260 N_B_M1029_g N_VGND_c_882_n 0.00422898f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_261 N_B_M1012_g N_VGND_c_883_n 0.00669028f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_262 N_B_M1015_g N_VGND_c_883_n 0.00573607f $X=0.89 $Y=0.56 $X2=0 $Y2=0
cc_263 N_B_M1016_g N_VGND_c_883_n 0.00573607f $X=1.31 $Y=0.56 $X2=0 $Y2=0
cc_264 N_B_M1018_g N_VGND_c_883_n 0.00573607f $X=1.73 $Y=0.56 $X2=0 $Y2=0
cc_265 N_B_M1020_g N_VGND_c_883_n 0.00573607f $X=2.15 $Y=0.56 $X2=0 $Y2=0
cc_266 N_B_M1025_g N_VGND_c_883_n 0.00573607f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_267 N_B_M1026_g N_VGND_c_883_n 0.00573607f $X=2.99 $Y=0.56 $X2=0 $Y2=0
cc_268 N_B_M1029_g N_VGND_c_883_n 0.00577235f $X=3.41 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A_M1002_g N_VPWR_c_438_n 0.00146448f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_270 N_A_M1003_g N_VPWR_c_439_n 0.00146448f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_271 N_A_M1006_g N_VPWR_c_439_n 0.00146448f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_M1006_g N_VPWR_c_440_n 0.00541359f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_273 N_A_M1010_g N_VPWR_c_440_n 0.00541359f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_M1010_g N_VPWR_c_441_n 0.00146448f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A_M1011_g N_VPWR_c_441_n 0.00146448f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_276 N_A_M1013_g N_VPWR_c_442_n 0.00146448f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_M1014_g N_VPWR_c_442_n 0.00268723f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_278 N_A_M1017_g N_VPWR_c_444_n 0.0268969f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_279 N_A_M1002_g N_VPWR_c_453_n 0.00541359f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_280 N_A_M1003_g N_VPWR_c_453_n 0.00541359f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_M1011_g N_VPWR_c_455_n 0.00541359f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_282 N_A_M1013_g N_VPWR_c_455_n 0.00541359f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_283 N_A_M1014_g N_VPWR_c_457_n 0.00541359f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_284 N_A_M1017_g N_VPWR_c_457_n 0.00541359f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_285 N_A_M1002_g N_VPWR_c_432_n 0.00952874f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_286 N_A_M1003_g N_VPWR_c_432_n 0.00950154f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_287 N_A_M1006_g N_VPWR_c_432_n 0.00950154f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_288 N_A_M1010_g N_VPWR_c_432_n 0.00950154f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_289 N_A_M1011_g N_VPWR_c_432_n 0.00950154f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_290 N_A_M1013_g N_VPWR_c_432_n 0.00950154f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_291 N_A_M1014_g N_VPWR_c_432_n 0.00950154f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_292 N_A_M1017_g N_VPWR_c_432_n 0.0107188f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_293 N_A_M1002_g N_Y_c_599_n 6.1949e-19 $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_294 N_A_M1000_g N_Y_c_620_n 0.00325271f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A_M1000_g N_Y_c_552_n 0.00314663f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A_M1005_g N_Y_c_552_n 0.00302963f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A_c_310_n N_Y_c_552_n 0.00603353f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_M1002_g N_Y_c_553_n 0.0163272f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_299 N_A_M1003_g N_Y_c_553_n 0.00647727f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_300 A N_Y_c_553_n 0.0163282f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_301 N_A_c_310_n N_Y_c_553_n 0.0184365f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_M1002_g N_Y_c_606_n 0.00975139f $X=3.83 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A_M1003_g N_Y_c_606_n 0.00975139f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_304 N_A_M1006_g N_Y_c_606_n 6.1949e-19 $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_305 N_A_M1005_g N_Y_c_554_n 0.0120487f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_M1007_g N_Y_c_554_n 0.0107009f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_M1021_g N_Y_c_554_n 0.0107009f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A_M1023_g N_Y_c_554_n 0.0107009f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_M1024_g N_Y_c_554_n 0.0107009f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A_M1030_g N_Y_c_554_n 0.0121073f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_311 A N_Y_c_554_n 0.147814f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A_c_310_n N_Y_c_554_n 0.010373f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_M1003_g N_Y_c_562_n 0.0125389f $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_314 N_A_M1006_g N_Y_c_562_n 0.0116113f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_315 A N_Y_c_562_n 0.0280381f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_316 N_A_c_310_n N_Y_c_562_n 0.00196602f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_M1003_g N_Y_c_643_n 6.1949e-19 $X=4.25 $Y=1.985 $X2=0 $Y2=0
cc_318 N_A_M1006_g N_Y_c_643_n 0.00975139f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_319 N_A_M1010_g N_Y_c_643_n 0.00975139f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_M1011_g N_Y_c_643_n 6.1949e-19 $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_321 N_A_M1010_g N_Y_c_563_n 0.0116113f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_322 N_A_M1011_g N_Y_c_563_n 0.0116113f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_323 A N_Y_c_563_n 0.0334099f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_324 N_A_c_310_n N_Y_c_563_n 0.00196602f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_M1010_g N_Y_c_651_n 6.1949e-19 $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_M1011_g N_Y_c_651_n 0.00975139f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_327 N_A_M1013_g N_Y_c_651_n 0.00975139f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_328 N_A_M1014_g N_Y_c_651_n 6.1949e-19 $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_M1013_g N_Y_c_564_n 0.0116113f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_330 N_A_M1014_g N_Y_c_564_n 0.0125941f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_331 A N_Y_c_564_n 0.0277202f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_332 N_A_c_310_n N_Y_c_564_n 0.00196602f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_M1013_g N_Y_c_659_n 6.1949e-19 $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_334 N_A_M1014_g N_Y_c_659_n 0.00975139f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_335 N_A_M1017_g N_Y_c_659_n 0.00943894f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_336 N_A_M1031_g N_Y_c_662_n 0.00339728f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_337 N_A_M1030_g N_Y_c_555_n 0.00306065f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_338 N_A_M1014_g N_Y_c_555_n 0.00434664f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_339 N_A_M1031_g N_Y_c_555_n 0.00604668f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A_M1017_g N_Y_c_555_n 0.00860884f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_341 A N_Y_c_555_n 0.0154944f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_342 N_A_c_310_n N_Y_c_555_n 0.0272316f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_343 N_A_M1006_g N_Y_c_569_n 0.0012288f $X=4.67 $Y=1.985 $X2=0 $Y2=0
cc_344 N_A_M1010_g N_Y_c_569_n 0.0012288f $X=5.09 $Y=1.985 $X2=0 $Y2=0
cc_345 A N_Y_c_569_n 0.0244853f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_346 N_A_c_310_n N_Y_c_569_n 0.0020448f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_M1011_g N_Y_c_570_n 0.0012288f $X=5.51 $Y=1.985 $X2=0 $Y2=0
cc_348 N_A_M1013_g N_Y_c_570_n 0.0012288f $X=5.93 $Y=1.985 $X2=0 $Y2=0
cc_349 A N_Y_c_570_n 0.0244853f $X=6.13 $Y=1.105 $X2=0 $Y2=0
cc_350 N_A_c_310_n N_Y_c_570_n 0.0020448f $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_351 N_A_M1014_g N_Y_c_571_n 0.00153652f $X=6.35 $Y=1.985 $X2=0 $Y2=0
cc_352 N_A_M1017_g N_Y_c_571_n 0.0036105f $X=6.77 $Y=1.985 $X2=0 $Y2=0
cc_353 N_A_M1000_g N_A_27_47#_c_799_n 0.0107976f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A_M1005_g N_A_27_47#_c_799_n 0.00918728f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_M1007_g N_A_27_47#_c_799_n 0.00918728f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_M1021_g N_A_27_47#_c_799_n 0.00918728f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_M1023_g N_A_27_47#_c_799_n 0.00918728f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_M1024_g N_A_27_47#_c_799_n 0.00918728f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_M1030_g N_A_27_47#_c_799_n 0.00918728f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_M1031_g N_A_27_47#_c_799_n 0.0180277f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_c_310_n N_A_27_47#_c_799_n 5.98765e-19 $X=6.77 $Y=1.16 $X2=0 $Y2=0
cc_362 N_A_M1031_g N_A_27_47#_c_749_n 0.00815319f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_M1000_g N_VGND_c_882_n 0.00357877f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_M1005_g N_VGND_c_882_n 0.00357877f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_365 N_A_M1007_g N_VGND_c_882_n 0.00357877f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_366 N_A_M1021_g N_VGND_c_882_n 0.00357877f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_M1023_g N_VGND_c_882_n 0.00357877f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_M1024_g N_VGND_c_882_n 0.00357877f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_369 N_A_M1030_g N_VGND_c_882_n 0.00357877f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_370 N_A_M1031_g N_VGND_c_882_n 0.00357877f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_M1000_g N_VGND_c_883_n 0.00525237f $X=3.83 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_M1005_g N_VGND_c_883_n 0.00522516f $X=4.25 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A_M1007_g N_VGND_c_883_n 0.00522516f $X=4.67 $Y=0.56 $X2=0 $Y2=0
cc_374 N_A_M1021_g N_VGND_c_883_n 0.00522516f $X=5.09 $Y=0.56 $X2=0 $Y2=0
cc_375 N_A_M1023_g N_VGND_c_883_n 0.00522516f $X=5.51 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A_M1024_g N_VGND_c_883_n 0.00522516f $X=5.93 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_M1030_g N_VGND_c_883_n 0.00522516f $X=6.35 $Y=0.56 $X2=0 $Y2=0
cc_378 N_A_M1031_g N_VGND_c_883_n 0.00635551f $X=6.77 $Y=0.56 $X2=0 $Y2=0
cc_379 N_VPWR_c_432_n N_Y_M1001_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_432_n N_Y_M1008_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_432_n N_Y_M1019_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_432_n N_Y_M1027_d 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_432_n N_Y_M1002_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_432_n N_Y_M1006_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_432_n N_Y_M1011_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_c_432_n N_Y_M1014_s 0.00215201f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_445_n N_Y_c_576_n 0.0189039f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_432_n N_Y_c_576_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_389 N_VPWR_M1004_s N_Y_c_557_n 0.00166664f $X=0.965 $Y=1.485 $X2=0 $Y2=0
cc_390 N_VPWR_c_435_n N_Y_c_557_n 0.0128323f $X=1.1 $Y=2 $X2=0 $Y2=0
cc_391 N_VPWR_c_447_n N_Y_c_583_n 0.0189039f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_432_n N_Y_c_583_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_M1009_s N_Y_c_558_n 0.00166664f $X=1.805 $Y=1.485 $X2=0 $Y2=0
cc_394 N_VPWR_c_436_n N_Y_c_558_n 0.0128323f $X=1.94 $Y=2 $X2=0 $Y2=0
cc_395 N_VPWR_c_449_n N_Y_c_591_n 0.0189039f $X=2.695 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_432_n N_Y_c_591_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_M1022_s N_Y_c_559_n 0.00166664f $X=2.645 $Y=1.485 $X2=0 $Y2=0
cc_398 N_VPWR_c_437_n N_Y_c_559_n 0.0128323f $X=2.78 $Y=2 $X2=0 $Y2=0
cc_399 N_VPWR_c_451_n N_Y_c_599_n 0.0189039f $X=3.535 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_432_n N_Y_c_599_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_M1028_s N_Y_c_560_n 0.00103631f $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_402 N_VPWR_c_438_n N_Y_c_560_n 0.00802394f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_M1028_s N_Y_c_553_n 6.39069e-19 $X=3.485 $Y=1.485 $X2=0 $Y2=0
cc_404 N_VPWR_c_438_n N_Y_c_553_n 0.0051749f $X=3.62 $Y=2 $X2=0 $Y2=0
cc_405 N_VPWR_c_453_n N_Y_c_606_n 0.0189039f $X=4.375 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_c_432_n N_Y_c_606_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_407 N_VPWR_M1003_d N_Y_c_562_n 0.00166664f $X=4.325 $Y=1.485 $X2=0 $Y2=0
cc_408 N_VPWR_c_439_n N_Y_c_562_n 0.0128323f $X=4.46 $Y=2 $X2=0 $Y2=0
cc_409 N_VPWR_c_440_n N_Y_c_643_n 0.0189039f $X=5.215 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_432_n N_Y_c_643_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_M1010_d N_Y_c_563_n 0.00166664f $X=5.165 $Y=1.485 $X2=0 $Y2=0
cc_412 N_VPWR_c_441_n N_Y_c_563_n 0.0128323f $X=5.3 $Y=2 $X2=0 $Y2=0
cc_413 N_VPWR_c_455_n N_Y_c_651_n 0.0189039f $X=6.055 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_432_n N_Y_c_651_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_M1013_d N_Y_c_564_n 0.00166664f $X=6.005 $Y=1.485 $X2=0 $Y2=0
cc_416 N_VPWR_c_442_n N_Y_c_564_n 0.0128323f $X=6.14 $Y=2 $X2=0 $Y2=0
cc_417 N_VPWR_c_444_n N_Y_c_659_n 0.0572868f $X=7.08 $Y=1.66 $X2=0 $Y2=0
cc_418 N_VPWR_c_457_n N_Y_c_659_n 0.0189039f $X=6.915 $Y=2.72 $X2=0 $Y2=0
cc_419 N_VPWR_c_432_n N_Y_c_659_n 0.0122217f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_444_n N_Y_c_571_n 0.0129178f $X=7.08 $Y=1.66 $X2=0 $Y2=0
cc_421 N_VPWR_c_434_n N_A_27_47#_c_743_n 0.00938479f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_422 N_VPWR_c_444_n N_A_27_47#_c_749_n 0.0132088f $X=7.08 $Y=1.66 $X2=0 $Y2=0
cc_423 N_Y_c_554_n N_A_27_47#_M1005_d 0.00162409f $X=6.475 $Y=0.78 $X2=0 $Y2=0
cc_424 N_Y_c_554_n N_A_27_47#_M1021_d 0.00162409f $X=6.475 $Y=0.78 $X2=0 $Y2=0
cc_425 N_Y_c_554_n N_A_27_47#_M1024_d 0.00162409f $X=6.475 $Y=0.78 $X2=0 $Y2=0
cc_426 N_Y_c_560_n N_A_27_47#_c_746_n 0.00229229f $X=3.64 $Y=1.565 $X2=0 $Y2=0
cc_427 N_Y_c_560_n N_A_27_47#_c_747_n 0.00659652f $X=3.64 $Y=1.565 $X2=0 $Y2=0
cc_428 N_Y_c_620_n N_A_27_47#_c_747_n 0.00808483f $X=3.997 $Y=0.905 $X2=0 $Y2=0
cc_429 N_Y_c_553_n N_A_27_47#_c_747_n 0.00600544f $X=4.04 $Y=1.665 $X2=0 $Y2=0
cc_430 N_Y_M1000_s N_A_27_47#_c_799_n 0.00305588f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_431 N_Y_M1007_s N_A_27_47#_c_799_n 0.0030596f $X=4.745 $Y=0.235 $X2=0 $Y2=0
cc_432 N_Y_M1023_s N_A_27_47#_c_799_n 0.0030596f $X=5.585 $Y=0.235 $X2=0 $Y2=0
cc_433 N_Y_M1030_s N_A_27_47#_c_799_n 0.00305588f $X=6.425 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Y_c_620_n N_A_27_47#_c_799_n 0.014471f $X=3.997 $Y=0.905 $X2=0 $Y2=0
cc_435 N_Y_c_553_n N_A_27_47#_c_799_n 0.00423797f $X=4.04 $Y=1.665 $X2=0 $Y2=0
cc_436 N_Y_c_554_n N_A_27_47#_c_799_n 0.117609f $X=6.475 $Y=0.78 $X2=0 $Y2=0
cc_437 N_Y_c_662_n N_A_27_47#_c_799_n 0.014471f $X=6.6 $Y=0.905 $X2=0 $Y2=0
cc_438 N_Y_c_662_n N_A_27_47#_c_749_n 0.0113403f $X=6.6 $Y=0.905 $X2=0 $Y2=0
cc_439 N_Y_M1000_s N_VGND_c_883_n 0.00216833f $X=3.905 $Y=0.235 $X2=0 $Y2=0
cc_440 N_Y_M1007_s N_VGND_c_883_n 0.00216833f $X=4.745 $Y=0.235 $X2=0 $Y2=0
cc_441 N_Y_M1023_s N_VGND_c_883_n 0.00216833f $X=5.585 $Y=0.235 $X2=0 $Y2=0
cc_442 N_Y_M1030_s N_VGND_c_883_n 0.00216833f $X=6.425 $Y=0.235 $X2=0 $Y2=0
cc_443 N_A_27_47#_c_742_n N_VGND_M1012_s 0.00162006f $X=0.935 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_444 N_A_27_47#_c_744_n N_VGND_M1016_s 0.00162006f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_c_745_n N_VGND_M1020_s 0.00162006f $X=2.615 $Y=0.82 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_746_n N_VGND_M1026_s 0.00162006f $X=3.455 $Y=0.82 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_742_n N_VGND_c_870_n 0.0122414f $X=0.935 $Y=0.82 $X2=0 $Y2=0
cc_448 N_A_27_47#_c_744_n N_VGND_c_871_n 0.0122414f $X=1.775 $Y=0.82 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_745_n N_VGND_c_872_n 0.0122414f $X=2.615 $Y=0.82 $X2=0 $Y2=0
cc_450 N_A_27_47#_c_746_n N_VGND_c_873_n 0.0122414f $X=3.455 $Y=0.82 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_741_n N_VGND_c_874_n 0.0213324f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_742_n N_VGND_c_874_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_453 N_A_27_47#_c_742_n N_VGND_c_876_n 0.00193763f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_c_760_n N_VGND_c_876_n 0.0188551f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_455 N_A_27_47#_c_744_n N_VGND_c_876_n 0.00193763f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_c_744_n N_VGND_c_878_n 0.00193763f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_768_n N_VGND_c_878_n 0.0188551f $X=1.94 $Y=0.4 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_745_n N_VGND_c_878_n 0.00193763f $X=2.615 $Y=0.82 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_745_n N_VGND_c_880_n 0.00193763f $X=2.615 $Y=0.82 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_776_n N_VGND_c_880_n 0.0188551f $X=2.78 $Y=0.4 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_746_n N_VGND_c_880_n 0.00193763f $X=3.455 $Y=0.82 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_746_n N_VGND_c_882_n 0.00193763f $X=3.455 $Y=0.82 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_784_n N_VGND_c_882_n 0.0152108f $X=3.58 $Y=0.485 $X2=0 $Y2=0
cc_464 N_A_27_47#_c_799_n N_VGND_c_882_n 0.177444f $X=6.895 $Y=0.37 $X2=0 $Y2=0
cc_465 N_A_27_47#_c_748_n N_VGND_c_882_n 0.0261024f $X=7.082 $Y=0.485 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1012_d N_VGND_c_883_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_M1015_d N_VGND_c_883_n 0.00215201f $X=0.965 $Y=0.235 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_M1018_d N_VGND_c_883_n 0.00215201f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_M1025_d N_VGND_c_883_n 0.00215201f $X=2.645 $Y=0.235 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_M1029_d N_VGND_c_883_n 0.00215206f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_M1005_d N_VGND_c_883_n 0.00215227f $X=4.325 $Y=0.235 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_M1021_d N_VGND_c_883_n 0.00215227f $X=5.165 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_M1024_d N_VGND_c_883_n 0.00215227f $X=6.005 $Y=0.235 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_M1031_d N_VGND_c_883_n 0.00308503f $X=6.845 $Y=0.235 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_741_n N_VGND_c_883_n 0.0126042f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_742_n N_VGND_c_883_n 0.00825759f $X=0.935 $Y=0.82 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_760_n N_VGND_c_883_n 0.0122069f $X=1.1 $Y=0.4 $X2=0 $Y2=0
cc_478 N_A_27_47#_c_744_n N_VGND_c_883_n 0.00825759f $X=1.775 $Y=0.82 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_768_n N_VGND_c_883_n 0.0122069f $X=1.94 $Y=0.4 $X2=0 $Y2=0
cc_480 N_A_27_47#_c_745_n N_VGND_c_883_n 0.00825759f $X=2.615 $Y=0.82 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_776_n N_VGND_c_883_n 0.0122069f $X=2.78 $Y=0.4 $X2=0 $Y2=0
cc_482 N_A_27_47#_c_746_n N_VGND_c_883_n 0.00825759f $X=3.455 $Y=0.82 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_784_n N_VGND_c_883_n 0.00940698f $X=3.58 $Y=0.485 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_c_799_n N_VGND_c_883_n 0.113624f $X=6.895 $Y=0.37 $X2=0 $Y2=0
cc_485 N_A_27_47#_c_748_n N_VGND_c_883_n 0.0144249f $X=7.082 $Y=0.485 $X2=0
+ $Y2=0

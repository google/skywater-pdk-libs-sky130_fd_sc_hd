* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__lpflow_decapkapwr_6 KAPWR VGND VNB VPB VPWR
M1000 KAPWR VGND KAPWR VPB phighvt w=870000u l=1.97e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND KAPWR VGND VNB nshort w=550000u l=1.97e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_hd__dlxtn_1.pex.spice
* Created: Tue Sep  1 19:06:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLXTN_1%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%A_27_47# 1 2 9 13 15 17 19 21 25 29 30 31 35
+ 41 44 46 52 56 57 60 63 64 68
c168 52 0 8.44901e-20 $X=3.2 $Y=1.745
c169 15 0 2.5173e-20 $X=2.725 $Y=0.73
c170 13 0 2.6965e-20 $X=0.89 $Y=2.135
c171 9 0 2.6965e-20 $X=0.89 $Y=0.445
r172 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.035 $Y=1.53
+ $X2=3.035 $Y2=1.53
r173 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r175 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.89 $Y=1.53
+ $X2=3.035 $Y2=1.53
r176 56 57 2.53712 $w=1.4e-07 $l=2.05e-06 $layer=MET1_cond $X=2.89 $Y=1.53
+ $X2=0.84 $Y2=1.53
r177 54 64 1.09756 $w=3.13e-07 $l=3e-08 $layer=LI1_cond $X=3.107 $Y=1.56
+ $X2=3.107 $Y2=1.53
r178 52 54 6.41959 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=3.117 $Y=1.745
+ $X2=3.117 $Y2=1.56
r179 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.745 $X2=3.2 $Y2=1.745
r180 49 64 17.9269 $w=3.13e-07 $l=4.9e-07 $layer=LI1_cond $X=3.107 $Y=1.04
+ $X2=3.107 $Y2=1.53
r181 48 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r182 47 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r183 45 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r184 44 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r185 44 46 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r186 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r187 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.745
+ $Y=0.91 $X2=2.745 $Y2=0.91
r188 35 49 6.8188 $w=3.05e-07 $l=2.20613e-07 $layer=LI1_cond $X=2.95 $Y=0.887
+ $X2=3.107 $Y2=1.04
r189 35 37 7.74593 $w=3.03e-07 $l=2.05e-07 $layer=LI1_cond $X=2.95 $Y=0.887
+ $X2=2.745 $Y2=0.887
r190 33 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r191 32 41 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r192 31 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r193 31 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r194 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r195 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r196 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r197 23 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r198 19 53 34.1986 $w=3.29e-07 $l=1.60156e-07 $layer=POLY_cond $X=3.145 $Y=1.88
+ $X2=3.2 $Y2=1.745
r199 19 21 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.145 $Y=1.88
+ $X2=3.145 $Y2=2.275
r200 15 38 40.7947 $w=3.35e-07 $l=1.84932e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.735 $Y2=0.91
r201 15 17 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=2.725 $Y=0.73
+ $X2=2.725 $Y2=0.415
r202 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r203 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r204 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r206 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%D 2 3 5 6 8 10 13 16 18 21 22
c57 16 0 5.59029e-20 $X=1.83 $Y=1.695
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.04 $X2=1.6 $Y2=1.04
r59 18 22 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.6 $Y=1.19 $X2=1.6
+ $Y2=1.04
r60 14 16 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.66 $Y=1.695
+ $X2=1.83 $Y2=1.695
r61 12 21 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=1.6 $Y=1.07 $X2=1.6
+ $Y2=1.04
r62 12 13 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=1.6 $Y=1.07 $X2=1.6
+ $Y2=1.205
r63 10 21 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.6 $Y=0.88 $X2=1.6
+ $Y2=1.04
r64 6 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=1.77 $X2=1.83
+ $Y2=1.695
r65 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.83 $Y=1.77 $X2=1.83
+ $Y2=2.165
r66 3 10 106.596 $w=1.04e-07 $l=2.3e-07 $layer=POLY_cond $X=1.83 $Y=0.805
+ $X2=1.6 $Y2=0.805
r67 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.83 $Y=0.73 $X2=1.83
+ $Y2=0.445
r68 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.66 $Y=1.62 $X2=1.66
+ $Y2=1.695
r69 2 13 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.66 $Y=1.62
+ $X2=1.66 $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%A_299_47# 1 2 9 11 13 17 19 22 24 27 30 35
c94 35 0 4.8632e-21 $X=2.215 $Y=1.07
c95 19 0 2.5173e-20 $X=1.945 $Y=0.7
r96 35 37 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.132 $Y=1.07
+ $X2=2.132 $Y2=1.235
r97 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.215
+ $Y=1.07 $X2=2.215 $Y2=1.07
r98 30 32 10.8065 $w=1.93e-07 $l=1.9e-07 $layer=LI1_cond $X=1.607 $Y=0.51
+ $X2=1.607 $Y2=0.7
r99 24 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.58
r100 24 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.235
r101 22 35 0.6761 $w=3.73e-07 $l=2.2e-08 $layer=LI1_cond $X=2.132 $Y=1.048
+ $X2=2.132 $Y2=1.07
r102 21 22 8.08247 $w=3.73e-07 $l=2.63e-07 $layer=LI1_cond $X=2.132 $Y=0.785
+ $X2=2.132 $Y2=1.048
r103 20 32 1.54022 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.607 $Y2=0.7
r104 19 21 34.7438 $w=6.3e-08 $l=2.2553e-07 $layer=LI1_cond $X=1.945 $Y=0.7
+ $X2=2.132 $Y2=0.785
r105 19 20 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.945 $Y=0.7
+ $X2=1.705 $Y2=0.7
r106 15 27 27.5968 $w=1.68e-07 $l=4.23e-07 $layer=LI1_cond $X=1.607 $Y=1.58
+ $X2=2.03 $Y2=1.58
r107 15 17 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=1.607 $Y=1.665
+ $X2=1.607 $Y2=1.99
r108 11 36 38.9235 $w=2.69e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.25 $Y=1.235
+ $X2=2.215 $Y2=1.07
r109 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.25 $Y=1.235
+ $X2=2.25 $Y2=2.165
r110 7 36 38.9235 $w=2.69e-07 $l=1.81659e-07 $layer=POLY_cond $X=2.25 $Y=0.905
+ $X2=2.215 $Y2=1.07
r111 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.25 $Y=0.905
+ $X2=2.25 $Y2=0.445
r112 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r113 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%A_193_47# 1 2 9 11 13 15 18 20 22 23 26 29
+ 34 35
c109 35 0 1.84897e-19 $X=2.725 $Y=1.42
c110 18 0 5.59029e-20 $X=1.1 $Y=0.51
r111 33 35 6.29478 $w=2.68e-07 $l=3.5e-08 $layer=POLY_cond $X=2.69 $Y=1.42
+ $X2=2.725 $Y2=1.42
r112 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.52 $X2=2.69 $Y2=1.52
r113 30 34 12.0404 $w=3.33e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r114 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=1.87
+ $X2=2.53 $Y2=1.87
r115 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r116 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r117 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=2.53 $Y2=1.87
r118 22 23 1.34282 $w=1.4e-07 $l=1.085e-06 $layer=MET1_cond $X=2.385 $Y=1.87
+ $X2=1.3 $Y2=1.87
r119 20 26 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r120 20 21 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r121 18 21 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r122 15 35 87.2276 $w=2.68e-07 $l=5.95021e-07 $layer=POLY_cond $X=3.21 $Y=1.175
+ $X2=2.725 $Y2=1.42
r123 14 15 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.21 $Y=0.785
+ $X2=3.21 $Y2=1.175
r124 11 14 28.5207 $w=1.69e-07 $l=1.16189e-07 $layer=POLY_cond $X=3.175 $Y=0.685
+ $X2=3.21 $Y2=0.785
r125 11 13 86.76 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.175 $Y=0.685
+ $X2=3.175 $Y2=0.415
r126 7 35 16.3317 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.725 $Y=1.685
+ $X2=2.725 $Y2=1.42
r127 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.725 $Y=1.685
+ $X2=2.725 $Y2=2.275
r128 2 26 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r129 1 18 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%A_715_21# 1 2 9 13 17 20 22 25 29 33 36 38
+ 41 42 44 46 47 53
c83 42 0 1.06502e-19 $X=5.01 $Y=1.16
c84 13 0 8.44901e-20 $X=3.65 $Y=2.275
r85 42 54 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.022 $Y=1.16
+ $X2=5.022 $Y2=1.325
r86 42 53 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.022 $Y=1.16
+ $X2=5.022 $Y2=0.995
r87 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.16 $X2=5.01 $Y2=1.16
r88 39 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=1.16
+ $X2=4.455 $Y2=1.16
r89 39 41 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.54 $Y=1.16
+ $X2=5.01 $Y2=1.16
r90 38 46 7.45506 $w=2.07e-07 $l=1.83016e-07 $layer=LI1_cond $X=4.455 $Y=1.535
+ $X2=4.417 $Y2=1.7
r91 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=1.325
+ $X2=4.455 $Y2=1.16
r92 37 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.455 $Y=1.325
+ $X2=4.455 $Y2=1.535
r93 36 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0.995
+ $X2=4.455 $Y2=1.16
r94 36 44 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.455 $Y=0.995
+ $X2=4.455 $Y2=0.72
r95 31 46 7.45506 $w=2.07e-07 $l=1.65e-07 $layer=LI1_cond $X=4.417 $Y=1.865
+ $X2=4.417 $Y2=1.7
r96 31 33 19.0506 $w=2.43e-07 $l=4.05e-07 $layer=LI1_cond $X=4.417 $Y=1.865
+ $X2=4.417 $Y2=2.27
r97 27 44 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=4.417 $Y=0.598
+ $X2=4.417 $Y2=0.72
r98 27 29 8.13766 $w=2.43e-07 $l=1.73e-07 $layer=LI1_cond $X=4.417 $Y=0.598
+ $X2=4.417 $Y2=0.425
r99 25 48 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.9 $Y=1.7 $X2=3.65
+ $Y2=1.7
r100 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.7 $X2=3.9 $Y2=1.7
r101 22 46 0.261258 $w=3.3e-07 $l=1.22e-07 $layer=LI1_cond $X=4.295 $Y=1.7
+ $X2=4.417 $Y2=1.7
r102 22 24 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.295 $Y=1.7
+ $X2=3.9 $Y2=1.7
r103 20 54 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.05 $Y=1.985
+ $X2=5.05 $Y2=1.325
r104 17 53 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.05 $Y=0.56
+ $X2=5.05 $Y2=0.995
r105 11 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.865
+ $X2=3.65 $Y2=1.7
r106 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.65 $Y=1.865
+ $X2=3.65 $Y2=2.275
r107 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.535
+ $X2=3.65 $Y2=1.7
r108 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.65 $Y=1.535
+ $X2=3.65 $Y2=0.445
r109 2 46 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.485 $X2=4.38 $Y2=1.755
r110 2 33 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.485 $X2=4.38 $Y2=2.27
r111 1 29 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.235 $X2=4.38 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%A_560_47# 1 2 7 9 12 14 15 16 20 25 27 30 34
c90 34 0 3.17665e-20 $X=3.54 $Y=1.222
c91 30 0 1.06502e-19 $X=4.115 $Y=1.16
c92 20 0 1.48267e-19 $X=3.435 $Y=0.45
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r94 28 34 0.718145 $w=3.3e-07 $l=1.3242e-07 $layer=LI1_cond $X=3.645 $Y=1.16
+ $X2=3.54 $Y2=1.222
r95 28 30 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=3.645 $Y=1.16
+ $X2=4.115 $Y2=1.16
r96 27 33 15.1613 $w=2.96e-07 $l=3.67831e-07 $layer=LI1_cond $X=3.55 $Y=2.01
+ $X2=3.47 $Y2=2.34
r97 26 34 8.26956 $w=1.8e-07 $l=2.32946e-07 $layer=LI1_cond $X=3.55 $Y=1.45
+ $X2=3.54 $Y2=1.222
r98 26 27 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.55 $Y=1.45 $X2=3.55
+ $Y2=2.01
r99 25 34 8.26956 $w=1.8e-07 $l=2.36789e-07 $layer=LI1_cond $X=3.52 $Y=0.995
+ $X2=3.54 $Y2=1.222
r100 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.52 $Y=0.535
+ $X2=3.52 $Y2=0.995
r101 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=3.52 $Y2=0.535
r102 20 22 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.435 $Y=0.45
+ $X2=2.935 $Y2=0.45
r103 16 33 3.98214 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=2.34
+ $X2=3.47 $Y2=2.34
r104 16 18 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.295 $Y=2.34
+ $X2=2.935 $Y2=2.34
r105 14 31 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=4.515 $Y=1.16
+ $X2=4.115 $Y2=1.16
r106 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.515 $Y=1.16
+ $X2=4.59 $Y2=1.16
r107 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.16
r108 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.59 $Y=1.325
+ $X2=4.59 $Y2=1.985
r109 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=1.16
r110 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.59 $Y=0.995
+ $X2=4.59 $Y2=0.56
r111 2 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=2.065 $X2=2.935 $Y2=2.34
r112 1 22 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.235 $X2=2.935 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%VPWR 1 2 3 4 15 19 23 27 29 31 36 41 49 56
+ 57 60 63 66 69
r92 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r93 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r95 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r96 57 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r97 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 54 69 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=4.862 $Y2=2.72
r99 54 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.005 $Y=2.72
+ $X2=5.29 $Y2=2.72
r100 53 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r101 53 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r102 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 50 66 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=3.935 $Y2=2.72
r104 50 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 49 69 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.862 $Y2=2.72
r106 49 52 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.72 $Y=2.72
+ $X2=4.37 $Y2=2.72
r107 48 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r108 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r109 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r110 45 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 44 47 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r112 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r113 42 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.1 $Y2=2.72
r114 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.245 $Y=2.72
+ $X2=2.53 $Y2=2.72
r115 41 66 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.775 $Y=2.72
+ $X2=3.935 $Y2=2.72
r116 41 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.775 $Y=2.72
+ $X2=3.45 $Y2=2.72
r117 40 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r118 40 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r120 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r121 37 39 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 36 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.1 $Y2=2.72
r123 36 39 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r124 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r125 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 29 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 29 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r128 25 69 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.862 $Y=2.635
+ $X2=4.862 $Y2=2.72
r129 25 27 36.3929 $w=2.83e-07 $l=9e-07 $layer=LI1_cond $X=4.862 $Y=2.635
+ $X2=4.862 $Y2=1.735
r130 21 66 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=2.635
+ $X2=3.935 $Y2=2.72
r131 21 23 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.935 $Y=2.635
+ $X2=3.935 $Y2=2.34
r132 17 63 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2.72
r133 17 19 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=2.1 $Y=2.635
+ $X2=2.1 $Y2=2
r134 13 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r135 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r136 4 27 300 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.485 $X2=4.84 $Y2=1.735
r137 3 23 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.725
+ $Y=2.065 $X2=3.86 $Y2=2.34
r138 2 19 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r139 1 15 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%Q 1 2 9 10 11 19 30
r16 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.35 $Y=0.745
+ $X2=5.35 $Y2=1.67
r17 16 19 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.305 $Y=1.8
+ $X2=5.305 $Y2=1.835
r18 10 16 0.354598 $w=2.58e-07 $l=8e-09 $layer=LI1_cond $X=5.305 $Y=1.792
+ $X2=5.305 $Y2=1.8
r19 10 30 6.78766 $w=2.58e-07 $l=1.22e-07 $layer=LI1_cond $X=5.305 $Y=1.792
+ $X2=5.305 $Y2=1.67
r20 10 11 14.7601 $w=2.58e-07 $l=3.33e-07 $layer=LI1_cond $X=5.305 $Y=1.877
+ $X2=5.305 $Y2=2.21
r21 10 19 1.86164 $w=2.58e-07 $l=4.2e-08 $layer=LI1_cond $X=5.305 $Y=1.877
+ $X2=5.305 $Y2=1.835
r22 9 28 11.7964 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=5.305 $Y=0.51
+ $X2=5.305 $Y2=0.745
r23 2 19 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.125
+ $Y=1.485 $X2=5.26 $Y2=1.835
r24 1 9 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.26 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HD__DLXTN_1%VGND 1 2 3 4 15 19 23 25 29 31 33 38 43 53
+ 54 57 60 63 66
c86 54 0 2.71124e-20 $X=5.29 $Y=0
r87 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r88 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r89 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r90 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r91 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r92 54 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r93 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r94 51 66 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=4.867
+ $Y2=0
r95 51 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=5.29
+ $Y2=0
r96 50 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r97 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r98 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r99 47 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r100 46 49 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r101 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r102 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r103 44 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r104 43 63 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=3.91
+ $Y2=0
r105 43 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=3.45 $Y2=0
r106 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r107 42 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r108 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r109 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r110 39 41 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r111 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r112 38 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r113 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r114 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r115 31 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 27 66 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.867 $Y=0.085
+ $X2=4.867 $Y2=0
r118 27 29 23.8172 $w=2.23e-07 $l=4.65e-07 $layer=LI1_cond $X=4.867 $Y=0.085
+ $X2=4.867 $Y2=0.55
r119 26 63 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.045 $Y=0 $X2=3.91
+ $Y2=0
r120 25 66 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=4.867 $Y2=0
r121 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=4.045 $Y2=0
r122 21 63 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0
r123 21 23 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.91 $Y=0.085
+ $X2=3.91 $Y2=0.38
r124 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r125 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r126 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r127 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r128 4 29 182 $w=1.7e-07 $l=3.92874e-07 $layer=licon1_NDIFF $count=1 $X=4.665
+ $Y=0.235 $X2=4.84 $Y2=0.55
r129 3 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.725
+ $Y=0.235 $X2=3.86 $Y2=0.38
r130 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r131 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


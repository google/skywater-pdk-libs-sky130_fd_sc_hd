* File: sky130_fd_sc_hd__clkdlybuf4s18_1.spice.SKY130_FD_SC_HD__CLKDLYBUF4S18_1.pxi
* Created: Thu Aug 27 14:11:31 2020
* 
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A N_A_M1002_g N_A_M1004_g A N_A_c_67_n
+ N_A_c_68_n N_A_c_71_n PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_27_47# N_A_27_47#_M1002_s
+ N_A_27_47#_M1004_s N_A_27_47#_M1000_g N_A_27_47#_M1006_g N_A_27_47#_c_98_n
+ N_A_27_47#_c_99_n N_A_27_47#_c_100_n N_A_27_47#_c_107_n N_A_27_47#_c_101_n
+ N_A_27_47#_c_102_n N_A_27_47#_c_108_n N_A_27_47#_c_109_n N_A_27_47#_c_103_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_27_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_282_47# N_A_282_47#_M1000_d
+ N_A_282_47#_M1006_d N_A_282_47#_M1005_g N_A_282_47#_M1001_g
+ N_A_282_47#_c_163_n N_A_282_47#_c_164_n N_A_282_47#_c_165_n
+ N_A_282_47#_c_166_n N_A_282_47#_c_167_n N_A_282_47#_c_172_n
+ N_A_282_47#_c_168_n N_A_282_47#_c_169_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_282_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_394_47# N_A_394_47#_M1005_s
+ N_A_394_47#_M1001_s N_A_394_47#_M1003_g N_A_394_47#_M1007_g
+ N_A_394_47#_c_225_n N_A_394_47#_c_230_n N_A_394_47#_c_226_n
+ N_A_394_47#_c_227_n N_A_394_47#_c_231_n N_A_394_47#_c_232_n
+ N_A_394_47#_c_228_n N_A_394_47#_c_229_n N_A_394_47#_c_235_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%A_394_47#
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VPWR N_VPWR_M1004_d N_VPWR_M1001_d
+ N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n VPWR
+ N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_290_n N_VPWR_c_298_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VPWR
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%X N_X_M1003_d N_X_M1007_d X X X X X X
+ N_X_c_332_n X PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%X
x_PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VGND N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_c_347_n N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n VGND
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n
+ PM_SKY130_FD_SC_HD__CLKDLYBUF4S18_1%VGND
cc_1 VNB N_A_M1002_g 0.043678f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_c_67_n 0.0258591f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_3 VNB N_A_c_68_n 0.0123004f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.16
cc_4 VNB N_A_27_47#_M1000_g 0.0260315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_c_98_n 0.0305278f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_6 VNB N_A_27_47#_c_99_n 0.0135529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_100_n 0.0182375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_101_n 0.00275349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_102_n 0.00988333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_103_n 0.00445545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_282_47#_M1005_g 0.0266102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_282_47#_c_163_n 0.00453903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_282_47#_c_164_n 0.00503371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_282_47#_c_165_n 0.0138999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_282_47#_c_166_n 0.046472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_282_47#_c_167_n 0.00192115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_282_47#_c_168_n 0.00131782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_282_47#_c_169_n 0.00281555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_394_47#_M1003_g 0.0375015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_394_47#_c_225_n 0.00430508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_394_47#_c_226_n 0.0012699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_394_47#_c_227_n 0.00326801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_394_47#_c_228_n 0.00385296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_394_47#_c_229_n 0.0229123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_290_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0366411f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.985
cc_27 VNB N_X_c_332_n 0.0125801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_347_n 0.0055024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_348_n 0.00558109f $X=-0.19 $Y=-0.24 $X2=0.385 $Y2=1.025
cc_30 VNB N_VGND_c_349_n 0.0474987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_350_n 0.00631567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_351_n 0.0172145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_352_n 0.0182402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_353_n 0.208683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_354_n 0.00602727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_c_67_n 0.0109012f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_37 VPB N_A_c_68_n 0.00196302f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_38 VPB N_A_c_71_n 0.0248709f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.375
cc_39 VPB N_A_27_47#_M1006_g 0.0367872f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.025
cc_40 VPB N_A_27_47#_c_98_n 0.0179428f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_41 VPB N_A_27_47#_c_99_n 0.0033884f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_107_n 0.031185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_108_n 0.00223288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_109_n 0.00756198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_103_n 0.00279737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_282_47#_M1001_g 0.0376316f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.025
cc_47 VPB N_A_282_47#_c_166_n 0.0211298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_282_47#_c_172_n 0.00707847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_282_47#_c_168_n 0.00982875f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_394_47#_c_230_n 0.00817407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_394_47#_c_231_n 0.0104266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_394_47#_c_232_n 0.00409921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_394_47#_c_228_n 0.0012917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_394_47#_c_229_n 0.00886211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_394_47#_c_235_n 0.021413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_291_n 0.00558649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_292_n 0.00563065f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.025
cc_58 VPB N_VPWR_c_293_n 0.0498889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_294_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_295_n 0.0178539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_296_n 0.0189199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_290_n 0.0528294f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_298_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB X 0.0194334f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_65 VPB X 0.0292395f $X=-0.19 $Y=1.305 $X2=0.385 $Y2=1.16
cc_66 N_A_M1002_g N_A_27_47#_M1000_g 0.0100164f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_67 N_A_c_71_n N_A_27_47#_M1006_g 0.0146572f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_68 N_A_c_67_n N_A_27_47#_c_98_n 0.0225951f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_68_n N_A_27_47#_c_98_n 3.0562e-19 $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_M1002_g N_A_27_47#_c_100_n 0.0134301f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_c_71_n N_A_27_47#_c_107_n 0.0163421f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_A_27_47#_c_101_n 0.0101783f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A_c_68_n N_A_27_47#_c_101_n 0.00875068f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_A_27_47#_c_102_n 0.00418154f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A_c_67_n N_A_27_47#_c_102_n 0.00438111f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_27_47#_c_102_n 0.0272348f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_68_n N_A_27_47#_c_108_n 0.00875068f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_c_71_n N_A_27_47#_c_108_n 0.0125516f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_A_27_47#_c_109_n 0.00431459f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_c_68_n N_A_27_47#_c_109_n 0.0243826f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_c_71_n N_A_27_47#_c_109_n 0.00419718f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_A_27_47#_c_103_n 0.0048366f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_c_67_n N_A_27_47#_c_103_n 0.00570434f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_c_68_n N_A_27_47#_c_103_n 0.0225095f $X=0.385 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_71_n N_VPWR_c_291_n 0.00916932f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_86 N_A_c_71_n N_VPWR_c_295_n 0.0054895f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_87 N_A_c_71_n N_VPWR_c_290_n 0.0114789f $X=0.385 $Y=1.375 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_VGND_c_347_n 0.00341797f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VGND_c_351_n 0.00424868f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VGND_c_353_n 0.00741185f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1000_g N_A_282_47#_c_163_n 0.00977878f $X=1.32 $Y=0.56 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_M1000_g N_A_282_47#_c_164_n 0.00363648f $X=1.32 $Y=0.56 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_c_103_n N_A_282_47#_c_164_n 0.00784898f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_M1000_g N_A_282_47#_c_166_n 0.00493946f $X=1.32 $Y=0.56 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_M1000_g N_A_282_47#_c_167_n 0.0058351f $X=1.32 $Y=0.56 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_M1006_g N_A_282_47#_c_172_n 0.0131002f $X=1.32 $Y=2.075 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_99_n N_A_282_47#_c_168_n 0.012754f $X=1.32 $Y=1.2 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_108_n N_A_282_47#_c_168_n 0.00825693f $X=0.72 $Y=1.58 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_103_n N_A_282_47#_c_168_n 0.0109765f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_99_n N_A_282_47#_c_169_n 0.00290025f $X=1.32 $Y=1.2 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_103_n N_A_282_47#_c_169_n 0.00936769f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_108_n N_VPWR_M1004_d 0.0202644f $X=0.72 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_27_47#_M1006_g N_VPWR_c_291_n 0.0091189f $X=1.32 $Y=2.075 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_98_n N_VPWR_c_291_n 6.91023e-19 $X=1.23 $Y=1.2 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_108_n N_VPWR_c_291_n 0.027505f $X=0.72 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1006_g N_VPWR_c_293_n 0.00666027f $X=1.32 $Y=2.075 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_107_n N_VPWR_c_295_n 0.0210489f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1004_s N_VPWR_c_290_n 0.00213418f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1006_g N_VPWR_c_290_n 0.0138366f $X=1.32 $Y=2.075 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_107_n N_VPWR_c_290_n 0.0124497f $X=0.26 $Y=1.965 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_101_n N_VGND_M1002_d 0.0121993f $X=0.72 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_27_47#_M1000_g N_VGND_c_347_n 0.00539845f $X=1.32 $Y=0.56 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_98_n N_VGND_c_347_n 5.9826e-19 $X=1.23 $Y=1.2 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_101_n N_VGND_c_347_n 0.0255398f $X=0.72 $Y=0.8 $X2=0 $Y2=0
cc_115 N_A_27_47#_M1000_g N_VGND_c_349_n 0.00666027f $X=1.32 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_101_n N_VGND_c_349_n 0.00463496f $X=0.72 $Y=0.8 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_100_n N_VGND_c_351_n 0.0209424f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_101_n N_VGND_c_351_n 0.00239555f $X=0.72 $Y=0.8 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1002_s N_VGND_c_353_n 0.00213418f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_120 N_A_27_47#_M1000_g N_VGND_c_353_n 0.0138366f $X=1.32 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_100_n N_VGND_c_353_n 0.0124245f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_101_n N_VGND_c_353_n 0.01386f $X=0.72 $Y=0.8 $X2=0 $Y2=0
cc_123 N_A_282_47#_M1005_g N_A_394_47#_M1003_g 0.0120269f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_124 N_A_282_47#_M1005_g N_A_394_47#_c_225_n 0.0157423f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_125 N_A_282_47#_c_163_n N_A_394_47#_c_225_n 0.0385933f $X=1.55 $Y=0.38 $X2=0
+ $Y2=0
cc_126 N_A_282_47#_M1001_g N_A_394_47#_c_230_n 0.0241909f $X=2.325 $Y=2.075
+ $X2=0 $Y2=0
cc_127 N_A_282_47#_c_168_n N_A_394_47#_c_230_n 0.072274f $X=1.572 $Y=1.835 $X2=0
+ $Y2=0
cc_128 N_A_282_47#_M1005_g N_A_394_47#_c_226_n 0.0118486f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_129 N_A_282_47#_c_165_n N_A_394_47#_c_226_n 0.0276647f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_282_47#_c_166_n N_A_394_47#_c_226_n 0.00765601f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_131 N_A_282_47#_M1005_g N_A_394_47#_c_227_n 0.00418154f $X=2.325 $Y=0.56
+ $X2=0 $Y2=0
cc_132 N_A_282_47#_c_165_n N_A_394_47#_c_227_n 0.0239186f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_133 N_A_282_47#_c_166_n N_A_394_47#_c_227_n 0.00522157f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_282_47#_c_167_n N_A_394_47#_c_227_n 0.0148501f $X=1.572 $Y=0.825
+ $X2=0 $Y2=0
cc_135 N_A_282_47#_M1001_g N_A_394_47#_c_231_n 0.0147962f $X=2.325 $Y=2.075
+ $X2=0 $Y2=0
cc_136 N_A_282_47#_c_165_n N_A_394_47#_c_231_n 0.0300881f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_282_47#_c_166_n N_A_394_47#_c_231_n 0.00868919f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_282_47#_M1001_g N_A_394_47#_c_232_n 0.00419718f $X=2.325 $Y=2.075
+ $X2=0 $Y2=0
cc_139 N_A_282_47#_c_165_n N_A_394_47#_c_232_n 0.0270768f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_282_47#_c_166_n N_A_394_47#_c_232_n 0.00605921f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_282_47#_c_168_n N_A_394_47#_c_232_n 0.014358f $X=1.572 $Y=1.835 $X2=0
+ $Y2=0
cc_142 N_A_282_47#_M1005_g N_A_394_47#_c_228_n 0.00266247f $X=2.325 $Y=0.56
+ $X2=0 $Y2=0
cc_143 N_A_282_47#_M1001_g N_A_394_47#_c_228_n 8.74243e-19 $X=2.325 $Y=2.075
+ $X2=0 $Y2=0
cc_144 N_A_282_47#_c_165_n N_A_394_47#_c_228_n 0.0162311f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_282_47#_c_166_n N_A_394_47#_c_228_n 0.00546854f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_146 N_A_282_47#_c_166_n N_A_394_47#_c_229_n 0.0233501f $X=2.52 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_282_47#_M1001_g N_A_394_47#_c_235_n 0.0149063f $X=2.325 $Y=2.075
+ $X2=0 $Y2=0
cc_148 N_A_282_47#_c_172_n N_VPWR_c_291_n 0.0228359f $X=1.55 $Y=1.97 $X2=0 $Y2=0
cc_149 N_A_282_47#_M1001_g N_VPWR_c_292_n 0.0100242f $X=2.325 $Y=2.075 $X2=0
+ $Y2=0
cc_150 N_A_282_47#_M1001_g N_VPWR_c_293_n 0.00666027f $X=2.325 $Y=2.075 $X2=0
+ $Y2=0
cc_151 N_A_282_47#_c_172_n N_VPWR_c_293_n 0.0242182f $X=1.55 $Y=1.97 $X2=0 $Y2=0
cc_152 N_A_282_47#_M1006_d N_VPWR_c_290_n 0.00213418f $X=1.41 $Y=1.665 $X2=0
+ $Y2=0
cc_153 N_A_282_47#_M1001_g N_VPWR_c_290_n 0.0138366f $X=2.325 $Y=2.075 $X2=0
+ $Y2=0
cc_154 N_A_282_47#_c_172_n N_VPWR_c_290_n 0.0141671f $X=1.55 $Y=1.97 $X2=0 $Y2=0
cc_155 N_A_282_47#_c_163_n N_VGND_c_347_n 0.0102124f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_156 N_A_282_47#_M1005_g N_VGND_c_348_n 0.0056082f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_157 N_A_282_47#_M1005_g N_VGND_c_349_n 0.00512166f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_158 N_A_282_47#_c_163_n N_VGND_c_349_n 0.0241445f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_159 N_A_282_47#_M1000_d N_VGND_c_353_n 0.00213418f $X=1.41 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_282_47#_M1005_g N_VGND_c_353_n 0.00889447f $X=2.325 $Y=0.56 $X2=0
+ $Y2=0
cc_161 N_A_282_47#_c_163_n N_VGND_c_353_n 0.0141471f $X=1.55 $Y=0.38 $X2=0 $Y2=0
cc_162 N_A_394_47#_c_231_n N_VPWR_M1001_d 0.00879448f $X=2.855 $Y=1.505 $X2=0
+ $Y2=0
cc_163 N_A_394_47#_c_230_n N_VPWR_c_292_n 0.0257926f $X=2.095 $Y=1.965 $X2=0
+ $Y2=0
cc_164 N_A_394_47#_c_231_n N_VPWR_c_292_n 0.0281787f $X=2.855 $Y=1.505 $X2=0
+ $Y2=0
cc_165 N_A_394_47#_c_229_n N_VPWR_c_292_n 4.5311e-19 $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_394_47#_c_235_n N_VPWR_c_292_n 0.0096431f $X=3.095 $Y=1.375 $X2=0
+ $Y2=0
cc_167 N_A_394_47#_c_230_n N_VPWR_c_293_n 0.0210489f $X=2.095 $Y=1.965 $X2=0
+ $Y2=0
cc_168 N_A_394_47#_c_235_n N_VPWR_c_296_n 0.0054895f $X=3.095 $Y=1.375 $X2=0
+ $Y2=0
cc_169 N_A_394_47#_M1001_s N_VPWR_c_290_n 0.00213418f $X=1.97 $Y=1.665 $X2=0
+ $Y2=0
cc_170 N_A_394_47#_c_230_n N_VPWR_c_290_n 0.0124497f $X=2.095 $Y=1.965 $X2=0
+ $Y2=0
cc_171 N_A_394_47#_c_235_n N_VPWR_c_290_n 0.0115355f $X=3.095 $Y=1.375 $X2=0
+ $Y2=0
cc_172 N_A_394_47#_M1003_g X 0.0310689f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A_394_47#_c_226_n X 0.0138643f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_174 N_A_394_47#_c_231_n X 0.0137182f $X=2.855 $Y=1.505 $X2=0 $Y2=0
cc_175 N_A_394_47#_c_228_n X 0.0410231f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A_394_47#_c_235_n X 0.00933827f $X=3.095 $Y=1.375 $X2=0 $Y2=0
cc_177 N_A_394_47#_M1003_g N_X_c_332_n 0.00516929f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A_394_47#_c_226_n N_VGND_M1005_d 0.0143915f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_179 N_A_394_47#_M1003_g N_VGND_c_348_n 0.00604549f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_394_47#_c_225_n N_VGND_c_348_n 0.0106097f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_181 N_A_394_47#_c_226_n N_VGND_c_348_n 0.0271231f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_182 N_A_394_47#_c_229_n N_VGND_c_348_n 3.7903e-19 $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_394_47#_c_225_n N_VGND_c_349_n 0.0209424f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_184 N_A_394_47#_c_226_n N_VGND_c_349_n 0.00607688f $X=2.855 $Y=0.8 $X2=0
+ $Y2=0
cc_185 N_A_394_47#_M1003_g N_VGND_c_352_n 0.00432943f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_186 N_A_394_47#_c_226_n N_VGND_c_352_n 0.0024529f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_187 N_A_394_47#_M1005_s N_VGND_c_353_n 0.00213418f $X=1.97 $Y=0.235 $X2=0
+ $Y2=0
cc_188 N_A_394_47#_M1003_g N_VGND_c_353_n 0.0079683f $X=3.17 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_A_394_47#_c_225_n N_VGND_c_353_n 0.0124245f $X=2.095 $Y=0.38 $X2=0
+ $Y2=0
cc_190 N_A_394_47#_c_226_n N_VGND_c_353_n 0.0164916f $X=2.855 $Y=0.8 $X2=0 $Y2=0
cc_191 N_VPWR_c_290_n N_X_M1007_d 0.00213418f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_296_n X 0.0239326f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_290_n X 0.0139953f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_194 N_X_c_332_n N_VGND_c_352_n 0.0232369f $X=3.477 $Y=0.4 $X2=0 $Y2=0
cc_195 N_X_M1003_d N_VGND_c_353_n 0.00213443f $X=3.245 $Y=0.235 $X2=0 $Y2=0
cc_196 N_X_c_332_n N_VGND_c_353_n 0.0140906f $X=3.477 $Y=0.4 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__a2111oi_4.spice
* Created: Tue Sep  1 18:50:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a2111oi_4.pex.spice"
.subckt sky130_fd_sc_hd__a2111oi_4  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_D1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.182
+ AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2 SB=75005.1
+ A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_D1_M1009_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.08775 PD=0.93 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6 SB=75004.7
+ A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1009_d N_D1_M1016_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1 SB=75004.3
+ A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_D1_M1027_g N_Y_M1016_s VNB NSHORT L=0.15 W=0.65 AD=0.117
+ AS=0.091 PD=1.01 PS=0.93 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75001.5 SB=75003.8
+ A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1008_d N_C1_M1008_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.117 PD=0.93 PS=1.01 NRD=0 NRS=0 M=1 R=4.33333 SA=75002 SB=75003.3
+ A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1008_d N_C1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4 SB=75002.9
+ A=0.0975 P=1.6 MULT=1
MM1021 N_Y_M1021_d N_C1_M1021_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9 SB=75002.5
+ A=0.0975 P=1.6 MULT=1
MM1036 N_Y_M1021_d N_C1_M1036_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.12675 PD=0.93 PS=1.04 NRD=0 NRS=11.076 M=1 R=4.33333 SA=75003.3 SB=75002
+ A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1036_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.12675 PD=0.93 PS=1.04 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75003.8 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1001_d N_B1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.3 SB=75001.1
+ A=0.0975 P=1.6 MULT=1
MM1029 N_Y_M1029_d N_B1_M1029_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75004.7 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1037 N_Y_M1029_d N_B1_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.182 PD=0.93 PS=1.86 NRD=0 NRS=0 M=1 R=4.33333 SA=75005.1 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1017 N_A_1205_47#_M1017_d N_A1_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.091 PD=1.86 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1020 N_A_1205_47#_M1020_d N_A1_M1020_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1034 N_A_1205_47#_M1020_d N_A1_M1034_g N_Y_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1038 N_A_1205_47#_M1038_d N_A1_M1038_g N_Y_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.121875 AS=0.091 PD=1.025 PS=0.93 NRD=16.608 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75002 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_1205_47#_M1038_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.121875 PD=0.93 PS=1.025 NRD=0 NRS=0.912 M=1 R=4.33333 SA=75002
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1022 N_VGND_M1006_d N_A2_M1022_g N_A_1205_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_A2_M1024_g N_A_1205_47#_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1039 N_VGND_M1024_d N_A2_M1039_g N_A_1205_47#_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.17225 PD=0.93 PS=1.83 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_28_297#_M1003_d N_D1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75003.2 A=0.15 P=2.3 MULT=1
MM1014 N_A_28_297#_M1014_d N_D1_M1014_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75002.8 A=0.15 P=2.3 MULT=1
MM1015 N_A_28_297#_M1014_d N_D1_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75002.3
+ A=0.15 P=2.3 MULT=1
MM1032 N_A_28_297#_M1032_d N_D1_M1032_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1005 N_A_28_297#_M1032_d N_C1_M1005_g N_A_455_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75001.5 A=0.15 P=2.3 MULT=1
MM1011 N_A_28_297#_M1011_d N_C1_M1011_g N_A_455_297#_M1005_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3
+ SB=75001 A=0.15 P=2.3 MULT=1
MM1023 N_A_28_297#_M1011_d N_C1_M1023_g N_A_455_297#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1028 N_A_28_297#_M1028_d N_C1_M1028_g N_A_455_297#_M1023_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75003.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
MM1012 N_A_821_297#_M1012_d N_B1_M1012_g N_A_455_297#_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.26 AS=0.14 PD=2.52 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75005.2 A=0.15 P=2.3 MULT=1
MM1013 N_A_821_297#_M1013_d N_B1_M1013_g N_A_455_297#_M1012_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75004.7 A=0.15 P=2.3 MULT=1
MM1025 N_A_821_297#_M1013_d N_B1_M1025_g N_A_455_297#_M1025_s VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001
+ SB=75004.3 A=0.15 P=2.3 MULT=1
MM1031 N_A_821_297#_M1031_d N_B1_M1031_g N_A_455_297#_M1025_s VPB PHIGHVT L=0.15
+ W=1 AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=1.9503 NRS=0 M=1 R=6.66667 SA=75001.5
+ SB=75003.9 A=0.15 P=2.3 MULT=1
MM1018 N_A_821_297#_M1031_d N_A1_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.9
+ SB=75003.4 A=0.15 P=2.3 MULT=1
MM1026 N_A_821_297#_M1026_d N_A1_M1026_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.3 SB=75003
+ A=0.15 P=2.3 MULT=1
MM1033 N_A_821_297#_M1026_d N_A1_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.8 SB=75002.6
+ A=0.15 P=2.3 MULT=1
MM1035 N_A_821_297#_M1035_d N_A1_M1035_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2 AS=0.15 PD=1.4 PS=1.3 NRD=4.9053 NRS=3.9203 M=1 R=6.66667 SA=75003.2
+ SB=75002.1 A=0.15 P=2.3 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_821_297#_M1035_d VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.2 PD=1.28 PS=1.4 NRD=0 NRS=18.715 M=1 R=6.66667 SA=75003.8
+ SB=75001.6 A=0.15 P=2.3 MULT=1
MM1004 N_VPWR_M1000_d N_A2_M1004_g N_A_821_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.185 PD=1.28 PS=1.37 NRD=0 NRS=7.8603 M=1 R=6.66667 SA=75004.2
+ SB=75001.1 A=0.15 P=2.3 MULT=1
MM1019 N_VPWR_M1019_d N_A2_M1019_g N_A_821_297#_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.185 PD=1.28 PS=1.37 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75004.7
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1030 N_VPWR_M1019_d N_A2_M1030_g N_A_821_297#_M1030_s VPB PHIGHVT L=0.15 W=1
+ AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=6.66667 SA=75005.2
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX40_noxref VNB VPB NWDIODE A=16.8525 P=24.21
*
.include "sky130_fd_sc_hd__a2111oi_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__nand2_2.spice
* Created: Tue Sep  1 19:15:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__nand2_2.pex.spice"
.subckt sky130_fd_sc_hd__nand2_2  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_B_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1007_d N_B_M1007_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_47#_M1007_d N_A_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_A_M1004_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.26
+ AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2 SB=75001.4
+ A=0.15 P=2.3 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6 SB=75001 A=0.15
+ P=2.3 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=6.66667 SA=75001 SB=75000.6 A=0.15
+ P=2.3 MULT=1
MM1006 N_Y_M1000_d N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1 AD=0.135
+ AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=6.66667 SA=75001.4 SB=75000.2 A=0.15
+ P=2.3 MULT=1
DX8_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hd__nand2_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_hd__o2bb2a_2.spice
* Created: Thu Aug 27 14:38:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__o2bb2a_2.pex.spice"
.subckt sky130_fd_sc_hd__o2bb2a_2  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_84_21#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.08775 PD=1.87 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_84_21#_M1004_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.119825 AS=0.08775 PD=1.19065 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1003 A_294_47# N_A1_N_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0774252 PD=0.735 PS=0.769346 NRD=29.28 NRS=8.568 M=1 R=2.8
+ SA=75001.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_295_369#_M1007_d N_A2_N_M1007_g A_294_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.06615 PD=1.36 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_581_47#_M1013_d N_A_295_369#_M1013_g N_A_84_21#_M1013_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B2_M1005_g N_A_581_47#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_581_47#_M1008_d N_B1_M1008_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_84_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.285 PD=1.27 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 N_X_M1002_d N_A_84_21#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1
+ AD=0.135 AS=0.187805 PD=1.27 PS=1.62805 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.6
+ SB=75001.9 A=0.15 P=2.3 MULT=1
MM1001 N_A_295_369#_M1001_d N_A1_N_M1001_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.173 AS=0.120195 PD=1.4 PS=1.04195 NRD=66.2708 NRS=18.4589 M=1
+ R=4.26667 SA=75001.1 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A2_N_M1006_g N_A_295_369#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2272 AS=0.173 PD=1.35 PS=1.4 NRD=61.5625 NRS=66.2708 M=1 R=4.26667
+ SA=75001.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1009 N_A_84_21#_M1009_d N_A_295_369#_M1009_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0928 AS=0.2272 PD=0.93 PS=1.35 NRD=0 NRS=70.7821 M=1 R=4.26667
+ SA=75002.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1012 A_665_369# N_B2_M1012_g N_A_84_21#_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0864 AS=0.0928 PD=0.91 PS=0.93 NRD=24.625 NRS=4.6098 M=1 R=4.26667
+ SA=75003 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_B1_M1011_g A_665_369# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=24.625 M=1 R=4.26667 SA=75003.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hd__o2bb2a_2.pxi.spice"
*
.ends
*
*

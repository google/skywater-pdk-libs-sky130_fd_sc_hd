* File: sky130_fd_sc_hd__and3_1.pex.spice
* Created: Tue Sep  1 18:57:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND3_1%A 3 6 8 11 13
r27 11 14 67.3385 $w=4.2e-07 $l=3.25e-07 $layer=POLY_cond $X=0.335 $Y=0.93
+ $X2=0.335 $Y2=1.255
r28 11 13 50.7863 $w=4.2e-07 $l=2e-07 $layer=POLY_cond $X=0.335 $Y=0.93
+ $X2=0.335 $Y2=0.73
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=0.93 $X2=0.26 $Y2=0.93
r30 6 14 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.71
+ $X2=0.47 $Y2=1.255
r31 3 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.445 $X2=0.47
+ $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%B 3 8 10 11 14
r39 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.295
+ $X2=0.95 $Y2=2.13
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.295 $X2=0.95 $Y2=2.295
r41 11 15 6.77908 $w=3.38e-07 $l=2e-07 $layer=LI1_cond $X=1.15 $Y=2.295 $X2=0.95
+ $Y2=2.295
r42 9 10 39.4735 $w=2.1e-07 $l=1.25e-07 $layer=POLY_cond $X=0.86 $Y=1.285
+ $X2=0.86 $Y2=1.41
r43 8 16 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.89 $Y=1.71 $X2=0.89
+ $Y2=2.13
r44 8 10 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.89 $Y=1.71 $X2=0.89
+ $Y2=1.41
r45 3 9 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.83 $Y=0.445 $X2=0.83
+ $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%C 1 3 4 6 8 17 18
c46 4 0 2.56587e-19 $X=1.355 $Y=1.295
r47 17 18 3.37884 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.31 $Y=0.85 $X2=1.31
+ $Y2=0.79
r48 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.13 $X2=1.31 $Y2=1.13
r49 8 13 9.35923 $w=3.28e-07 $l=2.68e-07 $layer=LI1_cond $X=1.31 $Y=0.862
+ $X2=1.31 $Y2=1.13
r50 8 17 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=1.31 $Y=0.862
+ $X2=1.31 $Y2=0.85
r51 8 18 0.720909 $w=2.2e-07 $l=1.3e-08 $layer=LI1_cond $X=1.255 $Y=0.777
+ $X2=1.255 $Y2=0.79
r52 4 12 39.2307 $w=2.57e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.28 $Y2=1.13
r53 4 6 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.355 $Y2=1.71
r54 1 12 83.3047 $w=2.57e-07 $l=4.42719e-07 $layer=POLY_cond $X=1.19 $Y=0.73
+ $X2=1.28 $Y2=1.13
r55 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.19 $Y=0.73 $X2=1.19
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%A_27_47# 1 2 3 12 15 17 23 25 26 28 29 30 35
+ 36 40
c87 28 0 1.71644e-19 $X=0.89 $Y=1.19
r88 36 41 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=1.79 $Y2=1.325
r89 36 40 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.16
+ $X2=1.79 $Y2=0.995
r90 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.16 $X2=1.79 $Y2=1.16
r91 33 35 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.76 $Y=1.385
+ $X2=1.76 $Y2=1.16
r92 30 38 6.20793 $w=5e-07 $l=2.54323e-07 $layer=LI1_cond $X=1.1 $Y=1.635
+ $X2=0.89 $Y2=1.537
r93 30 32 1.07647 $w=4.98e-07 $l=4.5e-08 $layer=LI1_cond $X=1.1 $Y=1.635
+ $X2=1.145 $Y2=1.635
r94 29 33 5.10332 $w=5.79e-07 $l=3.02076e-07 $layer=LI1_cond $X=1.645 $Y=1.635
+ $X2=1.76 $Y2=1.385
r95 29 32 11.9608 $w=4.98e-07 $l=5e-07 $layer=LI1_cond $X=1.645 $Y=1.635
+ $X2=1.145 $Y2=1.635
r96 28 38 5.00804 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=0.89 $Y=1.19
+ $X2=0.89 $Y2=1.537
r97 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.89 $Y=0.465
+ $X2=0.89 $Y2=1.19
r98 25 38 9.51026 $w=3.52e-07 $l=3.403e-07 $layer=LI1_cond $X=0.71 $Y=1.275
+ $X2=0.89 $Y2=1.537
r99 25 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.71 $Y=1.275
+ $X2=0.345 $Y2=1.275
r100 21 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=1.36
+ $X2=0.345 $Y2=1.275
r101 21 23 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=0.215 $Y=1.36
+ $X2=0.215 $Y2=1.645
r102 17 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=0.38
+ $X2=0.89 $Y2=0.465
r103 17 19 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.805 $Y=0.38
+ $X2=0.26 $Y2=0.38
r104 15 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.83 $Y=1.985
+ $X2=1.83 $Y2=1.325
r105 12 40 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.83 $Y=0.56
+ $X2=1.83 $Y2=0.995
r106 3 32 600 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=1.5 $X2=1.145 $Y2=1.7
r107 2 23 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.5 $X2=0.26 $Y2=1.645
r108 1 19 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%VPWR 1 2 9 11 13 20 21 26 29
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 24 26 20.6307 $w=5.47e-07 $l=1.04608e-06 $layer=LI1_cond $X=0.68 $Y=1.795
+ $X2=0.422 $Y2=2.72
r35 21 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 18 29 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.77 $Y=2.72
+ $X2=1.642 $Y2=2.72
r38 18 20 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.77 $Y=2.72 $X2=2.07
+ $Y2=2.72
r39 17 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 16 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r42 13 29 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.642 $Y2=2.72
r43 13 16 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.515 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 11 17 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r45 11 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 7 29 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.642 $Y=2.635
+ $X2=1.642 $Y2=2.72
r47 7 9 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.642 $Y=2.635
+ $X2=1.642 $Y2=2.34
r48 2 9 600 $w=1.7e-07 $l=9.30161e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.5 $X2=1.62 $Y2=2.34
r49 1 24 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.5 $X2=0.68 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%X 1 2 9 10 12 13 14 22
r18 14 22 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=2.077 $Y=2.21
+ $X2=2.077 $Y2=1.93
r19 11 13 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=2.085 $Y=0.605
+ $X2=2.085 $Y2=0.51
r20 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.085 $Y=0.605
+ $X2=2.085 $Y2=0.735
r21 10 12 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.13 $Y=1.765
+ $X2=2.13 $Y2=0.735
r22 9 22 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.077 $Y=1.902
+ $X2=2.077 $Y2=1.93
r23 9 10 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.077 $Y=1.902
+ $X2=2.077 $Y2=1.765
r24 2 22 300 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.485 $X2=2.04 $Y2=1.93
r25 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__AND3_1%VGND 1 6 8 10 17 18 21
c31 10 0 8.49422e-20 $X=1.535 $Y=0
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r33 18 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r34 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r35 15 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.66
+ $Y2=0
r36 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.07
+ $Y2=0
r37 10 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.66
+ $Y2=0
r38 10 12 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=1.535 $Y=0 $X2=0.23
+ $Y2=0
r39 8 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r40 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r41 4 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0
r42 4 6 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.66 $Y=0.085
+ $X2=1.66 $Y2=0.46
r43 1 6 182 $w=1.7e-07 $l=4.53762e-07 $layer=licon1_NDIFF $count=1 $X=1.265
+ $Y=0.235 $X2=1.62 $Y2=0.46
.ends


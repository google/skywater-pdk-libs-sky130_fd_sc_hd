* File: sky130_fd_sc_hd__o21a_2.pex.spice
* Created: Tue Sep  1 19:21:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O21A_2%A_79_21# 1 2 7 9 12 14 16 19 24 27 28 29 30
+ 32 34 36 42 46
c75 34 0 1.12844e-19 $X=2.095 $Y=2.005
r76 45 46 60.9673 $w=3.36e-07 $l=4.25e-07 $layer=POLY_cond $X=0.47 $Y=1.165
+ $X2=0.895 $Y2=1.165
r77 34 44 3.15253 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=2.095 $Y=2.005
+ $X2=2.095 $Y2=1.895
r78 34 36 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.095 $Y=2.005
+ $X2=2.095 $Y2=2.3
r79 30 32 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.63 $Y=0.635
+ $X2=1.63 $Y2=0.385
r80 28 44 3.72571 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.965 $Y=1.895
+ $X2=2.095 $Y2=1.895
r81 28 29 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=1.965 $Y=1.895
+ $X2=1.275 $Y2=1.895
r82 27 29 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.19 $Y=1.785
+ $X2=1.275 $Y2=1.895
r83 27 42 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.19 $Y=1.785
+ $X2=1.19 $Y2=1.33
r84 25 46 30.8423 $w=3.36e-07 $l=2.15e-07 $layer=POLY_cond $X=1.11 $Y=1.165
+ $X2=0.895 $Y2=1.165
r85 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.16 $X2=1.11 $Y2=1.16
r86 22 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=1.165
+ $X2=1.11 $Y2=1.33
r87 22 24 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.11 $Y=1.165
+ $X2=1.11 $Y2=1.16
r88 21 30 28.133 $w=2.03e-07 $l=5.2e-07 $layer=LI1_cond $X=1.11 $Y=0.737
+ $X2=1.63 $Y2=0.737
r89 21 24 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.11 $Y=0.84
+ $X2=1.11 $Y2=1.16
r90 17 46 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.895 $Y=1.335
+ $X2=0.895 $Y2=1.165
r91 17 19 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.895 $Y=1.335
+ $X2=0.895 $Y2=1.985
r92 14 46 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=1.165
r93 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.895 $Y=0.995
+ $X2=0.895 $Y2=0.56
r94 10 45 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.47 $Y=1.335
+ $X2=0.47 $Y2=1.165
r95 10 12 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.47 $Y=1.335
+ $X2=0.47 $Y2=1.985
r96 7 45 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.165
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
r98 2 44 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.485 $X2=2.06 $Y2=1.92
r99 2 36 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.485 $X2=2.06 $Y2=2.3
r100 1 32 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.63 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%B1 3 6 8 11 12 13
r36 11 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.722 $Y=1.16
+ $X2=1.722 $Y2=1.325
r37 11 13 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.722 $Y=1.16
+ $X2=1.722 $Y2=0.995
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.16 $X2=1.69 $Y2=1.16
r39 8 12 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=1.53 $X2=1.65
+ $Y2=1.16
r40 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.845 $Y=1.985
+ $X2=1.845 $Y2=1.325
r41 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.845 $Y=0.56
+ $X2=1.845 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%A2 3 6 8 11 14 17
r44 13 14 25.4279 $w=2.03e-07 $l=4.7e-07 $layer=LI1_cond $X=2.507 $Y=1.4
+ $X2=2.507 $Y2=1.87
r45 11 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.16
+ $X2=2.295 $Y2=1.325
r46 11 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.16
+ $X2=2.295 $Y2=0.995
r47 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.16 $X2=2.295 $Y2=1.16
r48 8 13 7.60723 $w=3.75e-07 $l=2.33495e-07 $layer=LI1_cond $X=2.405 $Y=1.212
+ $X2=2.507 $Y2=1.4
r49 8 10 3.3805 $w=3.73e-07 $l=1.1e-07 $layer=LI1_cond $X=2.405 $Y=1.212
+ $X2=2.295 $Y2=1.212
r50 6 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.275 $Y=1.985
+ $X2=2.275 $Y2=1.325
r51 3 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.275 $Y=0.56
+ $X2=2.275 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%A1 1 3 6 8 13
c26 6 0 1.12844e-19 $X=2.745 $Y=1.985
r27 10 13 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.745 $Y=1.16
+ $X2=2.975 $Y2=1.16
r28 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.16 $X2=2.975 $Y2=1.16
r29 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.16
r30 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.745 $Y=1.325
+ $X2=2.745 $Y2=1.985
r31 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=0.995
+ $X2=2.745 $Y2=1.16
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.745 $Y=0.995
+ $X2=2.745 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%VPWR 1 2 3 10 12 14 16 18 25 36 39 42
r49 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 38 39 10.2865 $w=6.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.495
+ $X2=1.795 $Y2=2.495
r51 34 38 0.385832 $w=6.18e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=2.495
+ $X2=1.63 $Y2=2.495
r52 34 36 19.9323 $w=6.18e-07 $l=6.65e-07 $layer=LI1_cond $X=1.61 $Y=2.495
+ $X2=0.945 $Y2=2.495
r53 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 29 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 29 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 28 39 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=1.795 $Y2=2.72
r57 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 25 41 4.719 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.007 $Y2=2.72
r59 25 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 24 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 23 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=0.945 $Y2=2.72
r62 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 21 31 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r64 21 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 18 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 14 41 3.00502 $w=3.25e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.957 $Y=2.635
+ $X2=3.007 $Y2=2.72
r68 14 16 28.1905 $w=3.23e-07 $l=7.95e-07 $layer=LI1_cond $X=2.957 $Y=2.635
+ $X2=2.957 $Y2=1.84
r69 10 31 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r70 10 12 37.059 $w=2.53e-07 $l=8.2e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=1.815
r71 3 16 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=1.485 $X2=2.96 $Y2=1.84
r72 2 38 300 $w=1.7e-07 $l=1.13812e-06 $layer=licon1_PDIFF $count=2 $X=0.97
+ $Y=1.485 $X2=1.63 $Y2=2.34
r73 1 12 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%X 1 2 7 10
r15 10 13 65.3835 $w=2.43e-07 $l=1.39e-06 $layer=LI1_cond $X=0.652 $Y=0.42
+ $X2=0.652 $Y2=1.81
r16 7 13 18.8154 $w=2.43e-07 $l=4e-07 $layer=LI1_cond $X=0.652 $Y=2.21 $X2=0.652
+ $Y2=1.81
r17 2 13 300 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_PDIFF $count=2 $X=0.545
+ $Y=1.485 $X2=0.68 $Y2=1.81
r18 1 10 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r54 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r55 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.51
+ $Y2=0
r56 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.99
+ $Y2=0
r57 33 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r58 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r59 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r60 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.11
+ $Y2=0
r61 30 32 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=2.07
+ $Y2=0
r62 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.51
+ $Y2=0
r63 29 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.07
+ $Y2=0
r64 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r65 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r66 25 40 3.93736 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r67 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r68 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.11
+ $Y2=0
r69 24 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.69
+ $Y2=0
r70 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r71 22 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r72 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0
r73 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.51 $Y=0.085
+ $X2=2.51 $Y2=0.38
r74 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0
r75 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0.38
r76 10 40 3.14078 $w=2.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.172 $Y2=0
r77 10 12 14.1654 $w=2.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=0.085
+ $X2=0.225 $Y2=0.38
r78 3 20 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.51 $Y2=0.38
r79 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.11 $Y2=0.38
r80 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O21A_2%A_384_47# 1 2 7 10 15
r20 10 12 3.69697 $w=2.08e-07 $l=7e-08 $layer=LI1_cond $X=2.07 $Y=0.66 $X2=2.07
+ $Y2=0.73
r21 8 12 1.31963 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=2.175 $Y=0.73
+ $X2=2.07 $Y2=0.73
r22 7 15 2.93349 $w=2.73e-07 $l=7e-08 $layer=LI1_cond $X=2.982 $Y=0.73 $X2=2.982
+ $Y2=0.66
r23 7 8 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=2.845 $Y=0.73 $X2=2.175
+ $Y2=0.73
r24 2 15 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.96 $Y2=0.66
r25 1 10 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.06 $Y2=0.66
.ends


* File: sky130_fd_sc_hd__maj3_4.pxi.spice
* Created: Thu Aug 27 14:27:21 2020
* 
x_PM_SKY130_FD_SC_HD__MAJ3_4%C N_C_M1002_g N_C_M1011_g N_C_M1016_g N_C_M1001_g
+ N_C_c_83_n N_C_c_94_n N_C_c_100_p N_C_c_122_p N_C_c_110_p N_C_c_172_p
+ N_C_c_84_n N_C_c_85_n N_C_c_86_n N_C_c_87_n C N_C_c_88_n N_C_c_89_n N_C_c_90_n
+ N_C_c_91_n C PM_SKY130_FD_SC_HD__MAJ3_4%C
x_PM_SKY130_FD_SC_HD__MAJ3_4%A N_A_c_188_n N_A_M1013_g N_A_M1017_g N_A_c_189_n
+ N_A_M1012_g N_A_M1008_g A A N_A_c_198_n N_A_c_190_n
+ PM_SKY130_FD_SC_HD__MAJ3_4%A
x_PM_SKY130_FD_SC_HD__MAJ3_4%B N_B_c_231_n N_B_M1015_g N_B_M1004_g N_B_c_232_n
+ N_B_M1014_g N_B_M1019_g B N_B_c_233_n PM_SKY130_FD_SC_HD__MAJ3_4%B
x_PM_SKY130_FD_SC_HD__MAJ3_4%A_47_297# N_A_47_297#_M1002_s N_A_47_297#_M1015_d
+ N_A_47_297#_M1011_s N_A_47_297#_M1004_d N_A_47_297#_c_271_n
+ N_A_47_297#_M1003_g N_A_47_297#_M1000_g N_A_47_297#_c_272_n
+ N_A_47_297#_M1005_g N_A_47_297#_M1006_g N_A_47_297#_c_273_n
+ N_A_47_297#_M1007_g N_A_47_297#_M1009_g N_A_47_297#_c_274_n
+ N_A_47_297#_M1018_g N_A_47_297#_M1010_g N_A_47_297#_c_285_n
+ N_A_47_297#_c_294_n N_A_47_297#_c_275_n N_A_47_297#_c_301_n
+ N_A_47_297#_c_302_n N_A_47_297#_c_276_n N_A_47_297#_c_277_n
+ N_A_47_297#_c_369_p N_A_47_297#_c_278_n N_A_47_297#_c_287_n
+ N_A_47_297#_c_279_n N_A_47_297#_c_323_n N_A_47_297#_c_280_n
+ PM_SKY130_FD_SC_HD__MAJ3_4%A_47_297#
x_PM_SKY130_FD_SC_HD__MAJ3_4%VPWR N_VPWR_M1017_d N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1010_d N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n
+ N_VPWR_c_448_n N_VPWR_c_449_n VPWR N_VPWR_c_450_n N_VPWR_c_451_n
+ N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_443_n
+ VPWR PM_SKY130_FD_SC_HD__MAJ3_4%VPWR
x_PM_SKY130_FD_SC_HD__MAJ3_4%X N_X_M1003_s N_X_M1007_s N_X_M1000_s N_X_M1009_s
+ N_X_c_535_n N_X_c_543_n N_X_c_531_n N_X_c_532_n N_X_c_536_n N_X_c_558_n
+ N_X_c_561_n N_X_c_564_n X X X N_X_c_534_n N_X_c_538_n
+ PM_SKY130_FD_SC_HD__MAJ3_4%X
x_PM_SKY130_FD_SC_HD__MAJ3_4%VGND N_VGND_M1013_d N_VGND_M1016_d N_VGND_M1005_d
+ N_VGND_M1018_d N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n
+ N_VGND_c_609_n N_VGND_c_610_n VGND N_VGND_c_611_n N_VGND_c_612_n
+ N_VGND_c_613_n N_VGND_c_614_n N_VGND_c_615_n N_VGND_c_616_n N_VGND_c_617_n
+ VGND PM_SKY130_FD_SC_HD__MAJ3_4%VGND
cc_1 VNB N_C_c_83_n 0.00255713f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.285
cc_2 VNB N_C_c_84_n 3.40629e-19 $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=2.225
cc_3 VNB N_C_c_85_n 0.00254731f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.16
cc_4 VNB N_C_c_86_n 0.00110173f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=1.16
cc_5 VNB N_C_c_87_n 0.023781f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=1.16
cc_6 VNB N_C_c_88_n 0.0276542f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_7 VNB N_C_c_89_n 0.0206149f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=0.995
cc_8 VNB N_C_c_90_n 0.017509f $X=-0.19 $Y=-0.24 $X2=2.782 $Y2=0.995
cc_9 VNB N_C_c_91_n 0.00194057f $X=-0.19 $Y=-0.24 $X2=0.72 $Y2=1.18
cc_10 VNB N_A_c_188_n 0.0157238f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_11 VNB N_A_c_189_n 0.0159353f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=0.995
cc_12 VNB N_A_c_190_n 0.0324824f $X=-0.19 $Y=-0.24 $X2=2.545 $Y2=2.225
cc_13 VNB N_B_c_231_n 0.0161625f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.995
cc_14 VNB N_B_c_232_n 0.015595f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=0.995
cc_15 VNB N_B_c_233_n 0.032028f $X=-0.19 $Y=-0.24 $X2=1.79 $Y2=2.31
cc_16 VNB N_A_47_297#_c_271_n 0.0172678f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=1.985
cc_17 VNB N_A_47_297#_c_272_n 0.0157937f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=2.225
cc_18 VNB N_A_47_297#_c_273_n 0.0157835f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=1.16
cc_19 VNB N_A_47_297#_c_274_n 0.0191475f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_20 VNB N_A_47_297#_c_275_n 0.007427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_47_297#_c_276_n 0.00196953f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_47_297#_c_277_n 0.00516934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_47_297#_c_278_n 0.0353894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_47_297#_c_279_n 0.0200405f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_47_297#_c_280_n 0.0649906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_443_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_531_n 0.00188062f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=2
cc_28 VNB N_X_c_532_n 0.00218282f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=2.085
cc_29 VNB X 0.0210201f $X=-0.19 $Y=-0.24 $X2=2.782 $Y2=0.995
cc_30 VNB N_X_c_534_n 0.0123721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_605_n 4.89148e-19 $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.285
cc_32 VNB N_VGND_c_606_n 0.00514051f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=2.085
cc_33 VNB N_VGND_c_607_n 0.0169962f $X=-0.19 $Y=-0.24 $X2=2.46 $Y2=2.31
cc_34 VNB N_VGND_c_608_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=2.63 $Y2=1.16
cc_35 VNB N_VGND_c_609_n 0.0106809f $X=-0.19 $Y=-0.24 $X2=2.78 $Y2=1.16
cc_36 VNB N_VGND_c_610_n 0.00416524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_611_n 0.0293937f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_38 VNB N_VGND_c_612_n 0.0361197f $X=-0.19 $Y=-0.24 $X2=2.782 $Y2=1.16
cc_39 VNB N_VGND_c_613_n 0.0166611f $X=-0.19 $Y=-0.24 $X2=0.805 $Y2=1.18
cc_40 VNB N_VGND_c_614_n 0.00436303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_615_n 0.00660408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_616_n 0.00323604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_617_n 0.258201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_C_M1011_g 0.0225842f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.985
cc_45 VPB N_C_M1001_g 0.0195084f $X=-0.19 $Y=1.305 $X2=2.695 $Y2=1.985
cc_46 VPB N_C_c_94_n 0.00105639f $X=-0.19 $Y=1.305 $X2=0.805 $Y2=1.915
cc_47 VPB N_C_c_84_n 0.00161927f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=2.225
cc_48 VPB N_C_c_87_n 0.00751915f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=1.16
cc_49 VPB N_C_c_88_n 0.00953913f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_50 VPB N_A_M1017_g 0.0175904f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.985
cc_51 VPB N_A_M1008_g 0.0178759f $X=-0.19 $Y=1.305 $X2=2.695 $Y2=1.985
cc_52 VPB N_A_c_190_n 0.00451192f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=2.225
cc_53 VPB N_B_M1004_g 0.0187785f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.985
cc_54 VPB N_B_M1019_g 0.0180762f $X=-0.19 $Y=1.305 $X2=2.695 $Y2=1.985
cc_55 VPB N_B_c_233_n 0.004171f $X=-0.19 $Y=1.305 $X2=1.79 $Y2=2.31
cc_56 VPB N_A_47_297#_M1000_g 0.0207373f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=2
cc_57 VPB N_A_47_297#_M1006_g 0.0182176f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.16
cc_58 VPB N_A_47_297#_M1009_g 0.0181992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_47_297#_M1010_g 0.0218907f $X=-0.19 $Y=1.305 $X2=2.782 $Y2=0.995
cc_60 VPB N_A_47_297#_c_285_n 0.0366532f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.19
cc_61 VPB N_A_47_297#_c_275_n 0.00312718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_47_297#_c_287_n 0.0111995f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_47_297#_c_279_n 0.00724139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_47_297#_c_280_n 0.0103056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_444_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0.805 $Y2=1.285
cc_66 VPB N_VPWR_c_445_n 0.0102498f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=2.085
cc_67 VPB N_VPWR_c_446_n 0.0189004f $X=-0.19 $Y=1.305 $X2=2.545 $Y2=1.245
cc_68 VPB N_VPWR_c_447_n 0.00410835f $X=-0.19 $Y=1.305 $X2=2.78 $Y2=1.16
cc_69 VPB N_VPWR_c_448_n 0.0105174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_449_n 0.00438892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_450_n 0.0313984f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_72 VPB N_VPWR_c_451_n 0.0342412f $X=-0.19 $Y=1.305 $X2=2.782 $Y2=1.325
cc_73 VPB N_VPWR_c_452_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_453_n 0.00436154f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_454_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_455_n 0.00323736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_443_n 0.0461355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_X_c_535_n 0.0022339f $X=-0.19 $Y=1.305 $X2=2.695 $Y2=1.985
cc_79 VPB N_X_c_536_n 0.00218546f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=2.31
cc_80 VPB X 0.00831516f $X=-0.19 $Y=1.305 $X2=2.782 $Y2=0.995
cc_81 VPB N_X_c_538_n 0.0125274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 N_C_c_89_n N_A_c_188_n 0.0435952f $X=0.59 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_83 N_C_M1011_g N_A_M1017_g 0.0435952f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_84 N_C_c_100_p N_A_M1017_g 0.0134418f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_85 N_C_c_100_p N_A_M1008_g 0.0147922f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_86 N_C_c_83_n N_A_c_198_n 0.0173748f $X=0.805 $Y=1.285 $X2=0 $Y2=0
cc_87 N_C_c_94_n N_A_c_198_n 0.0263696f $X=0.805 $Y=1.915 $X2=0 $Y2=0
cc_88 N_C_c_100_p N_A_c_198_n 0.0145635f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_89 N_C_c_88_n N_A_c_198_n 5.0881e-19 $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_90 N_C_c_83_n N_A_c_190_n 0.00160717f $X=0.805 $Y=1.285 $X2=0 $Y2=0
cc_91 N_C_c_94_n N_A_c_190_n 0.00817523f $X=0.805 $Y=1.915 $X2=0 $Y2=0
cc_92 N_C_c_100_p N_A_c_190_n 3.22614e-19 $X=1.62 $Y=2 $X2=0 $Y2=0
cc_93 N_C_c_88_n N_A_c_190_n 0.0435952f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_94 N_C_c_110_p N_B_M1004_g 0.0108531f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_95 N_C_c_90_n N_B_c_232_n 0.0518917f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_96 N_C_M1001_g N_B_M1019_g 0.0518917f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_97 N_C_c_110_p N_B_M1019_g 0.0132508f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_98 N_C_c_84_n B 0.00592804f $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_99 N_C_c_85_n B 0.0139301f $X=2.63 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C_c_84_n N_B_c_233_n 0.00495375f $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_101 N_C_c_85_n N_B_c_233_n 0.0013712f $X=2.63 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C_c_87_n N_B_c_233_n 0.0518917f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_103 N_C_c_110_p N_A_47_297#_M1004_d 0.00335253f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_104 N_C_c_90_n N_A_47_297#_c_271_n 0.0181763f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C_M1001_g N_A_47_297#_M1000_g 0.0224466f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_106 N_C_c_122_p N_A_47_297#_c_285_n 0.0103497f $X=0.89 $Y=2 $X2=0 $Y2=0
cc_107 N_C_c_83_n N_A_47_297#_c_294_n 0.0110378f $X=0.805 $Y=1.285 $X2=0 $Y2=0
cc_108 N_C_c_89_n N_A_47_297#_c_294_n 0.0101286f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_109 N_C_c_91_n N_A_47_297#_c_294_n 0.00544125f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_110 N_C_M1001_g N_A_47_297#_c_275_n 3.96997e-19 $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_111 N_C_c_100_p N_A_47_297#_c_275_n 0.0137112f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_112 N_C_c_110_p N_A_47_297#_c_275_n 0.019506f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_113 N_C_c_84_n N_A_47_297#_c_275_n 0.00452226f $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_114 N_C_c_90_n N_A_47_297#_c_301_n 0.00142909f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C_c_85_n N_A_47_297#_c_302_n 0.0108187f $X=2.63 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_c_86_n N_A_47_297#_c_302_n 0.0180199f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_117 N_C_c_87_n N_A_47_297#_c_302_n 0.00410162f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_118 N_C_c_90_n N_A_47_297#_c_302_n 0.0127166f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C_c_87_n N_A_47_297#_c_276_n 0.00171871f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_c_90_n N_A_47_297#_c_276_n 0.00199392f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_121 N_C_c_84_n N_A_47_297#_c_277_n 0.00145926f $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_122 N_C_c_86_n N_A_47_297#_c_277_n 0.0146215f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_123 N_C_c_87_n N_A_47_297#_c_277_n 0.00119787f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C_c_88_n N_A_47_297#_c_278_n 0.00434498f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_125 N_C_c_89_n N_A_47_297#_c_278_n 0.00915574f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_126 N_C_c_91_n N_A_47_297#_c_278_n 0.0128103f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_127 N_C_M1011_g N_A_47_297#_c_287_n 0.0257076f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_128 N_C_c_94_n N_A_47_297#_c_287_n 0.0252423f $X=0.805 $Y=1.915 $X2=0 $Y2=0
cc_129 N_C_c_88_n N_A_47_297#_c_287_n 9.5351e-19 $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_130 N_C_c_91_n N_A_47_297#_c_287_n 0.00319035f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_131 N_C_M1011_g N_A_47_297#_c_279_n 0.00140958f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_132 N_C_c_94_n N_A_47_297#_c_279_n 0.00401274f $X=0.805 $Y=1.915 $X2=0 $Y2=0
cc_133 N_C_c_88_n N_A_47_297#_c_279_n 0.00556899f $X=0.59 $Y=1.16 $X2=0 $Y2=0
cc_134 N_C_c_89_n N_A_47_297#_c_279_n 0.00168233f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_135 N_C_c_91_n N_A_47_297#_c_279_n 0.0161301f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_136 N_C_c_90_n N_A_47_297#_c_323_n 2.70861e-19 $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C_c_84_n N_A_47_297#_c_280_n 9.17807e-19 $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_138 N_C_c_87_n N_A_47_297#_c_280_n 0.0133549f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_139 N_C_c_94_n A_151_297# 0.00436024f $X=0.805 $Y=1.915 $X2=-0.19 $Y2=-0.24
cc_140 N_C_c_100_p A_151_297# 0.00289102f $X=1.62 $Y=2 $X2=-0.19 $Y2=-0.24
cc_141 N_C_c_122_p A_151_297# 0.00140764f $X=0.89 $Y=2 $X2=-0.19 $Y2=-0.24
cc_142 N_C_c_100_p N_VPWR_M1017_d 0.00355609f $X=1.62 $Y=2 $X2=-0.19 $Y2=-0.24
cc_143 N_C_M1011_g N_VPWR_c_444_n 0.00182394f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_144 N_C_c_100_p N_VPWR_c_444_n 0.0159625f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_145 N_C_M1001_g N_VPWR_c_445_n 0.0152069f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_146 N_C_c_110_p N_VPWR_c_445_n 0.0116785f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_147 N_C_c_84_n N_VPWR_c_445_n 0.0475996f $X=2.545 $Y=2.225 $X2=0 $Y2=0
cc_148 N_C_c_86_n N_VPWR_c_445_n 0.00682027f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_149 N_C_c_87_n N_VPWR_c_445_n 0.00249055f $X=2.78 $Y=1.16 $X2=0 $Y2=0
cc_150 N_C_M1011_g N_VPWR_c_450_n 0.00547949f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_151 N_C_c_100_p N_VPWR_c_450_n 0.00343154f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_152 N_C_c_122_p N_VPWR_c_450_n 0.00267754f $X=0.89 $Y=2 $X2=0 $Y2=0
cc_153 N_C_M1001_g N_VPWR_c_451_n 0.00571152f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_154 N_C_c_100_p N_VPWR_c_451_n 0.00244309f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_155 N_C_c_110_p N_VPWR_c_451_n 0.0316032f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_156 N_C_c_172_p N_VPWR_c_451_n 0.00771938f $X=1.79 $Y=2.31 $X2=0 $Y2=0
cc_157 N_C_M1011_g N_VPWR_c_443_n 0.0107683f $X=0.68 $Y=1.985 $X2=0 $Y2=0
cc_158 N_C_M1001_g N_VPWR_c_443_n 0.0107347f $X=2.695 $Y=1.985 $X2=0 $Y2=0
cc_159 N_C_c_100_p N_VPWR_c_443_n 0.0116255f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_160 N_C_c_122_p N_VPWR_c_443_n 0.00492202f $X=0.89 $Y=2 $X2=0 $Y2=0
cc_161 N_C_c_110_p N_VPWR_c_443_n 0.0287047f $X=2.46 $Y=2.31 $X2=0 $Y2=0
cc_162 N_C_c_172_p N_VPWR_c_443_n 0.00623193f $X=1.79 $Y=2.31 $X2=0 $Y2=0
cc_163 N_C_c_100_p A_314_297# 0.00190901f $X=1.62 $Y=2 $X2=-0.19 $Y2=-0.24
cc_164 N_C_c_172_p A_314_297# 0.00197209f $X=1.79 $Y=2.31 $X2=-0.19 $Y2=-0.24
cc_165 N_C_c_110_p A_482_297# 0.00108703f $X=2.46 $Y=2.31 $X2=-0.19 $Y2=-0.24
cc_166 N_C_c_89_n N_VGND_c_605_n 0.0018479f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_167 N_C_c_90_n N_VGND_c_606_n 0.00775599f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_168 N_C_c_89_n N_VGND_c_611_n 0.00416048f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C_c_90_n N_VGND_c_612_n 0.00436487f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C_c_89_n N_VGND_c_617_n 0.00682124f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_171 N_C_c_90_n N_VGND_c_617_n 0.00640166f $X=2.782 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_189_n N_B_c_231_n 0.0367288f $X=1.495 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_173 N_A_M1008_g N_B_M1004_g 0.0367288f $X=1.495 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A_c_190_n N_B_c_233_n 0.0367288f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_c_188_n N_A_47_297#_c_294_n 0.0153627f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_189_n N_A_47_297#_c_294_n 0.0174342f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_198_n N_A_47_297#_c_294_n 0.0238047f $X=1.285 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_190_n N_A_47_297#_c_294_n 0.00220502f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_189_n N_A_47_297#_c_275_n 0.00807776f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_M1008_g N_A_47_297#_c_275_n 9.48716e-19 $X=1.495 $Y=1.985 $X2=0 $Y2=0
cc_181 N_A_c_198_n N_A_47_297#_c_275_n 0.0334418f $X=1.285 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_189_n N_A_47_297#_c_301_n 0.00153014f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_c_188_n N_A_47_297#_c_278_n 0.00161843f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_198_n N_VPWR_M1017_d 0.00216303f $X=1.285 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_185 N_A_M1017_g N_VPWR_c_444_n 0.00973976f $X=1.075 $Y=1.985 $X2=0 $Y2=0
cc_186 N_A_M1008_g N_VPWR_c_444_n 0.00840395f $X=1.495 $Y=1.985 $X2=0 $Y2=0
cc_187 N_A_M1017_g N_VPWR_c_450_n 0.00339367f $X=1.075 $Y=1.985 $X2=0 $Y2=0
cc_188 N_A_M1008_g N_VPWR_c_451_n 0.00339367f $X=1.495 $Y=1.985 $X2=0 $Y2=0
cc_189 N_A_M1017_g N_VPWR_c_443_n 0.0039496f $X=1.075 $Y=1.985 $X2=0 $Y2=0
cc_190 N_A_M1008_g N_VPWR_c_443_n 0.00401529f $X=1.495 $Y=1.985 $X2=0 $Y2=0
cc_191 N_A_c_188_n N_VGND_c_605_n 0.00961653f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_189_n N_VGND_c_605_n 0.00975027f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_188_n N_VGND_c_611_n 0.00342263f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_189_n N_VGND_c_612_n 0.00342263f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_188_n N_VGND_c_617_n 0.00399861f $X=1.075 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_189_n N_VGND_c_617_n 0.0040643f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B_c_231_n N_A_47_297#_c_275_n 0.00905542f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B_M1004_g N_A_47_297#_c_275_n 0.016362f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_199 N_B_M1019_g N_A_47_297#_c_275_n 0.0061734f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_200 B N_A_47_297#_c_275_n 0.0358593f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_201 N_B_c_233_n N_A_47_297#_c_275_n 0.00201841f $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B_c_231_n N_A_47_297#_c_301_n 0.0075627f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B_c_232_n N_A_47_297#_c_301_n 0.00759048f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_204 N_B_c_232_n N_A_47_297#_c_302_n 0.0116364f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B_c_231_n N_A_47_297#_c_323_n 0.0124771f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B_c_232_n N_A_47_297#_c_323_n 0.00208195f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_207 B N_A_47_297#_c_323_n 0.0181722f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_208 N_B_c_233_n N_A_47_297#_c_323_n 0.00220628f $X=2.335 $Y=1.16 $X2=0 $Y2=0
cc_209 N_B_M1004_g N_VPWR_c_444_n 0.00159208f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_210 N_B_M1004_g N_VPWR_c_451_n 0.0037209f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_211 N_B_M1019_g N_VPWR_c_451_n 0.0037209f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_212 N_B_M1004_g N_VPWR_c_443_n 0.00532914f $X=1.915 $Y=1.985 $X2=0 $Y2=0
cc_213 N_B_M1019_g N_VPWR_c_443_n 0.00516633f $X=2.335 $Y=1.985 $X2=0 $Y2=0
cc_214 N_B_c_231_n N_VGND_c_605_n 0.00182905f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_231_n N_VGND_c_612_n 0.00415003f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B_c_232_n N_VGND_c_612_n 0.00421197f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_231_n N_VGND_c_617_n 0.00579681f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_232_n N_VGND_c_617_n 0.00572905f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_47_297#_c_285_n N_VPWR_c_444_n 0.00564305f $X=0.38 $Y=2.3 $X2=0 $Y2=0
cc_220 N_A_47_297#_M1000_g N_VPWR_c_445_n 0.0135283f $X=3.33 $Y=1.985 $X2=0
+ $Y2=0
cc_221 N_A_47_297#_c_302_n N_VPWR_c_445_n 0.00590988f $X=3.115 $Y=0.8 $X2=0
+ $Y2=0
cc_222 N_A_47_297#_c_277_n N_VPWR_c_445_n 0.00545579f $X=3.285 $Y=1.18 $X2=0
+ $Y2=0
cc_223 N_A_47_297#_M1000_g N_VPWR_c_446_n 0.00541359f $X=3.33 $Y=1.985 $X2=0
+ $Y2=0
cc_224 N_A_47_297#_M1006_g N_VPWR_c_446_n 0.00541359f $X=3.75 $Y=1.985 $X2=0
+ $Y2=0
cc_225 N_A_47_297#_M1006_g N_VPWR_c_447_n 0.00268723f $X=3.75 $Y=1.985 $X2=0
+ $Y2=0
cc_226 N_A_47_297#_M1009_g N_VPWR_c_447_n 0.00146448f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_227 N_A_47_297#_M1010_g N_VPWR_c_449_n 0.0031902f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_228 N_A_47_297#_c_285_n N_VPWR_c_450_n 0.026786f $X=0.38 $Y=2.3 $X2=0 $Y2=0
cc_229 N_A_47_297#_M1009_g N_VPWR_c_452_n 0.00541359f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_230 N_A_47_297#_M1010_g N_VPWR_c_452_n 0.00541359f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_231 N_A_47_297#_M1011_s N_VPWR_c_443_n 0.00789791f $X=0.235 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_47_297#_M1004_d N_VPWR_c_443_n 0.00222735f $X=1.99 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_47_297#_M1000_g N_VPWR_c_443_n 0.0101378f $X=3.33 $Y=1.985 $X2=0
+ $Y2=0
cc_234 N_A_47_297#_M1006_g N_VPWR_c_443_n 0.00950154f $X=3.75 $Y=1.985 $X2=0
+ $Y2=0
cc_235 N_A_47_297#_M1009_g N_VPWR_c_443_n 0.00950154f $X=4.17 $Y=1.985 $X2=0
+ $Y2=0
cc_236 N_A_47_297#_M1010_g N_VPWR_c_443_n 0.0104557f $X=4.59 $Y=1.985 $X2=0
+ $Y2=0
cc_237 N_A_47_297#_c_285_n N_VPWR_c_443_n 0.0145574f $X=0.38 $Y=2.3 $X2=0 $Y2=0
cc_238 N_A_47_297#_c_275_n A_314_297# 0.00205406f $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_239 N_A_47_297#_M1000_g N_X_c_535_n 0.0027286f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_47_297#_M1006_g N_X_c_535_n 0.00123753f $X=3.75 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_47_297#_c_369_p N_X_c_535_n 0.0267295f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_47_297#_c_280_n N_X_c_535_n 0.00220041f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_47_297#_M1000_g N_X_c_543_n 0.00985325f $X=3.33 $Y=1.985 $X2=0 $Y2=0
cc_244 N_A_47_297#_M1006_g N_X_c_543_n 0.0101686f $X=3.75 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_47_297#_M1009_g N_X_c_543_n 6.31279e-19 $X=4.17 $Y=1.985 $X2=0 $Y2=0
cc_246 N_A_47_297#_c_272_n N_X_c_531_n 0.00461054f $X=3.75 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_47_297#_c_276_n N_X_c_531_n 0.00153275f $X=3.2 $Y=1.075 $X2=0 $Y2=0
cc_248 N_A_47_297#_c_369_p N_X_c_531_n 0.0202409f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_47_297#_c_280_n N_X_c_531_n 0.00230339f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_47_297#_c_272_n N_X_c_532_n 0.00890471f $X=3.75 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_47_297#_c_273_n N_X_c_532_n 0.0088553f $X=4.17 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_47_297#_c_369_p N_X_c_532_n 0.0603554f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_47_297#_c_280_n N_X_c_532_n 0.00222429f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_47_297#_M1006_g N_X_c_536_n 0.0107189f $X=3.75 $Y=1.985 $X2=0 $Y2=0
cc_255 N_A_47_297#_M1009_g N_X_c_536_n 0.0107189f $X=4.17 $Y=1.985 $X2=0 $Y2=0
cc_256 N_A_47_297#_c_369_p N_X_c_536_n 0.0598351f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_47_297#_c_280_n N_X_c_536_n 0.00211509f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_47_297#_c_272_n N_X_c_558_n 5.2007e-19 $X=3.75 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_47_297#_c_273_n N_X_c_558_n 0.00631111f $X=4.17 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_47_297#_c_274_n N_X_c_558_n 0.0109535f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_47_297#_M1006_g N_X_c_561_n 6.32068e-19 $X=3.75 $Y=1.985 $X2=0 $Y2=0
cc_262 N_A_47_297#_M1009_g N_X_c_561_n 0.0102742f $X=4.17 $Y=1.985 $X2=0 $Y2=0
cc_263 N_A_47_297#_M1010_g N_X_c_561_n 0.0151316f $X=4.59 $Y=1.985 $X2=0 $Y2=0
cc_264 N_A_47_297#_c_271_n N_X_c_564_n 0.00352607f $X=3.33 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_47_297#_c_272_n N_X_c_564_n 0.00269075f $X=3.75 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_47_297#_c_273_n N_X_c_564_n 5.20035e-19 $X=4.17 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_47_297#_c_369_p N_X_c_564_n 0.00135981f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_47_297#_c_274_n X 0.0213848f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_47_297#_c_369_p X 0.0171439f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_47_297#_c_273_n N_X_c_534_n 0.0012996f $X=4.17 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_47_297#_c_274_n N_X_c_534_n 0.0133172f $X=4.59 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_47_297#_c_280_n N_X_c_534_n 0.00222429f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_47_297#_M1009_g N_X_c_538_n 0.00128444f $X=4.17 $Y=1.985 $X2=0 $Y2=0
cc_274 N_A_47_297#_M1010_g N_X_c_538_n 0.0149864f $X=4.59 $Y=1.985 $X2=0 $Y2=0
cc_275 N_A_47_297#_c_280_n N_X_c_538_n 0.00211509f $X=4.59 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_47_297#_c_294_n A_151_47# 0.00534239f $X=1.62 $Y=0.772 $X2=-0.19
+ $Y2=-0.24
cc_277 N_A_47_297#_c_294_n N_VGND_M1013_d 0.00313547f $X=1.62 $Y=0.772 $X2=-0.19
+ $Y2=-0.24
cc_278 N_A_47_297#_c_302_n N_VGND_M1016_d 0.00958334f $X=3.115 $Y=0.8 $X2=0
+ $Y2=0
cc_279 N_A_47_297#_c_294_n N_VGND_c_605_n 0.0163859f $X=1.62 $Y=0.772 $X2=0
+ $Y2=0
cc_280 N_A_47_297#_c_301_n N_VGND_c_605_n 0.00718914f $X=2.125 $Y=0.38 $X2=0
+ $Y2=0
cc_281 N_A_47_297#_c_278_n N_VGND_c_605_n 0.00781685f $X=0.47 $Y=0.38 $X2=0
+ $Y2=0
cc_282 N_A_47_297#_c_271_n N_VGND_c_606_n 0.00394292f $X=3.33 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_47_297#_c_301_n N_VGND_c_606_n 0.008733f $X=2.125 $Y=0.38 $X2=0 $Y2=0
cc_284 N_A_47_297#_c_302_n N_VGND_c_606_n 0.0268661f $X=3.115 $Y=0.8 $X2=0 $Y2=0
cc_285 N_A_47_297#_c_271_n N_VGND_c_607_n 0.00511552f $X=3.33 $Y=0.995 $X2=0
+ $Y2=0
cc_286 N_A_47_297#_c_272_n N_VGND_c_607_n 0.00422241f $X=3.75 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_47_297#_c_302_n N_VGND_c_607_n 8.37243e-19 $X=3.115 $Y=0.8 $X2=0
+ $Y2=0
cc_288 N_A_47_297#_c_272_n N_VGND_c_608_n 0.00146448f $X=3.75 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_47_297#_c_273_n N_VGND_c_608_n 0.00146448f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_47_297#_c_274_n N_VGND_c_610_n 0.00316354f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_47_297#_c_294_n N_VGND_c_611_n 0.0070234f $X=1.62 $Y=0.772 $X2=0
+ $Y2=0
cc_292 N_A_47_297#_c_278_n N_VGND_c_611_n 0.0366566f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_293 N_A_47_297#_c_294_n N_VGND_c_612_n 0.00747719f $X=1.62 $Y=0.772 $X2=0
+ $Y2=0
cc_294 N_A_47_297#_c_301_n N_VGND_c_612_n 0.018363f $X=2.125 $Y=0.38 $X2=0 $Y2=0
cc_295 N_A_47_297#_c_302_n N_VGND_c_612_n 0.00694641f $X=3.115 $Y=0.8 $X2=0
+ $Y2=0
cc_296 N_A_47_297#_c_273_n N_VGND_c_613_n 0.00421248f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_47_297#_c_274_n N_VGND_c_613_n 0.00421248f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_47_297#_M1002_s N_VGND_c_617_n 0.00225715f $X=0.325 $Y=0.235 $X2=0
+ $Y2=0
cc_299 N_A_47_297#_M1015_d N_VGND_c_617_n 0.00215201f $X=1.99 $Y=0.235 $X2=0
+ $Y2=0
cc_300 N_A_47_297#_c_271_n N_VGND_c_617_n 0.00911441f $X=3.33 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_47_297#_c_272_n N_VGND_c_617_n 0.00569656f $X=3.75 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_47_297#_c_273_n N_VGND_c_617_n 0.00571103f $X=4.17 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_47_297#_c_274_n N_VGND_c_617_n 0.00666524f $X=4.59 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_47_297#_c_294_n N_VGND_c_617_n 0.0270673f $X=1.62 $Y=0.772 $X2=0
+ $Y2=0
cc_305 N_A_47_297#_c_301_n N_VGND_c_617_n 0.0120598f $X=2.125 $Y=0.38 $X2=0
+ $Y2=0
cc_306 N_A_47_297#_c_302_n N_VGND_c_617_n 0.0173286f $X=3.115 $Y=0.8 $X2=0 $Y2=0
cc_307 N_A_47_297#_c_278_n N_VGND_c_617_n 0.0208703f $X=0.47 $Y=0.38 $X2=0 $Y2=0
cc_308 N_A_47_297#_c_275_n A_314_47# 4.61277e-19 $X=1.705 $Y=1.545 $X2=-0.19
+ $Y2=-0.24
cc_309 N_A_47_297#_c_323_n A_314_47# 0.00328779f $X=2.29 $Y=0.772 $X2=-0.19
+ $Y2=-0.24
cc_310 N_A_47_297#_c_302_n A_482_47# 0.00289474f $X=3.115 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_311 A_151_297# N_VPWR_c_443_n 0.00285919f $X=0.755 $Y=1.485 $X2=0 $Y2=0
cc_312 N_VPWR_c_443_n A_314_297# 0.00239791f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_313 N_VPWR_c_443_n A_482_297# 0.00173156f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_314 N_VPWR_c_443_n N_X_M1000_s 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_443_n N_X_M1009_s 0.00215201f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_c_445_n N_X_c_535_n 0.0123957f $X=3.01 $Y=1.62 $X2=0 $Y2=0
cc_317 N_VPWR_c_445_n N_X_c_543_n 0.0575032f $X=3.01 $Y=1.62 $X2=0 $Y2=0
cc_318 N_VPWR_c_446_n N_X_c_543_n 0.0189039f $X=3.875 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_443_n N_X_c_543_n 0.0122217f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_M1006_d N_X_c_536_n 0.00165831f $X=3.825 $Y=1.485 $X2=0 $Y2=0
cc_321 N_VPWR_c_447_n N_X_c_536_n 0.0126919f $X=3.96 $Y=1.96 $X2=0 $Y2=0
cc_322 N_VPWR_c_452_n N_X_c_561_n 0.0189039f $X=4.715 $Y=2.72 $X2=0 $Y2=0
cc_323 N_VPWR_c_443_n N_X_c_561_n 0.0122217f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_M1010_d N_X_c_538_n 0.00276279f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_325 N_VPWR_c_449_n N_X_c_538_n 0.0164344f $X=4.8 $Y=1.96 $X2=0 $Y2=0
cc_326 N_X_c_532_n N_VGND_M1005_d 0.00162148f $X=4.215 $Y=0.81 $X2=0 $Y2=0
cc_327 N_X_c_534_n N_VGND_M1018_d 0.00319503f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_328 N_X_c_532_n N_VGND_c_607_n 0.00203746f $X=4.215 $Y=0.81 $X2=0 $Y2=0
cc_329 N_X_c_564_n N_VGND_c_607_n 0.0187247f $X=3.54 $Y=0.4 $X2=0 $Y2=0
cc_330 N_X_c_532_n N_VGND_c_608_n 0.0122675f $X=4.215 $Y=0.81 $X2=0 $Y2=0
cc_331 N_X_c_534_n N_VGND_c_609_n 0.00138263f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_332 N_X_c_534_n N_VGND_c_610_n 0.0127393f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_333 N_X_c_532_n N_VGND_c_613_n 0.0041083f $X=4.215 $Y=0.81 $X2=0 $Y2=0
cc_334 N_X_c_558_n N_VGND_c_613_n 0.0184921f $X=4.38 $Y=0.4 $X2=0 $Y2=0
cc_335 N_X_M1003_s N_VGND_c_617_n 0.00215201f $X=3.405 $Y=0.235 $X2=0 $Y2=0
cc_336 N_X_M1007_s N_VGND_c_617_n 0.00215201f $X=4.245 $Y=0.235 $X2=0 $Y2=0
cc_337 N_X_c_532_n N_VGND_c_617_n 0.0124122f $X=4.215 $Y=0.81 $X2=0 $Y2=0
cc_338 N_X_c_558_n N_VGND_c_617_n 0.012098f $X=4.38 $Y=0.4 $X2=0 $Y2=0
cc_339 N_X_c_564_n N_VGND_c_617_n 0.0121358f $X=3.54 $Y=0.4 $X2=0 $Y2=0
cc_340 N_X_c_534_n N_VGND_c_617_n 0.00310154f $X=4.845 $Y=0.905 $X2=0 $Y2=0
cc_341 A_151_47# N_VGND_c_617_n 0.00295002f $X=0.755 $Y=0.235 $X2=3.54 $Y2=1.16
cc_342 N_VGND_c_617_n A_314_47# 0.00325105f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_343 N_VGND_c_617_n A_482_47# 0.00269901f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24

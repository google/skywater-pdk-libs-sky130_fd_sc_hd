* File: sky130_fd_sc_hd__or4_1.spice.SKY130_FD_SC_HD__OR4_1.pxi
* Created: Thu Aug 27 14:43:59 2020
* 
x_PM_SKY130_FD_SC_HD__OR4_1%D N_D_M1005_g N_D_M1008_g D D N_D_c_62_n
+ PM_SKY130_FD_SC_HD__OR4_1%D
x_PM_SKY130_FD_SC_HD__OR4_1%C N_C_M1009_g N_C_M1000_g C C N_C_c_90_n
+ PM_SKY130_FD_SC_HD__OR4_1%C
x_PM_SKY130_FD_SC_HD__OR4_1%B N_B_M1002_g N_B_c_126_n N_B_M1004_g B B B
+ N_B_c_128_n N_B_c_129_n PM_SKY130_FD_SC_HD__OR4_1%B
x_PM_SKY130_FD_SC_HD__OR4_1%A N_A_M1003_g N_A_M1007_g A N_A_c_161_n N_A_c_162_n
+ PM_SKY130_FD_SC_HD__OR4_1%A
x_PM_SKY130_FD_SC_HD__OR4_1%A_27_297# N_A_27_297#_M1005_d N_A_27_297#_M1004_d
+ N_A_27_297#_M1008_s N_A_27_297#_M1006_g N_A_27_297#_M1001_g
+ N_A_27_297#_c_211_n N_A_27_297#_c_283_p N_A_27_297#_c_202_n
+ N_A_27_297#_c_203_n N_A_27_297#_c_292_p N_A_27_297#_c_204_n
+ N_A_27_297#_c_238_n N_A_27_297#_c_212_n N_A_27_297#_c_213_n
+ N_A_27_297#_c_205_n N_A_27_297#_c_214_n N_A_27_297#_c_206_n
+ N_A_27_297#_c_207_n N_A_27_297#_c_208_n N_A_27_297#_c_209_n
+ PM_SKY130_FD_SC_HD__OR4_1%A_27_297#
x_PM_SKY130_FD_SC_HD__OR4_1%VPWR N_VPWR_M1007_d N_VPWR_c_308_n VPWR
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_307_n N_VPWR_c_312_n
+ PM_SKY130_FD_SC_HD__OR4_1%VPWR
x_PM_SKY130_FD_SC_HD__OR4_1%X N_X_M1006_d N_X_M1001_d N_X_c_333_n N_X_c_335_n
+ N_X_c_334_n X PM_SKY130_FD_SC_HD__OR4_1%X
x_PM_SKY130_FD_SC_HD__OR4_1%VGND N_VGND_M1005_s N_VGND_M1009_d N_VGND_M1003_d
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n VGND
+ N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n
+ N_VGND_c_360_n PM_SKY130_FD_SC_HD__OR4_1%VGND
cc_1 VNB N_D_M1005_g 0.0343362f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_2 VNB D 0.0236217f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_c_62_n 0.0355361f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_4 VNB N_C_M1009_g 0.0257827f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_5 VNB C 0.00562839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_C_c_90_n 0.0180743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_M1002_g 0.0180611f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_126_n 0.0264562f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_9 VNB N_A_M1003_g 0.0266384f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.475
cc_10 VNB N_A_c_161_n 0.020616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_162_n 0.00317591f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_12 VNB N_A_27_297#_c_202_n 0.00394971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_297#_c_203_n 0.00296979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_297#_c_204_n 0.00109036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_297#_c_205_n 0.00147654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_206_n 0.00185986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_207_n 0.0237064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_208_n 0.00106882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_209_n 0.0197132f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_307_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_333_n 0.0137322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_334_n 0.0241466f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_23 VNB N_VGND_c_351_n 0.0105427f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_VGND_c_352_n 0.0168474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_353_n 8.05577e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_354_n 6.33941e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_355_n 0.014035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_356_n 0.0115649f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_357_n 0.0164993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_358_n 0.168482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_359_n 0.00472891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_360_n 0.0052385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_D_M1008_g 0.0267282f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_34 VPB D 0.00359125f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_35 VPB N_D_c_62_n 0.0095147f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_36 VPB N_C_M1000_g 0.01663f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_37 VPB C 0.0018547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_C_c_90_n 0.00440081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_B_M1002_g 0.0243546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_B_c_128_n 0.0369905f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_41 VPB N_B_c_129_n 0.047246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_M1007_g 0.021674f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_43 VPB N_A_c_161_n 0.00400696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_c_162_n 0.00154474f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_45 VPB N_A_27_297#_M1001_g 0.0244633f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_46 VPB N_A_27_297#_c_211_n 0.00536076f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_47 VPB N_A_27_297#_c_212_n 0.0015591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_297#_c_213_n 0.0209902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_297#_c_214_n 0.00201186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_297#_c_207_n 0.00559796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_308_n 0.0126559f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.695
cc_52 VPB N_VPWR_c_309_n 0.0489859f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_53 VPB N_VPWR_c_310_n 0.0176015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_307_n 0.0614133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_312_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_X_c_335_n 0.0051537f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_57 VPB N_X_c_334_n 0.00879484f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_58 VPB X 0.0321952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 N_D_M1005_g N_C_M1009_g 0.0171645f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_60 D N_C_M1009_g 8.90538e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_61 N_D_M1008_g N_C_M1000_g 0.0254979f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_62 D C 0.0279539f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_63 N_D_c_62_n C 0.00905747f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_64 D N_C_c_90_n 2.65685e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_65 N_D_c_62_n N_C_c_90_n 0.0207331f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_66 N_D_M1008_g N_B_c_129_n 0.00441071f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_67 N_D_M1008_g N_A_27_297#_c_211_n 0.0112539f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_68 D N_A_27_297#_c_211_n 9.67991e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_69 N_D_M1005_g N_A_27_297#_c_203_n 0.00368534f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_70 D N_A_27_297#_c_203_n 0.00556084f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_71 N_D_M1008_g N_A_27_297#_c_213_n 0.00686729f $X=0.47 $Y=1.695 $X2=0 $Y2=0
cc_72 D N_A_27_297#_c_213_n 0.0243507f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_73 N_D_c_62_n N_A_27_297#_c_213_n 0.00190153f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_74 N_D_M1005_g N_VGND_c_352_n 0.0102085f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_75 D N_VGND_c_352_n 0.0260059f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_76 N_D_c_62_n N_VGND_c_352_n 0.00113138f $X=0.47 $Y=1.16 $X2=0 $Y2=0
cc_77 N_D_M1005_g N_VGND_c_353_n 5.21337e-19 $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_78 N_D_M1005_g N_VGND_c_355_n 0.00430458f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_79 N_D_M1005_g N_VGND_c_358_n 0.00749122f $X=0.47 $Y=0.475 $X2=0 $Y2=0
cc_80 D N_VGND_c_358_n 0.00186827f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_81 C N_B_M1002_g 0.0186833f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_82 N_C_c_90_n N_B_M1002_g 0.0411537f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_M1009_g N_B_c_126_n 0.0548441f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_84 N_C_M1000_g N_B_c_129_n 0.00439246f $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_85 C N_A_M1007_g 8.9759e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_86 C N_A_c_161_n 2.88415e-19 $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_87 C N_A_c_162_n 0.0281805f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_88 N_C_M1000_g N_A_27_297#_c_211_n 0.00925462f $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_89 C N_A_27_297#_c_211_n 0.0421076f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_90 N_C_c_90_n N_A_27_297#_c_211_n 3.74254e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_91 N_C_M1009_g N_A_27_297#_c_202_n 0.0110261f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_92 C N_A_27_297#_c_202_n 0.0414766f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_93 N_C_c_90_n N_A_27_297#_c_202_n 0.00179145f $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_94 C N_A_27_297#_c_203_n 0.0152593f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_95 N_C_c_90_n N_A_27_297#_c_203_n 9.23324e-19 $X=0.89 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C_M1000_g N_A_27_297#_c_213_n 9.69529e-19 $X=0.95 $Y=1.695 $X2=0 $Y2=0
cc_97 C N_A_27_297#_c_213_n 0.0086791f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_98 C N_A_27_297#_c_214_n 0.00860775f $X=1.07 $Y=1.105 $X2=0 $Y2=0
cc_99 C A_109_297# 0.00398871f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_100 C A_205_297# 0.00106447f $X=1.07 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_101 N_C_M1009_g N_VGND_c_352_n 5.50577e-19 $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_102 N_C_M1009_g N_VGND_c_353_n 0.00712013f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_103 N_C_M1009_g N_VGND_c_355_n 0.00322006f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_104 N_C_M1009_g N_VGND_c_358_n 0.00401385f $X=0.95 $Y=0.475 $X2=0 $Y2=0
cc_105 N_B_M1002_g N_A_M1003_g 0.0033853f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_106 N_B_c_126_n N_A_M1003_g 0.0187897f $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_107 N_B_M1002_g N_A_M1007_g 0.0231912f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_108 N_B_c_129_n N_A_M1007_g 9.99953e-19 $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_109 N_B_M1002_g N_A_c_161_n 0.0154653f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_110 N_B_M1002_g N_A_c_162_n 0.00212328f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_111 N_B_M1002_g N_A_27_297#_c_211_n 0.0112861f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_112 N_B_c_128_n N_A_27_297#_c_211_n 0.00103679f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_113 N_B_c_129_n N_A_27_297#_c_211_n 0.0815054f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_114 N_B_c_126_n N_A_27_297#_c_202_n 0.0166807f $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_115 N_B_c_129_n N_A_27_297#_c_238_n 0.0017825f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_116 N_B_c_129_n N_A_27_297#_c_213_n 0.0260771f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_117 N_B_M1002_g N_A_27_297#_c_214_n 0.00491229f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_118 N_B_c_129_n N_A_27_297#_c_214_n 0.0138062f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_119 N_B_M1002_g N_VPWR_c_308_n 0.00249809f $X=1.31 $Y=1.695 $X2=0 $Y2=0
cc_120 N_B_c_128_n N_VPWR_c_308_n 7.14013e-19 $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_121 N_B_c_129_n N_VPWR_c_308_n 0.0251801f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_122 N_B_c_128_n N_VPWR_c_309_n 0.00736312f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_123 N_B_c_129_n N_VPWR_c_309_n 0.0833171f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_124 N_B_c_128_n N_VPWR_c_307_n 0.0106165f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_125 N_B_c_129_n N_VPWR_c_307_n 0.0603546f $X=1.37 $Y=2.28 $X2=0 $Y2=0
cc_126 N_B_c_126_n N_VGND_c_353_n 0.00695614f $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_127 N_B_c_126_n N_VGND_c_354_n 5.25642e-19 $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_128 N_B_c_126_n N_VGND_c_356_n 0.00322006f $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_129 N_B_c_126_n N_VGND_c_358_n 0.00390029f $X=1.37 $Y=0.76 $X2=0 $Y2=0
cc_130 N_A_M1007_g N_A_27_297#_M1001_g 0.0190165f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_131 N_A_c_162_n N_A_27_297#_c_211_n 7.66792e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_c_162_n N_A_27_297#_c_202_n 3.58777e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_M1003_g N_A_27_297#_c_204_n 0.0116543f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_134 N_A_c_161_n N_A_27_297#_c_204_n 0.0020649f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_162_n N_A_27_297#_c_204_n 0.0166868f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_M1007_g N_A_27_297#_c_238_n 0.013079f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_137 N_A_c_162_n N_A_27_297#_c_238_n 0.0131508f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_M1007_g N_A_27_297#_c_212_n 0.0034529f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_139 N_A_c_161_n N_A_27_297#_c_205_n 6.92547e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_162_n N_A_27_297#_c_205_n 0.0146048f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_M1007_g N_A_27_297#_c_214_n 0.00166288f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_142 N_A_c_161_n N_A_27_297#_c_214_n 9.54211e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_162_n N_A_27_297#_c_214_n 0.0130691f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_c_161_n N_A_27_297#_c_206_n 0.00184138f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_162_n N_A_27_297#_c_206_n 0.026066f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_161_n N_A_27_297#_c_207_n 0.0202834f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_162_n N_A_27_297#_c_207_n 3.64881e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_M1003_g N_A_27_297#_c_208_n 0.0034529f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_149 N_A_M1003_g N_A_27_297#_c_209_n 0.0172443f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_VPWR_c_308_n 0.00298728f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_151 N_A_M1007_g N_VPWR_c_309_n 0.00264561f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_152 N_A_M1007_g N_VPWR_c_307_n 0.00333991f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_153 N_A_M1003_g N_VGND_c_353_n 5.2354e-19 $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_154 N_A_M1003_g N_VGND_c_354_n 0.00709299f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_155 N_A_M1003_g N_VGND_c_356_n 0.00322006f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_VGND_c_358_n 0.00390029f $X=1.79 $Y=0.475 $X2=0 $Y2=0
cc_157 N_A_27_297#_c_211_n A_109_297# 0.00243923f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_27_297#_c_211_n A_205_297# 0.00102299f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_159 N_A_27_297#_c_211_n A_277_297# 0.00246778f $X=1.51 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_27_297#_c_214_n A_277_297# 0.00525557f $X=1.595 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_27_297#_c_238_n N_VPWR_M1007_d 0.00526233f $X=2.065 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_162 N_A_27_297#_M1001_g N_VPWR_c_308_n 0.00485906f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_163 N_A_27_297#_c_238_n N_VPWR_c_308_n 0.0190361f $X=2.065 $Y=1.58 $X2=0
+ $Y2=0
cc_164 N_A_27_297#_c_214_n N_VPWR_c_308_n 0.0030545f $X=1.595 $Y=1.58 $X2=0
+ $Y2=0
cc_165 N_A_27_297#_c_207_n N_VPWR_c_308_n 2.30657e-19 $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_27_297#_M1001_g N_VPWR_c_310_n 0.00585385f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_27_297#_M1001_g N_VPWR_c_307_n 0.0128394f $X=2.28 $Y=1.985 $X2=0
+ $Y2=0
cc_168 N_A_27_297#_M1001_g N_X_c_334_n 0.00350509f $X=2.28 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A_27_297#_c_204_n N_X_c_334_n 0.00357198f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_27_297#_c_212_n N_X_c_334_n 0.00852743f $X=2.15 $Y=1.495 $X2=0 $Y2=0
cc_171 N_A_27_297#_c_206_n N_X_c_334_n 0.024425f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_297#_c_207_n N_X_c_334_n 0.00760589f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_27_297#_c_208_n N_X_c_334_n 0.00848187f $X=2.2 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_27_297#_c_209_n N_X_c_334_n 0.00442426f $X=2.252 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_27_297#_c_202_n N_VGND_M1009_d 0.00160115f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_c_204_n N_VGND_M1003_d 0.00482895f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_208_n N_VGND_M1003_d 6.98847e-19 $X=2.2 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_27_297#_c_283_p N_VGND_c_352_n 0.0182384f $X=0.71 $Y=0.47 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_283_p N_VGND_c_353_n 0.0117247f $X=0.71 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_202_n N_VGND_c_353_n 0.0160613f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_181 N_A_27_297#_c_204_n N_VGND_c_354_n 0.020701f $X=2.065 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_207_n N_VGND_c_354_n 2.52562e-19 $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_A_27_297#_c_209_n N_VGND_c_354_n 0.0132447f $X=2.252 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_27_297#_c_283_p N_VGND_c_355_n 0.00876148f $X=0.71 $Y=0.47 $X2=0
+ $Y2=0
cc_185 N_A_27_297#_c_202_n N_VGND_c_355_n 0.00276686f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_202_n N_VGND_c_356_n 0.00232396f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_c_292_p N_VGND_c_356_n 0.00846569f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_c_204_n N_VGND_c_356_n 0.00232396f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_c_204_n N_VGND_c_357_n 3.34073e-19 $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_c_209_n N_VGND_c_357_n 0.00524631f $X=2.252 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_c_283_p N_VGND_c_358_n 0.00625722f $X=0.71 $Y=0.47 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_202_n N_VGND_c_358_n 0.0105423f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_193 N_A_27_297#_c_292_p N_VGND_c_358_n 0.00625722f $X=1.58 $Y=0.47 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_204_n N_VGND_c_358_n 0.00637905f $X=2.065 $Y=0.74 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_209_n N_VGND_c_358_n 0.00951256f $X=2.252 $Y=0.995 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_307_n N_X_M1001_d 0.0039537f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_197 N_VPWR_c_310_n X 0.0187043f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_307_n X 0.0103212f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_199 N_X_c_333_n N_VGND_c_357_n 0.00876347f $X=2.59 $Y=0.587 $X2=0 $Y2=0
cc_200 N_X_M1006_d N_VGND_c_358_n 0.00411498f $X=2.355 $Y=0.235 $X2=0 $Y2=0
cc_201 N_X_c_333_n N_VGND_c_358_n 0.00924648f $X=2.59 $Y=0.587 $X2=0 $Y2=0

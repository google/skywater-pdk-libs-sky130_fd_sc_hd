* File: sky130_fd_sc_hd__o211a_4.pex.spice
* Created: Thu Aug 27 14:34:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__O211A_4%A_79_21# 1 2 3 4 13 15 18 20 22 25 27 29 32
+ 34 36 39 41 50 52 53 55 57 58 61 63 67 69 73 74 75 77 88
r161 85 86 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.72 $Y=1.16 $X2=1.73
+ $Y2=1.16
r162 84 85 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.31 $Y=1.16
+ $X2=1.72 $Y2=1.16
r163 83 84 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.29 $Y=1.16 $X2=1.31
+ $Y2=1.16
r164 82 83 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=0.89 $Y=1.16 $X2=1.29
+ $Y2=1.16
r165 81 82 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.86 $Y=1.16 $X2=0.89
+ $Y2=1.16
r166 70 75 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.12 $Y=1.94
+ $X2=3.952 $Y2=1.94
r167 69 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=1.94
+ $X2=5.32 $Y2=1.94
r168 69 70 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=5.155 $Y=1.94
+ $X2=4.12 $Y2=1.94
r169 65 75 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.952 $Y=2.025
+ $X2=3.952 $Y2=1.94
r170 65 67 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=3.952 $Y=2.025
+ $X2=3.952 $Y2=2.3
r171 64 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.06 $Y=1.94
+ $X2=2.88 $Y2=1.94
r172 63 75 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.785 $Y=1.94
+ $X2=3.952 $Y2=1.94
r173 63 64 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.785 $Y=1.94
+ $X2=3.06 $Y2=1.94
r174 59 74 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=2.025
+ $X2=2.88 $Y2=1.94
r175 59 61 8.80338 $w=3.58e-07 $l=2.75e-07 $layer=LI1_cond $X=2.88 $Y=2.025
+ $X2=2.88 $Y2=2.3
r176 57 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.7 $Y=1.94 $X2=2.88
+ $Y2=1.94
r177 57 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.7 $Y=1.94
+ $X2=2.37 $Y2=1.94
r178 53 55 60.6919 $w=1.78e-07 $l=9.85e-07 $layer=LI1_cond $X=2.37 $Y=0.725
+ $X2=3.355 $Y2=0.725
r179 52 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.285 $Y=1.855
+ $X2=2.37 $Y2=1.94
r180 51 73 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.265
+ $X2=2.285 $Y2=1.165
r181 51 52 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.285 $Y=1.265
+ $X2=2.285 $Y2=1.855
r182 50 73 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.285 $Y=1.065
+ $X2=2.285 $Y2=1.165
r183 49 53 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.285 $Y=0.815
+ $X2=2.37 $Y2=0.725
r184 49 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.285 $Y=0.815
+ $X2=2.285 $Y2=1.065
r185 48 88 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=1.16 $X2=2.15
+ $Y2=1.16
r186 48 86 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.06 $Y=1.16
+ $X2=1.73 $Y2=1.16
r187 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.16 $X2=2.06 $Y2=1.16
r188 44 81 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.7 $Y=1.16
+ $X2=0.86 $Y2=1.16
r189 44 78 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.7 $Y=1.16
+ $X2=0.47 $Y2=1.16
r190 43 47 75.4182 $w=1.98e-07 $l=1.36e-06 $layer=LI1_cond $X=0.7 $Y=1.165
+ $X2=2.06 $Y2=1.165
r191 43 44 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.16 $X2=0.7 $Y2=1.16
r192 41 73 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=1.165
+ $X2=2.285 $Y2=1.165
r193 41 47 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=2.2 $Y=1.165
+ $X2=2.06 $Y2=1.165
r194 37 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.16
r195 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=1.325
+ $X2=2.15 $Y2=1.985
r196 34 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=1.16
r197 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.73 $Y=0.995
+ $X2=1.73 $Y2=0.56
r198 30 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.325
+ $X2=1.72 $Y2=1.16
r199 30 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.72 $Y=1.325
+ $X2=1.72 $Y2=1.985
r200 27 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=1.16
r201 27 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.31 $Y2=0.56
r202 23 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.325
+ $X2=1.29 $Y2=1.16
r203 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.29 $Y=1.325
+ $X2=1.29 $Y2=1.985
r204 20 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=1.16
r205 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.89 $Y=0.995
+ $X2=0.89 $Y2=0.56
r206 16 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.86 $Y=1.325
+ $X2=0.86 $Y2=1.16
r207 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.86 $Y=1.325
+ $X2=0.86 $Y2=1.985
r208 13 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.16
r209 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r210 4 77 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=5.18
+ $Y=1.485 $X2=5.32 $Y2=2.02
r211 3 67 600 $w=1.7e-07 $l=9.13989e-07 $layer=licon1_PDIFF $count=1 $X=3.74
+ $Y=1.485 $X2=3.95 $Y2=2.3
r212 2 61 600 $w=1.7e-07 $l=9.27268e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=1.485 $X2=2.895 $Y2=2.3
r213 1 55 182 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.355 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%B1 3 7 10 13 17 18 20 21 26 29 30 31 33 36
c94 30 0 1.29314e-19 $X=4.115 $Y=1.16
r95 33 36 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=3.95 $Y=1.565
+ $X2=3.905 $Y2=1.565
r96 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.16
+ $X2=4.115 $Y2=1.325
r97 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.16
+ $X2=4.115 $Y2=0.995
r98 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.16 $X2=4.115 $Y2=1.16
r99 21 33 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=4.115 $Y=1.565
+ $X2=3.95 $Y2=1.565
r100 21 30 9.03851 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.115 $Y=1.445
+ $X2=4.115 $Y2=1.16
r101 21 36 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=3.885 $Y=1.565
+ $X2=3.905 $Y2=1.565
r102 20 21 50.6595 $w=2.38e-07 $l=1.055e-06 $layer=LI1_cond $X=2.83 $Y=1.565
+ $X2=3.885 $Y2=1.565
r103 18 27 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.637 $Y=1.16
+ $X2=2.637 $Y2=1.325
r104 18 26 48.0119 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.637 $Y=1.16
+ $X2=2.637 $Y2=0.995
r105 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.16 $X2=2.625 $Y2=1.16
r106 15 20 6.8957 $w=2.4e-07 $l=1.96023e-07 $layer=LI1_cond $X=2.685 $Y=1.445
+ $X2=2.83 $Y2=1.565
r107 15 17 11.3257 $w=2.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.685 $Y=1.445
+ $X2=2.685 $Y2=1.16
r108 13 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.205 $Y=1.985
+ $X2=4.205 $Y2=1.325
r109 10 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.095 $Y=0.56
+ $X2=4.095 $Y2=0.995
r110 7 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.71 $Y=0.56
+ $X2=2.71 $Y2=0.995
r111 3 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.58 $Y=1.985
+ $X2=2.58 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%C1 1 3 6 8 10 13 15 22 23
r46 21 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.575 $Y=1.16
+ $X2=3.665 $Y2=1.16
r47 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.575
+ $Y=1.16 $X2=3.575 $Y2=1.16
r48 19 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.235 $Y=1.16
+ $X2=3.575 $Y2=1.16
r49 17 19 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.16
+ $X2=3.235 $Y2=1.16
r50 15 22 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=3.445 $Y=1.155
+ $X2=3.575 $Y2=1.155
r51 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.325
+ $X2=3.665 $Y2=1.16
r52 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.665 $Y=1.325
+ $X2=3.665 $Y2=1.985
r53 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=0.995
+ $X2=3.665 $Y2=1.16
r54 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.665 $Y=0.995
+ $X2=3.665 $Y2=0.56
r55 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.325
+ $X2=3.235 $Y2=1.16
r56 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.235 $Y=1.325
+ $X2=3.235 $Y2=1.985
r57 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=0.995
+ $X2=3.07 $Y2=1.16
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.07 $Y=0.995 $X2=3.07
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%A1 3 6 10 13 17 18 20 21 22 26 29 30 31 33
c82 17 0 1.99978e-19 $X=4.655 $Y=1.16
c83 6 0 1.29314e-19 $X=4.675 $Y=1.985
r84 29 32 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.09 $Y=1.16 $X2=6.09
+ $Y2=1.325
r85 29 31 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.09 $Y=1.16 $X2=6.09
+ $Y2=0.995
r86 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=1.16 $X2=6.085 $Y2=1.16
r87 22 33 2.57785 $w=4e-07 $l=9.5e-08 $layer=LI1_cond $X=6.09 $Y=1.59 $X2=6.09
+ $Y2=1.495
r88 22 33 0.720277 $w=3.98e-07 $l=2.5e-08 $layer=LI1_cond $X=6.09 $Y=1.47
+ $X2=6.09 $Y2=1.495
r89 22 30 8.93143 $w=3.98e-07 $l=3.1e-07 $layer=LI1_cond $X=6.09 $Y=1.47
+ $X2=6.09 $Y2=1.16
r90 20 22 5.42706 $w=1.9e-07 $l=2e-07 $layer=LI1_cond $X=5.89 $Y=1.59 $X2=6.09
+ $Y2=1.59
r91 20 21 61 $w=1.88e-07 $l=1.045e-06 $layer=LI1_cond $X=5.89 $Y=1.59 $X2=4.845
+ $Y2=1.59
r92 18 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.16
+ $X2=4.655 $Y2=1.325
r93 18 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.16
+ $X2=4.655 $Y2=0.995
r94 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.655
+ $Y=1.16 $X2=4.655 $Y2=1.16
r95 15 21 7.66236 $w=1.9e-07 $l=2.2044e-07 $layer=LI1_cond $X=4.667 $Y=1.495
+ $X2=4.845 $Y2=1.59
r96 15 17 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=4.667 $Y=1.495
+ $X2=4.667 $Y2=1.16
r97 13 32 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.965 $Y=1.985
+ $X2=5.965 $Y2=1.325
r98 10 31 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.965 $Y=0.56
+ $X2=5.965 $Y2=0.995
r99 6 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.675 $Y=1.985
+ $X2=4.675 $Y2=1.325
r100 3 26 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.565 $Y=0.56
+ $X2=4.565 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%A2 1 3 6 8 10 13 15 20 21
r52 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.535
+ $Y=1.16 $X2=5.535 $Y2=1.16
r53 17 20 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.105 $Y=1.16
+ $X2=5.535 $Y2=1.16
r54 15 21 9.93485 $w=2.88e-07 $l=2.5e-07 $layer=LI1_cond $X=5.285 $Y=1.18
+ $X2=5.535 $Y2=1.18
r55 11 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.16
r56 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.535 $Y=1.325
+ $X2=5.535 $Y2=1.985
r57 8 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=1.16
r58 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.535 $Y=0.995
+ $X2=5.535 $Y2=0.56
r59 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.325
+ $X2=5.105 $Y2=1.16
r60 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.105 $Y=1.325
+ $X2=5.105 $Y2=1.985
r61 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=0.995
+ $X2=5.105 $Y2=1.16
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.105 $Y=0.995
+ $X2=5.105 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%VPWR 1 2 3 4 5 6 21 25 29 33 35 39 41 43 46
+ 47 49 50 51 53 65 69 78 81 84 88
c109 5 0 8.47117e-20 $X=4.28 $Y=1.485
r110 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r112 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r113 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r114 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 76 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r116 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r117 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r118 73 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r119 72 75 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r120 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r121 70 84 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.422 $Y2=2.72
r122 70 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 69 87 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=6.015 $Y=2.72
+ $X2=6.227 $Y2=2.72
r124 69 75 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.015 $Y=2.72
+ $X2=5.75 $Y2=2.72
r125 68 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r127 65 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.45 $Y2=2.72
r128 65 67 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=2.99 $Y2=2.72
r129 64 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r130 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r131 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r132 61 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r133 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r134 58 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=2.72
+ $X2=0.645 $Y2=2.72
r135 58 60 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.81 $Y=2.72
+ $X2=1.15 $Y2=2.72
r136 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.48 $Y=2.72
+ $X2=0.645 $Y2=2.72
r137 53 55 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.48 $Y=2.72
+ $X2=0.23 $Y2=2.72
r138 51 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r139 51 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r140 49 63 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=2.72
+ $X2=2.365 $Y2=2.72
r142 48 67 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r143 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.365 $Y2=2.72
r144 46 60 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.34 $Y=2.72
+ $X2=1.15 $Y2=2.72
r145 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=2.72
+ $X2=1.505 $Y2=2.72
r146 45 63 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.67 $Y=2.72 $X2=2.07
+ $Y2=2.72
r147 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=2.72
+ $X2=1.505 $Y2=2.72
r148 41 87 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.18 $Y=2.635
+ $X2=6.227 $Y2=2.72
r149 41 43 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.18 $Y=2.635
+ $X2=6.18 $Y2=2
r150 37 84 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.422 $Y=2.635
+ $X2=4.422 $Y2=2.72
r151 37 39 11.9593 $w=2.63e-07 $l=2.75e-07 $layer=LI1_cond $X=4.422 $Y=2.635
+ $X2=4.422 $Y2=2.36
r152 36 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.45 $Y2=2.72
r153 35 84 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=4.422 $Y2=2.72
r154 35 36 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.29 $Y=2.72
+ $X2=3.615 $Y2=2.72
r155 31 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=2.635
+ $X2=3.45 $Y2=2.72
r156 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.45 $Y=2.635
+ $X2=3.45 $Y2=2.36
r157 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=2.635
+ $X2=2.365 $Y2=2.72
r158 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.365 $Y=2.635
+ $X2=2.365 $Y2=2.32
r159 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=2.635
+ $X2=1.505 $Y2=2.72
r160 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.505 $Y=2.635
+ $X2=1.505 $Y2=1.955
r161 19 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=2.635
+ $X2=0.645 $Y2=2.72
r162 19 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.645 $Y=2.635
+ $X2=0.645 $Y2=1.955
r163 6 43 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=6.04
+ $Y=1.485 $X2=6.18 $Y2=2
r164 5 39 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.485 $X2=4.42 $Y2=2.36
r165 4 33 600 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.485 $X2=3.45 $Y2=2.36
r166 3 29 600 $w=1.7e-07 $l=9.02289e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.485 $X2=2.365 $Y2=2.32
r167 2 25 300 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=2 $X=1.365
+ $Y=1.485 $X2=1.505 $Y2=1.955
r168 1 21 300 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_PDIFF $count=2 $X=0.52
+ $Y=1.485 $X2=0.645 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%X 1 2 3 4 13 15 16 19 21 25 27 31 35 38 39
+ 40 43 45
r58 43 45 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.225 $Y=0.805
+ $X2=0.225 $Y2=0.85
r59 40 43 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=0.72
+ $X2=0.225 $Y2=0.805
r60 40 45 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=0.225 $Y=0.87
+ $X2=0.225 $Y2=0.85
r61 37 40 23.2547 $w=2.78e-07 $l=5.65e-07 $layer=LI1_cond $X=0.225 $Y=1.435
+ $X2=0.225 $Y2=0.87
r62 33 35 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.935 $Y=1.7
+ $X2=1.935 $Y2=1.845
r63 29 31 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.52 $Y=0.615
+ $X2=1.52 $Y2=0.42
r64 28 39 3.70371 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.16 $Y=1.567 $X2=1.07
+ $Y2=1.567
r65 27 33 7.06018 $w=2.65e-07 $l=1.74138e-07 $layer=LI1_cond $X=1.84 $Y=1.567
+ $X2=1.935 $Y2=1.7
r66 27 28 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=1.84 $Y=1.567
+ $X2=1.16 $Y2=1.567
r67 23 39 2.76582 $w=1.8e-07 $l=1.33e-07 $layer=LI1_cond $X=1.07 $Y=1.7 $X2=1.07
+ $Y2=1.567
r68 23 25 8.93434 $w=1.78e-07 $l=1.45e-07 $layer=LI1_cond $X=1.07 $Y=1.7
+ $X2=1.07 $Y2=1.845
r69 22 38 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.71
+ $X2=0.68 $Y2=0.71
r70 21 29 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.435 $Y=0.71
+ $X2=1.52 $Y2=0.615
r71 21 22 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=1.435 $Y=0.71
+ $X2=0.765 $Y2=0.71
r72 17 38 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.68 $Y=0.615
+ $X2=0.68 $Y2=0.71
r73 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.68 $Y=0.615
+ $X2=0.68 $Y2=0.42
r74 16 37 6.82321 $w=2.65e-07 $l=1.95141e-07 $layer=LI1_cond $X=0.365 $Y=1.567
+ $X2=0.225 $Y2=1.435
r75 15 39 3.70371 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=0.98 $Y=1.567 $X2=1.07
+ $Y2=1.567
r76 15 16 26.7454 $w=2.63e-07 $l=6.15e-07 $layer=LI1_cond $X=0.98 $Y=1.567
+ $X2=0.365 $Y2=1.567
r77 14 40 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=0.72
+ $X2=0.225 $Y2=0.72
r78 13 38 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.68 $Y2=0.71
r79 13 14 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.595 $Y=0.72
+ $X2=0.365 $Y2=0.72
r80 4 35 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=1.795
+ $Y=1.485 $X2=1.935 $Y2=1.845
r81 3 25 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=0.935
+ $Y=1.485 $X2=1.075 $Y2=1.845
r82 2 31 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.385
+ $Y=0.235 $X2=1.52 $Y2=0.42
r83 1 19 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 60 61 67 70 73 76
r102 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r103 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r104 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r105 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r106 61 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r107 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r108 58 76 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.845 $Y=0 $X2=5.75
+ $Y2=0
r109 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.845 $Y=0
+ $X2=6.21 $Y2=0
r110 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r111 57 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r112 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r113 54 73 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=4.985 $Y=0
+ $X2=4.827 $Y2=0
r114 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.985 $Y=0
+ $X2=5.29 $Y2=0
r115 53 76 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.75
+ $Y2=0
r116 53 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.655 $Y=0
+ $X2=5.29 $Y2=0
r117 52 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r118 52 71 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=2.07
+ $Y2=0
r119 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r120 49 70 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=1.957
+ $Y2=0
r121 49 51 145.487 $w=1.68e-07 $l=2.23e-06 $layer=LI1_cond $X=2.14 $Y=0 $X2=4.37
+ $Y2=0
r122 48 73 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.827
+ $Y2=0
r123 48 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.37
+ $Y2=0
r124 47 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r125 47 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r126 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r127 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r128 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.61
+ $Y2=0
r129 43 70 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.957 $Y2=0
r130 43 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=1.61 $Y2=0
r131 42 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r132 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r133 39 64 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r134 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r135 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r136 38 41 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.69
+ $Y2=0
r137 36 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r138 36 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r139 32 76 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.75 $Y=0.085
+ $X2=5.75 $Y2=0
r140 32 34 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=5.75 $Y=0.085
+ $X2=5.75 $Y2=0.36
r141 28 73 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.827 $Y=0.085
+ $X2=4.827 $Y2=0
r142 28 30 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=4.827 $Y=0.085
+ $X2=4.827 $Y2=0.36
r143 24 70 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0
r144 24 26 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.957 $Y=0.085
+ $X2=1.957 $Y2=0.38
r145 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r146 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.36
r147 16 64 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r148 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r149 5 34 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.235 $X2=5.75 $Y2=0.36
r150 4 30 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.64
+ $Y=0.235 $X2=4.82 $Y2=0.36
r151 3 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.235 $X2=1.94 $Y2=0.38
r152 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.36
r153 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HD__O211A_4%A_474_47# 1 2 3 4 13 17 18 19 20 23 25 29 33
r71 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.18 $Y=0.695
+ $X2=6.18 $Y2=0.38
r72 26 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.485 $Y=0.78
+ $X2=5.32 $Y2=0.78
r73 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.015 $Y=0.78
+ $X2=6.18 $Y2=0.695
r74 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.015 $Y=0.78
+ $X2=5.485 $Y2=0.78
r75 21 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.32 $Y=0.695
+ $X2=5.32 $Y2=0.78
r76 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.32 $Y=0.695
+ $X2=5.32 $Y2=0.36
r77 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0.78
+ $X2=5.32 $Y2=0.78
r78 19 20 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.155 $Y=0.78
+ $X2=4.5 $Y2=0.78
r79 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.335 $Y=0.695
+ $X2=4.5 $Y2=0.78
r80 17 32 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.335 $Y=0.465
+ $X2=4.335 $Y2=0.36
r81 17 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.335 $Y=0.465
+ $X2=4.335 $Y2=0.695
r82 13 32 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.17 $Y=0.36
+ $X2=4.335 $Y2=0.36
r83 13 15 88.4632 $w=2.08e-07 $l=1.675e-06 $layer=LI1_cond $X=4.17 $Y=0.36
+ $X2=2.495 $Y2=0.36
r84 4 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.04
+ $Y=0.235 $X2=6.18 $Y2=0.38
r85 3 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.18
+ $Y=0.235 $X2=5.32 $Y2=0.36
r86 2 32 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.17
+ $Y=0.235 $X2=4.335 $Y2=0.42
r87 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.37
+ $Y=0.235 $X2=2.495 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__ha_4.pxi.spice
* Created: Tue Sep  1 19:09:37 2020
* 
x_PM_SKY130_FD_SC_HD__HA_4%A_79_21# N_A_79_21#_M1015_s N_A_79_21#_M1002_d
+ N_A_79_21#_M1007_s N_A_79_21#_c_146_n N_A_79_21#_M1014_g N_A_79_21#_M1005_g
+ N_A_79_21#_c_147_n N_A_79_21#_M1020_g N_A_79_21#_M1011_g N_A_79_21#_c_148_n
+ N_A_79_21#_M1021_g N_A_79_21#_M1022_g N_A_79_21#_c_149_n N_A_79_21#_M1031_g
+ N_A_79_21#_M1030_g N_A_79_21#_c_150_n N_A_79_21#_c_151_n N_A_79_21#_c_152_n
+ N_A_79_21#_c_153_n N_A_79_21#_c_160_n N_A_79_21#_c_164_p N_A_79_21#_c_169_p
+ N_A_79_21#_c_213_p N_A_79_21#_c_166_p N_A_79_21#_c_162_p N_A_79_21#_c_167_p
+ N_A_79_21#_c_191_p N_A_79_21#_c_175_p N_A_79_21#_c_173_p
+ PM_SKY130_FD_SC_HD__HA_4%A_79_21#
x_PM_SKY130_FD_SC_HD__HA_4%A_514_199# N_A_514_199#_M1000_d N_A_514_199#_M1029_d
+ N_A_514_199#_M1018_d N_A_514_199#_M1002_g N_A_514_199#_c_286_n
+ N_A_514_199#_M1015_g N_A_514_199#_M1016_g N_A_514_199#_c_287_n
+ N_A_514_199#_M1017_g N_A_514_199#_c_288_n N_A_514_199#_M1001_g
+ N_A_514_199#_M1008_g N_A_514_199#_c_289_n N_A_514_199#_M1004_g
+ N_A_514_199#_M1019_g N_A_514_199#_c_290_n N_A_514_199#_M1010_g
+ N_A_514_199#_M1027_g N_A_514_199#_c_291_n N_A_514_199#_M1012_g
+ N_A_514_199#_M1035_g N_A_514_199#_c_303_n N_A_514_199#_c_304_n
+ N_A_514_199#_c_305_n N_A_514_199#_c_386_p N_A_514_199#_c_327_n
+ N_A_514_199#_c_329_n N_A_514_199#_c_411_p N_A_514_199#_c_363_p
+ N_A_514_199#_c_343_p N_A_514_199#_c_415_p N_A_514_199#_c_393_p
+ N_A_514_199#_c_348_p N_A_514_199#_c_345_p N_A_514_199#_c_368_p
+ N_A_514_199#_c_292_n N_A_514_199#_c_293_n N_A_514_199#_c_449_p
+ N_A_514_199#_c_365_p N_A_514_199#_c_379_p N_A_514_199#_c_294_n
+ N_A_514_199#_c_295_n N_A_514_199#_c_296_n PM_SKY130_FD_SC_HD__HA_4%A_514_199#
x_PM_SKY130_FD_SC_HD__HA_4%A N_A_c_506_n N_A_M1013_g N_A_M1026_g N_A_M1028_g
+ N_A_c_507_n N_A_M1024_g N_A_M1029_g N_A_c_508_n N_A_M1009_g N_A_c_509_n
+ N_A_M1033_g N_A_M1034_g N_A_c_510_n N_A_c_511_n N_A_c_520_n N_A_c_552_n
+ N_A_c_530_n N_A_c_521_n N_A_c_512_n N_A_c_554_n A A N_A_c_513_n N_A_c_514_n
+ N_A_c_575_n PM_SKY130_FD_SC_HD__HA_4%A
x_PM_SKY130_FD_SC_HD__HA_4%B N_B_c_662_n N_B_M1023_g N_B_M1007_g N_B_c_663_n
+ N_B_M1025_g N_B_M1032_g N_B_c_664_n N_B_M1000_g N_B_M1003_g N_B_c_665_n
+ N_B_M1006_g N_B_M1018_g N_B_c_666_n N_B_c_667_n N_B_c_723_n N_B_c_668_n
+ N_B_c_669_n N_B_c_670_n B B N_B_c_671_n N_B_c_698_n B
+ PM_SKY130_FD_SC_HD__HA_4%B
x_PM_SKY130_FD_SC_HD__HA_4%VPWR N_VPWR_M1005_s N_VPWR_M1011_s N_VPWR_M1030_s
+ N_VPWR_M1016_s N_VPWR_M1028_d N_VPWR_M1003_s N_VPWR_M1034_s N_VPWR_M1019_s
+ N_VPWR_M1035_s N_VPWR_c_791_n N_VPWR_c_792_n N_VPWR_c_793_n N_VPWR_c_794_n
+ N_VPWR_c_795_n N_VPWR_c_796_n N_VPWR_c_797_n N_VPWR_c_798_n N_VPWR_c_799_n
+ N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n
+ N_VPWR_c_805_n N_VPWR_c_806_n N_VPWR_c_807_n VPWR N_VPWR_c_808_n
+ N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n
+ N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_790_n
+ PM_SKY130_FD_SC_HD__HA_4%VPWR
x_PM_SKY130_FD_SC_HD__HA_4%SUM N_SUM_M1014_s N_SUM_M1021_s N_SUM_M1005_d
+ N_SUM_M1022_d N_SUM_c_936_n N_SUM_c_941_n N_SUM_c_935_n N_SUM_c_947_n
+ N_SUM_c_949_n N_SUM_c_952_n N_SUM_c_955_n N_SUM_c_937_n SUM SUM SUM SUM SUM
+ SUM N_SUM_c_966_n PM_SKY130_FD_SC_HD__HA_4%SUM
x_PM_SKY130_FD_SC_HD__HA_4%COUT N_COUT_M1001_s N_COUT_M1010_s N_COUT_M1008_d
+ N_COUT_M1027_d N_COUT_c_999_n N_COUT_c_1028_n N_COUT_c_996_n N_COUT_c_997_n
+ N_COUT_c_993_n N_COUT_c_994_n COUT COUT COUT COUT COUT COUT
+ PM_SKY130_FD_SC_HD__HA_4%COUT
x_PM_SKY130_FD_SC_HD__HA_4%VGND N_VGND_M1014_d N_VGND_M1020_d N_VGND_M1031_d
+ N_VGND_M1013_d N_VGND_M1025_d N_VGND_M1024_d N_VGND_M1033_s N_VGND_M1004_d
+ N_VGND_M1012_d N_VGND_c_1045_n N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n
+ N_VGND_c_1049_n N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n
+ N_VGND_c_1053_n N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n
+ N_VGND_c_1057_n N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n
+ N_VGND_c_1061_n N_VGND_c_1062_n N_VGND_c_1063_n N_VGND_c_1064_n VGND
+ N_VGND_c_1065_n N_VGND_c_1066_n N_VGND_c_1067_n N_VGND_c_1068_n
+ N_VGND_c_1069_n N_VGND_c_1070_n N_VGND_c_1071_n PM_SKY130_FD_SC_HD__HA_4%VGND
x_PM_SKY130_FD_SC_HD__HA_4%A_467_47# N_A_467_47#_M1015_d N_A_467_47#_M1017_d
+ N_A_467_47#_M1023_s N_A_467_47#_M1024_s N_A_467_47#_c_1196_n
+ N_A_467_47#_c_1208_n N_A_467_47#_c_1207_n N_A_467_47#_c_1237_n
+ N_A_467_47#_c_1197_n N_A_467_47#_c_1214_n N_A_467_47#_c_1198_n
+ PM_SKY130_FD_SC_HD__HA_4%A_467_47#
cc_1 VNB N_A_79_21#_c_146_n 0.0215085f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_147_n 0.0155244f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.995
cc_3 VNB N_A_79_21#_c_148_n 0.0155244f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_4 VNB N_A_79_21#_c_149_n 0.021952f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_5 VNB N_A_79_21#_c_150_n 0.0706848f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_6 VNB N_A_79_21#_c_151_n 0.0104117f $X=-0.19 $Y=-0.24 $X2=2.58 $Y2=1.16
cc_7 VNB N_A_79_21#_c_152_n 0.0422176f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.16
cc_8 VNB N_A_79_21#_c_153_n 0.0048714f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.075
cc_9 VNB N_A_514_199#_c_286_n 0.0194565f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_10 VNB N_A_514_199#_c_287_n 0.0162331f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_11 VNB N_A_514_199#_c_288_n 0.0168747f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_12 VNB N_A_514_199#_c_289_n 0.015773f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_13 VNB N_A_514_199#_c_290_n 0.0157605f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_14 VNB N_A_514_199#_c_291_n 0.0214956f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.16
cc_15 VNB N_A_514_199#_c_292_n 0.00322284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_514_199#_c_293_n 8.78812e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_514_199#_c_294_n 0.00102135f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_514_199#_c_295_n 0.0318455f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_514_199#_c_296_n 0.0753769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_c_506_n 0.016456f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=0.235
cc_21 VNB N_A_c_507_n 0.0212707f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_22 VNB N_A_c_508_n 0.015494f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=0.56
cc_23 VNB N_A_c_509_n 0.0171598f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_24 VNB N_A_c_510_n 0.00696273f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_25 VNB N_A_c_511_n 0.0202312f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_26 VNB N_A_c_512_n 0.044017f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.16
cc_27 VNB N_A_c_513_n 0.0210049f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=1.935
cc_28 VNB N_A_c_514_n 0.00244043f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=2.19
cc_29 VNB N_B_c_662_n 0.016213f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=0.235
cc_30 VNB N_B_c_663_n 0.0210871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B_c_664_n 0.0152697f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.985
cc_32 VNB N_B_c_665_n 0.0162222f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.985
cc_33 VNB N_B_c_666_n 0.0254277f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_34 VNB N_B_c_667_n 0.0088186f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.56
cc_35 VNB N_B_c_668_n 0.00158877f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_36 VNB N_B_c_669_n 0.02698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_B_c_670_n 9.76635e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_38 VNB N_B_c_671_n 0.0298886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB B 0.00108852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_790_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_SUM_c_935_n 0.00103446f $X=-0.19 $Y=-0.24 $X2=0.89 $Y2=1.325
cc_42 VNB N_COUT_c_993_n 0.00245684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_COUT_c_994_n 0.00187796f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.995
cc_44 VNB COUT 8.54099e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=0.56
cc_45 VNB N_VGND_c_1045_n 0.0105466f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.985
cc_46 VNB N_VGND_c_1046_n 0.00773781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_1047_n 0.00479928f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.325
cc_48 VNB N_VGND_c_1048_n 0.0137204f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.16
cc_49 VNB N_VGND_c_1049_n 3.95589e-19 $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.16
cc_50 VNB N_VGND_c_1050_n 0.00450741f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.16
cc_51 VNB N_VGND_c_1051_n 4.1623e-19 $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.075
cc_52 VNB N_VGND_c_1052_n 0.00504069f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=0.73
cc_53 VNB N_VGND_c_1053_n 0.0172422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1054_n 0.00377775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1055_n 0.0105466f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.85
cc_56 VNB N_VGND_c_1056_n 0.00769352f $X=-0.19 $Y=-0.24 $X2=3.615 $Y2=2.205
cc_57 VNB N_VGND_c_1057_n 0.018513f $X=-0.19 $Y=-0.24 $X2=4.165 $Y2=2.29
cc_58 VNB N_VGND_c_1058_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1059_n 0.0351166f $X=-0.19 $Y=-0.24 $X2=2.665 $Y2=1.85
cc_60 VNB N_VGND_c_1060_n 0.00469392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1061_n 0.0112489f $X=-0.19 $Y=-0.24 $X2=2.855 $Y2=1.85
cc_62 VNB N_VGND_c_1062_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=2.225 $Y2=1.16
cc_63 VNB N_VGND_c_1063_n 0.0154216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1064_n 0.00436154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1065_n 0.018513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1066_n 0.0327098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1067_n 0.0169941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1068_n 0.00461634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1069_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1070_n 0.00401244f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1071_n 0.441009f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_467_47#_c_1196_n 0.00288768f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.325
cc_73 VNB N_A_467_47#_c_1197_n 0.00544388f $X=-0.19 $Y=-0.24 $X2=1.31 $Y2=1.325
cc_74 VNB N_A_467_47#_c_1198_n 0.00567359f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.995
cc_75 VPB N_A_79_21#_M1005_g 0.025289f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.985
cc_76 VPB N_A_79_21#_M1011_g 0.0177497f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_77 VPB N_A_79_21#_M1022_g 0.0177497f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_78 VPB N_A_79_21#_M1030_g 0.0259414f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_79 VPB N_A_79_21#_c_150_n 0.0117672f $X=-0.19 $Y=1.305 $X2=1.805 $Y2=1.16
cc_80 VPB N_A_79_21#_c_152_n 0.0162404f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.16
cc_81 VPB N_A_79_21#_c_160_n 9.82205e-19 $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.765
cc_82 VPB N_A_514_199#_M1002_g 0.0252902f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_83 VPB N_A_514_199#_M1016_g 0.0180555f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.56
cc_84 VPB N_A_514_199#_M1008_g 0.0195672f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_85 VPB N_A_514_199#_M1019_g 0.0176322f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_86 VPB N_A_514_199#_M1027_g 0.0178427f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_87 VPB N_A_514_199#_M1035_g 0.025289f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.075
cc_88 VPB N_A_514_199#_c_303_n 6.03256e-19 $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.73
cc_89 VPB N_A_514_199#_c_304_n 0.00752569f $X=-0.19 $Y=1.305 $X2=2.855 $Y2=1.935
cc_90 VPB N_A_514_199#_c_305_n 3.73621e-19 $X=-0.19 $Y=1.305 $X2=2.855 $Y2=2.19
cc_91 VPB N_A_514_199#_c_293_n 0.00319264f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_514_199#_c_295_n 0.00527486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_514_199#_c_296_n 0.0112432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_M1026_g 0.0189695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_M1028_g 0.0235374f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_96 VPB N_A_M1029_g 0.0190815f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=0.995
cc_97 VPB N_A_M1034_g 0.0199143f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_98 VPB N_A_c_511_n 0.00406199f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.56
cc_99 VPB N_A_c_520_n 0.00132188f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_100 VPB N_A_c_521_n 0.00358543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_c_512_n 0.0112638f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.16
cc_102 VPB A 0.00180656f $X=-0.19 $Y=1.305 $X2=2.225 $Y2=1.16
cc_103 VPB N_A_c_513_n 0.00490685f $X=-0.19 $Y=1.305 $X2=2.855 $Y2=1.935
cc_104 VPB N_A_c_514_n 9.18598e-19 $X=-0.19 $Y=1.305 $X2=2.855 $Y2=2.19
cc_105 VPB N_B_M1007_g 0.018456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_B_M1032_g 0.0209159f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_107 VPB N_B_M1003_g 0.0185702f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.325
cc_108 VPB N_B_M1018_g 0.0176621f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.325
cc_109 VPB N_B_c_666_n 0.0043858f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_110 VPB N_B_c_668_n 0.00158877f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.16
cc_111 VPB N_B_c_669_n 0.0106819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_B_c_671_n 0.00400964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_791_n 0.0105207f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.985
cc_114 VPB N_VPWR_c_792_n 0.00440046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_793_n 0.00361209f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.985
cc_116 VPB N_VPWR_c_794_n 0.00606736f $X=-0.19 $Y=1.305 $X2=1.31 $Y2=1.16
cc_117 VPB N_VPWR_c_795_n 0.00470515f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_796_n 0.00503623f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.765
cc_119 VPB N_VPWR_c_797_n 0.0151348f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.73
cc_120 VPB N_VPWR_c_798_n 3.25223e-19 $X=-0.19 $Y=1.305 $X2=2.855 $Y2=2.19
cc_121 VPB N_VPWR_c_799_n 0.0136014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_800_n 0.00426714f $X=-0.19 $Y=1.305 $X2=3.615 $Y2=2.205
cc_123 VPB N_VPWR_c_801_n 0.00192314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_802_n 0.0105207f $X=-0.19 $Y=1.305 $X2=2.665 $Y2=1.85
cc_125 VPB N_VPWR_c_803_n 0.00435617f $X=-0.19 $Y=1.305 $X2=2.855 $Y2=1.85
cc_126 VPB N_VPWR_c_804_n 0.0184587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_805_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_806_n 0.0249151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_807_n 0.00324452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_808_n 0.0184587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_809_n 0.0498767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_810_n 0.0149139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_811_n 0.0176124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_812_n 0.00978383f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_813_n 0.00631736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_814_n 0.00436447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_815_n 0.00631736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_816_n 0.00430944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_790_n 0.047372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_SUM_c_936_n 0.00529213f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.325
cc_141 VPB N_SUM_c_937_n 0.00140122f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=0.995
cc_142 VPB N_COUT_c_996_n 0.00290698f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_143 VPB N_COUT_c_997_n 0.00180692f $X=-0.19 $Y=1.305 $X2=0.89 $Y2=1.985
cc_144 VPB COUT 8.54099e-19 $X=-0.19 $Y=1.305 $X2=1.31 $Y2=0.56
cc_145 N_A_79_21#_c_160_n N_A_514_199#_M1002_g 0.0152407f $X=2.665 $Y=1.765
+ $X2=0 $Y2=0
cc_146 N_A_79_21#_c_162_p N_A_514_199#_M1002_g 0.00685925f $X=2.94 $Y=1.85 $X2=0
+ $Y2=0
cc_147 N_A_79_21#_c_153_n N_A_514_199#_c_286_n 0.00529625f $X=2.665 $Y=1.075
+ $X2=0 $Y2=0
cc_148 N_A_79_21#_c_164_p N_A_514_199#_c_286_n 0.00692262f $X=2.75 $Y=0.73 $X2=0
+ $Y2=0
cc_149 N_A_79_21#_c_160_n N_A_514_199#_M1016_g 5.00502e-19 $X=2.665 $Y=1.765
+ $X2=0 $Y2=0
cc_150 N_A_79_21#_c_166_p N_A_514_199#_M1016_g 0.00985962f $X=3.53 $Y=1.85 $X2=0
+ $Y2=0
cc_151 N_A_79_21#_c_167_p N_A_514_199#_M1016_g 5.08404e-19 $X=3.615 $Y=2.205
+ $X2=0 $Y2=0
cc_152 N_A_79_21#_c_153_n N_A_514_199#_c_287_n 0.00200082f $X=2.665 $Y=1.075
+ $X2=0 $Y2=0
cc_153 N_A_79_21#_c_169_p N_A_514_199#_c_287_n 0.00255625f $X=2.88 $Y=0.73 $X2=0
+ $Y2=0
cc_154 N_A_79_21#_c_153_n N_A_514_199#_c_303_n 0.00538854f $X=2.665 $Y=1.075
+ $X2=0 $Y2=0
cc_155 N_A_79_21#_c_160_n N_A_514_199#_c_303_n 0.0128787f $X=2.665 $Y=1.765
+ $X2=0 $Y2=0
cc_156 N_A_79_21#_c_169_p N_A_514_199#_c_303_n 0.00713004f $X=2.88 $Y=0.73 $X2=0
+ $Y2=0
cc_157 N_A_79_21#_c_173_p N_A_514_199#_c_303_n 0.0129498f $X=2.665 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_79_21#_c_166_p N_A_514_199#_c_304_n 0.0317358f $X=3.53 $Y=1.85 $X2=0
+ $Y2=0
cc_159 N_A_79_21#_c_175_p N_A_514_199#_c_304_n 0.00342031f $X=4.165 $Y=2.29
+ $X2=0 $Y2=0
cc_160 N_A_79_21#_M1002_d N_A_514_199#_c_305_n 0.00110104f $X=2.72 $Y=1.485
+ $X2=0 $Y2=0
cc_161 N_A_79_21#_c_160_n N_A_514_199#_c_305_n 0.00996512f $X=2.665 $Y=1.765
+ $X2=0 $Y2=0
cc_162 N_A_79_21#_c_162_p N_A_514_199#_c_305_n 0.00851043f $X=2.94 $Y=1.85 $X2=0
+ $Y2=0
cc_163 N_A_79_21#_M1007_s N_A_514_199#_c_327_n 0.0041802f $X=4.03 $Y=1.485 $X2=0
+ $Y2=0
cc_164 N_A_79_21#_c_175_p N_A_514_199#_c_327_n 0.0121596f $X=4.165 $Y=2.29 $X2=0
+ $Y2=0
cc_165 N_A_79_21#_c_175_p N_A_514_199#_c_329_n 0.0102065f $X=4.165 $Y=2.29 $X2=0
+ $Y2=0
cc_166 N_A_79_21#_c_151_n N_A_514_199#_c_295_n 0.00223682f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_79_21#_c_152_n N_A_514_199#_c_295_n 0.0231397f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_79_21#_c_153_n N_A_514_199#_c_295_n 0.00355434f $X=2.665 $Y=1.075
+ $X2=0 $Y2=0
cc_169 N_A_79_21#_c_160_n N_A_514_199#_c_295_n 0.00326238f $X=2.665 $Y=1.765
+ $X2=0 $Y2=0
cc_170 N_A_79_21#_c_169_p N_A_514_199#_c_295_n 0.00327786f $X=2.88 $Y=0.73 $X2=0
+ $Y2=0
cc_171 N_A_79_21#_c_162_p N_A_514_199#_c_295_n 0.00261723f $X=2.94 $Y=1.85 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_c_173_p N_A_514_199#_c_295_n 0.00508446f $X=2.665 $Y=1.16
+ $X2=0 $Y2=0
cc_173 N_A_79_21#_c_166_p N_A_M1026_g 0.0098276f $X=3.53 $Y=1.85 $X2=0 $Y2=0
cc_174 N_A_79_21#_c_167_p N_A_M1026_g 0.00652432f $X=3.615 $Y=2.205 $X2=0 $Y2=0
cc_175 N_A_79_21#_c_191_p N_A_M1026_g 0.00485067f $X=3.7 $Y=2.29 $X2=0 $Y2=0
cc_176 N_A_79_21#_c_175_p N_A_M1028_g 7.02707e-19 $X=4.165 $Y=2.29 $X2=0 $Y2=0
cc_177 N_A_79_21#_M1007_s N_A_c_530_n 0.00183785f $X=4.03 $Y=1.485 $X2=0 $Y2=0
cc_178 N_A_79_21#_c_166_p N_B_M1007_g 6.77174e-19 $X=3.53 $Y=1.85 $X2=0 $Y2=0
cc_179 N_A_79_21#_c_167_p N_B_M1007_g 0.00396717f $X=3.615 $Y=2.205 $X2=0 $Y2=0
cc_180 N_A_79_21#_c_175_p N_B_M1007_g 0.00836886f $X=4.165 $Y=2.29 $X2=0 $Y2=0
cc_181 N_A_79_21#_c_175_p N_B_M1032_g 0.00496191f $X=4.165 $Y=2.29 $X2=0 $Y2=0
cc_182 N_A_79_21#_c_166_p N_VPWR_M1016_s 0.00395387f $X=3.53 $Y=1.85 $X2=0 $Y2=0
cc_183 N_A_79_21#_M1005_g N_VPWR_c_792_n 0.0031902f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_184 N_A_79_21#_M1011_g N_VPWR_c_793_n 0.00146448f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_79_21#_M1022_g N_VPWR_c_793_n 0.00146448f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_79_21#_c_150_n N_VPWR_c_793_n 6.89403e-19 $X=1.805 $Y=1.16 $X2=0
+ $Y2=0
cc_187 N_A_79_21#_M1030_g N_VPWR_c_794_n 0.00330958f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_79_21#_c_151_n N_VPWR_c_794_n 0.0296352f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_79_21#_c_152_n N_VPWR_c_794_n 0.0123655f $X=2.225 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_79_21#_c_160_n N_VPWR_c_794_n 0.017295f $X=2.665 $Y=1.765 $X2=0 $Y2=0
cc_191 N_A_79_21#_c_162_p N_VPWR_c_794_n 0.0119226f $X=2.94 $Y=1.85 $X2=0 $Y2=0
cc_192 N_A_79_21#_c_166_p N_VPWR_c_795_n 0.0128626f $X=3.53 $Y=1.85 $X2=0 $Y2=0
cc_193 N_A_79_21#_c_167_p N_VPWR_c_795_n 0.00698652f $X=3.615 $Y=2.205 $X2=0
+ $Y2=0
cc_194 N_A_79_21#_c_191_p N_VPWR_c_795_n 0.0133617f $X=3.7 $Y=2.29 $X2=0 $Y2=0
cc_195 N_A_79_21#_M1005_g N_VPWR_c_804_n 0.00543342f $X=0.47 $Y=1.985 $X2=0
+ $Y2=0
cc_196 N_A_79_21#_M1011_g N_VPWR_c_804_n 0.00543342f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_197 N_A_79_21#_c_213_p N_VPWR_c_806_n 0.00644334f $X=2.855 $Y=2.19 $X2=0
+ $Y2=0
cc_198 N_A_79_21#_M1022_g N_VPWR_c_808_n 0.00543342f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_199 N_A_79_21#_M1030_g N_VPWR_c_808_n 0.00543342f $X=1.73 $Y=1.985 $X2=0
+ $Y2=0
cc_200 N_A_79_21#_c_191_p N_VPWR_c_809_n 0.00620913f $X=3.7 $Y=2.29 $X2=0 $Y2=0
cc_201 N_A_79_21#_c_175_p N_VPWR_c_809_n 0.022136f $X=4.165 $Y=2.29 $X2=0 $Y2=0
cc_202 N_A_79_21#_M1002_d N_VPWR_c_790_n 0.00284428f $X=2.72 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_A_79_21#_M1007_s N_VPWR_c_790_n 0.00224151f $X=4.03 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_79_21#_M1005_g N_VPWR_c_790_n 0.0104596f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_79_21#_M1011_g N_VPWR_c_790_n 0.00950542f $X=0.89 $Y=1.985 $X2=0
+ $Y2=0
cc_206 N_A_79_21#_M1022_g N_VPWR_c_790_n 0.00950542f $X=1.31 $Y=1.985 $X2=0
+ $Y2=0
cc_207 N_A_79_21#_M1030_g N_VPWR_c_790_n 0.0108315f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_208 N_A_79_21#_c_213_p N_VPWR_c_790_n 0.00599338f $X=2.855 $Y=2.19 $X2=0
+ $Y2=0
cc_209 N_A_79_21#_c_166_p N_VPWR_c_790_n 0.00604207f $X=3.53 $Y=1.85 $X2=0 $Y2=0
cc_210 N_A_79_21#_c_162_p N_VPWR_c_790_n 0.0137051f $X=2.94 $Y=1.85 $X2=0 $Y2=0
cc_211 N_A_79_21#_c_191_p N_VPWR_c_790_n 0.00595251f $X=3.7 $Y=2.29 $X2=0 $Y2=0
cc_212 N_A_79_21#_c_175_p N_VPWR_c_790_n 0.0211574f $X=4.165 $Y=2.29 $X2=0 $Y2=0
cc_213 N_A_79_21#_M1011_g N_SUM_c_936_n 0.00573279f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_79_21#_M1022_g N_SUM_c_936_n 0.0057349f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_215 N_A_79_21#_c_150_n N_SUM_c_936_n 0.0312791f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_79_21#_c_147_n N_SUM_c_941_n 4.88724e-19 $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_79_21#_c_148_n N_SUM_c_941_n 0.00390226f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_79_21#_c_149_n N_SUM_c_941_n 0.00409685f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_79_21#_c_148_n N_SUM_c_935_n 0.00333484f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_79_21#_c_149_n N_SUM_c_935_n 0.00277126f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_79_21#_c_150_n N_SUM_c_935_n 0.00778176f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_79_21#_M1022_g N_SUM_c_947_n 0.00743608f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_79_21#_M1030_g N_SUM_c_947_n 0.007823f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_79_21#_c_148_n N_SUM_c_949_n 0.00172083f $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_79_21#_c_149_n N_SUM_c_949_n 0.00322066f $X=1.73 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_79_21#_c_150_n N_SUM_c_949_n 6.39166e-19 $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_79_21#_M1030_g N_SUM_c_952_n 2.92808e-19 $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_228 N_A_79_21#_c_150_n N_SUM_c_952_n 0.0138241f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_79_21#_c_151_n N_SUM_c_952_n 0.0142213f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_79_21#_M1022_g N_SUM_c_955_n 0.00172083f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_231 N_A_79_21#_M1030_g N_SUM_c_955_n 0.0032678f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_232 N_A_79_21#_c_150_n N_SUM_c_955_n 6.18329e-19 $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_79_21#_M1011_g N_SUM_c_937_n 7.2991e-19 $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_234 N_A_79_21#_M1022_g N_SUM_c_937_n 0.00475337f $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_235 N_A_79_21#_M1030_g N_SUM_c_937_n 0.00390686f $X=1.73 $Y=1.985 $X2=0 $Y2=0
cc_236 N_A_79_21#_M1005_g SUM 5.32291e-19 $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_237 N_A_79_21#_c_150_n SUM 0.0219283f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_79_21#_M1005_g SUM 0.0191001f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_239 N_A_79_21#_M1011_g SUM 0.0145306f $X=0.89 $Y=1.985 $X2=0 $Y2=0
cc_240 N_A_79_21#_M1022_g SUM 7.28419e-19 $X=1.31 $Y=1.985 $X2=0 $Y2=0
cc_241 N_A_79_21#_c_146_n N_SUM_c_966_n 0.0126101f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_79_21#_c_147_n N_SUM_c_966_n 0.00941625f $X=0.89 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_79_21#_c_148_n N_SUM_c_966_n 4.87931e-19 $X=1.31 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_79_21#_c_150_n N_SUM_c_966_n 0.00877399f $X=1.805 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_79_21#_c_166_p A_717_297# 0.00208389f $X=3.53 $Y=1.85 $X2=-0.19
+ $Y2=-0.24
cc_246 N_A_79_21#_c_167_p A_717_297# 0.00282757f $X=3.615 $Y=2.205 $X2=-0.19
+ $Y2=-0.24
cc_247 N_A_79_21#_c_191_p A_717_297# 6.80208e-19 $X=3.7 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_79_21#_c_175_p A_717_297# 0.00382668f $X=4.165 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_79_21#_c_146_n N_VGND_c_1046_n 0.0031902f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_79_21#_c_147_n N_VGND_c_1047_n 0.00146448f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_79_21#_c_148_n N_VGND_c_1047_n 0.00146448f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_79_21#_c_150_n N_VGND_c_1047_n 0.00227153f $X=1.805 $Y=1.16 $X2=0
+ $Y2=0
cc_253 N_A_79_21#_c_149_n N_VGND_c_1048_n 0.00320738f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A_79_21#_c_151_n N_VGND_c_1048_n 0.0170433f $X=2.58 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_79_21#_c_152_n N_VGND_c_1048_n 0.00602806f $X=2.225 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_A_79_21#_c_146_n N_VGND_c_1057_n 0.00543728f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_79_21#_c_147_n N_VGND_c_1057_n 0.00543728f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_79_21#_c_148_n N_VGND_c_1065_n 0.00543728f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_79_21#_c_149_n N_VGND_c_1065_n 0.00543728f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_79_21#_M1015_s N_VGND_c_1071_n 0.00220248f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_79_21#_c_146_n N_VGND_c_1071_n 0.010461f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A_79_21#_c_147_n N_VGND_c_1071_n 0.00950676f $X=0.89 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_79_21#_c_148_n N_VGND_c_1071_n 0.00950676f $X=1.31 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_79_21#_c_149_n N_VGND_c_1071_n 0.0108328f $X=1.73 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_79_21#_M1015_s N_A_467_47#_c_1196_n 0.00319408f $X=2.745 $Y=0.235
+ $X2=0 $Y2=0
cc_266 N_A_79_21#_c_151_n N_A_467_47#_c_1196_n 0.00836099f $X=2.58 $Y=1.16 $X2=0
+ $Y2=0
cc_267 N_A_79_21#_c_152_n N_A_467_47#_c_1196_n 0.00158376f $X=2.225 $Y=1.16
+ $X2=0 $Y2=0
cc_268 N_A_79_21#_c_164_p N_A_467_47#_c_1196_n 0.0107372f $X=2.75 $Y=0.73 $X2=0
+ $Y2=0
cc_269 N_A_79_21#_c_169_p N_A_467_47#_c_1196_n 0.0126745f $X=2.88 $Y=0.73 $X2=0
+ $Y2=0
cc_270 N_A_514_199#_c_287_n N_A_c_506_n 0.024085f $X=3.09 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_271 N_A_514_199#_M1016_g N_A_M1026_g 0.038544f $X=3.065 $Y=1.985 $X2=0 $Y2=0
cc_272 N_A_514_199#_c_303_n N_A_M1026_g 5.55475e-19 $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_514_199#_c_304_n N_A_M1026_g 0.0106329f $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_274 N_A_514_199#_c_327_n N_A_M1028_g 0.0142369f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_275 N_A_514_199#_c_327_n N_A_M1029_g 0.0125968f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_276 N_A_514_199#_c_343_p N_A_c_508_n 4.64299e-19 $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_277 N_A_514_199#_c_288_n N_A_c_509_n 0.017632f $X=7.47 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_514_199#_c_345_p N_A_c_509_n 0.0116653f $X=7.225 $Y=0.73 $X2=0 $Y2=0
cc_279 N_A_514_199#_c_292_n N_A_c_509_n 0.00378439f $X=7.31 $Y=1.075 $X2=0 $Y2=0
cc_280 N_A_514_199#_M1008_g N_A_M1034_g 0.0266311f $X=7.47 $Y=1.985 $X2=0 $Y2=0
cc_281 N_A_514_199#_c_348_p N_A_M1034_g 0.0137749f $X=7.225 $Y=1.94 $X2=0 $Y2=0
cc_282 N_A_514_199#_c_293_n N_A_M1034_g 0.00684364f $X=7.31 $Y=1.855 $X2=0 $Y2=0
cc_283 N_A_514_199#_c_303_n N_A_c_510_n 0.0108194f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_514_199#_c_304_n N_A_c_510_n 0.0505135f $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_285 N_A_514_199#_c_327_n N_A_c_510_n 0.00370407f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_286 N_A_514_199#_c_295_n N_A_c_510_n 0.00130709f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_514_199#_c_303_n N_A_c_511_n 0.00113351f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_514_199#_c_304_n N_A_c_511_n 0.00293883f $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_289 N_A_514_199#_c_295_n N_A_c_511_n 0.0224357f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_290 N_A_514_199#_c_304_n N_A_c_520_n 0.0057125f $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_291 N_A_514_199#_c_327_n N_A_c_552_n 0.0703877f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_292 N_A_514_199#_c_327_n N_A_c_530_n 0.00822338f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_293 N_A_514_199#_c_327_n N_A_c_554_n 0.0109114f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_294 N_A_514_199#_M1029_d A 0.00753638f $X=5.785 $Y=1.485 $X2=0 $Y2=0
cc_295 N_A_514_199#_M1018_d A 2.26939e-19 $X=6.625 $Y=1.485 $X2=0 $Y2=0
cc_296 N_A_514_199#_c_363_p A 0.0273367f $X=6.675 $Y=1.94 $X2=0 $Y2=0
cc_297 N_A_514_199#_c_293_n A 0.00737137f $X=7.31 $Y=1.855 $X2=0 $Y2=0
cc_298 N_A_514_199#_c_365_p A 0.0118617f $X=5.92 $Y=1.94 $X2=0 $Y2=0
cc_299 N_A_514_199#_c_348_p N_A_c_513_n 8.68669e-19 $X=7.225 $Y=1.94 $X2=0 $Y2=0
cc_300 N_A_514_199#_c_345_p N_A_c_513_n 0.00125203f $X=7.225 $Y=0.73 $X2=0 $Y2=0
cc_301 N_A_514_199#_c_368_p N_A_c_513_n 8.10017e-19 $X=6.875 $Y=0.73 $X2=0 $Y2=0
cc_302 N_A_514_199#_c_292_n N_A_c_513_n 5.5452e-19 $X=7.31 $Y=1.075 $X2=0 $Y2=0
cc_303 N_A_514_199#_c_293_n N_A_c_513_n 5.5452e-19 $X=7.31 $Y=1.855 $X2=0 $Y2=0
cc_304 N_A_514_199#_c_294_n N_A_c_513_n 0.0013108f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_305 N_A_514_199#_c_296_n N_A_c_513_n 0.0131619f $X=8.73 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_514_199#_c_343_p N_A_c_514_n 0.00312548f $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_307 N_A_514_199#_c_348_p N_A_c_514_n 0.0051099f $X=7.225 $Y=1.94 $X2=0 $Y2=0
cc_308 N_A_514_199#_c_345_p N_A_c_514_n 0.0113072f $X=7.225 $Y=0.73 $X2=0 $Y2=0
cc_309 N_A_514_199#_c_368_p N_A_c_514_n 0.0121557f $X=6.875 $Y=0.73 $X2=0 $Y2=0
cc_310 N_A_514_199#_c_292_n N_A_c_514_n 0.00609836f $X=7.31 $Y=1.075 $X2=0 $Y2=0
cc_311 N_A_514_199#_c_293_n N_A_c_514_n 0.00609836f $X=7.31 $Y=1.855 $X2=0 $Y2=0
cc_312 N_A_514_199#_c_379_p N_A_c_514_n 0.00115591f $X=6.76 $Y=1.94 $X2=0 $Y2=0
cc_313 N_A_514_199#_c_294_n N_A_c_514_n 0.0147729f $X=7.31 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_514_199#_M1018_d N_A_c_575_n 0.00356052f $X=6.625 $Y=1.485 $X2=0
+ $Y2=0
cc_315 N_A_514_199#_c_363_p N_A_c_575_n 0.00306305f $X=6.675 $Y=1.94 $X2=0 $Y2=0
cc_316 N_A_514_199#_c_293_n N_A_c_575_n 0.00713541f $X=7.31 $Y=1.855 $X2=0 $Y2=0
cc_317 N_A_514_199#_c_379_p N_A_c_575_n 0.0102507f $X=6.76 $Y=1.94 $X2=0 $Y2=0
cc_318 N_A_514_199#_c_304_n N_B_M1007_g 0.00720076f $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_319 N_A_514_199#_c_386_p N_B_M1007_g 0.0052929f $X=3.955 $Y=1.855 $X2=0 $Y2=0
cc_320 N_A_514_199#_c_329_n N_B_M1007_g 0.00717689f $X=4.04 $Y=1.94 $X2=0 $Y2=0
cc_321 N_A_514_199#_c_304_n N_B_M1032_g 2.68247e-19 $X=3.87 $Y=1.51 $X2=0 $Y2=0
cc_322 N_A_514_199#_c_327_n N_B_M1032_g 0.012916f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_323 N_A_514_199#_c_343_p N_B_c_664_n 0.00346885f $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_324 N_A_514_199#_c_363_p N_B_M1003_g 0.0113283f $X=6.675 $Y=1.94 $X2=0 $Y2=0
cc_325 N_A_514_199#_c_343_p N_B_c_665_n 0.0112217f $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_326 N_A_514_199#_c_393_p N_B_c_665_n 0.00410088f $X=6.79 $Y=0.645 $X2=0 $Y2=0
cc_327 N_A_514_199#_c_368_p N_B_c_665_n 0.00213225f $X=6.875 $Y=0.73 $X2=0 $Y2=0
cc_328 N_A_514_199#_c_363_p N_B_M1018_g 0.0113124f $X=6.675 $Y=1.94 $X2=0 $Y2=0
cc_329 N_A_514_199#_c_327_n N_B_c_666_n 0.00157032f $X=5.835 $Y=1.94 $X2=0 $Y2=0
cc_330 N_A_514_199#_c_343_p N_B_c_671_n 0.00188491f $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_331 N_A_514_199#_M1000_d N_B_c_698_n 0.00267273f $X=6.205 $Y=0.235 $X2=0
+ $Y2=0
cc_332 N_A_514_199#_c_343_p N_B_c_698_n 0.00561594f $X=6.705 $Y=0.38 $X2=0 $Y2=0
cc_333 N_A_514_199#_c_368_p N_B_c_698_n 0.00778845f $X=6.875 $Y=0.73 $X2=0 $Y2=0
cc_334 N_A_514_199#_M1000_d B 7.05201e-19 $X=6.205 $Y=0.235 $X2=0 $Y2=0
cc_335 N_A_514_199#_c_304_n N_VPWR_M1016_s 0.00192876f $X=3.87 $Y=1.51 $X2=0
+ $Y2=0
cc_336 N_A_514_199#_c_327_n N_VPWR_M1028_d 0.00815262f $X=5.835 $Y=1.94 $X2=0
+ $Y2=0
cc_337 N_A_514_199#_c_363_p N_VPWR_M1003_s 0.0032492f $X=6.675 $Y=1.94 $X2=0
+ $Y2=0
cc_338 N_A_514_199#_c_348_p N_VPWR_M1034_s 0.00812625f $X=7.225 $Y=1.94 $X2=0
+ $Y2=0
cc_339 N_A_514_199#_c_293_n N_VPWR_M1034_s 0.00668051f $X=7.31 $Y=1.855 $X2=0
+ $Y2=0
cc_340 N_A_514_199#_M1002_g N_VPWR_c_794_n 0.026282f $X=2.645 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_514_199#_M1016_g N_VPWR_c_795_n 0.00281065f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_342 N_A_514_199#_c_327_n N_VPWR_c_796_n 0.0242313f $X=5.835 $Y=1.94 $X2=0
+ $Y2=0
cc_343 N_A_514_199#_c_327_n N_VPWR_c_797_n 0.00314825f $X=5.835 $Y=1.94 $X2=0
+ $Y2=0
cc_344 N_A_514_199#_c_411_p N_VPWR_c_797_n 0.00651665f $X=5.92 $Y=2.19 $X2=0
+ $Y2=0
cc_345 N_A_514_199#_c_363_p N_VPWR_c_797_n 0.00211912f $X=6.675 $Y=1.94 $X2=0
+ $Y2=0
cc_346 N_A_514_199#_c_363_p N_VPWR_c_798_n 0.0154434f $X=6.675 $Y=1.94 $X2=0
+ $Y2=0
cc_347 N_A_514_199#_c_363_p N_VPWR_c_799_n 0.00211912f $X=6.675 $Y=1.94 $X2=0
+ $Y2=0
cc_348 N_A_514_199#_c_415_p N_VPWR_c_799_n 0.00651665f $X=6.76 $Y=2.19 $X2=0
+ $Y2=0
cc_349 N_A_514_199#_c_348_p N_VPWR_c_799_n 0.00263154f $X=7.225 $Y=1.94 $X2=0
+ $Y2=0
cc_350 N_A_514_199#_M1008_g N_VPWR_c_800_n 0.00168836f $X=7.47 $Y=1.985 $X2=0
+ $Y2=0
cc_351 N_A_514_199#_c_348_p N_VPWR_c_800_n 0.0182311f $X=7.225 $Y=1.94 $X2=0
+ $Y2=0
cc_352 N_A_514_199#_M1008_g N_VPWR_c_801_n 7.80338e-19 $X=7.47 $Y=1.985 $X2=0
+ $Y2=0
cc_353 N_A_514_199#_M1019_g N_VPWR_c_801_n 0.0123546f $X=7.89 $Y=1.985 $X2=0
+ $Y2=0
cc_354 N_A_514_199#_M1027_g N_VPWR_c_801_n 0.00178624f $X=8.31 $Y=1.985 $X2=0
+ $Y2=0
cc_355 N_A_514_199#_M1035_g N_VPWR_c_803_n 0.00314466f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_356 N_A_514_199#_M1002_g N_VPWR_c_806_n 0.00585385f $X=2.645 $Y=1.985 $X2=0
+ $Y2=0
cc_357 N_A_514_199#_M1016_g N_VPWR_c_806_n 0.00585385f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_358 N_A_514_199#_c_327_n N_VPWR_c_809_n 0.0125021f $X=5.835 $Y=1.94 $X2=0
+ $Y2=0
cc_359 N_A_514_199#_M1008_g N_VPWR_c_810_n 0.00585385f $X=7.47 $Y=1.985 $X2=0
+ $Y2=0
cc_360 N_A_514_199#_M1019_g N_VPWR_c_810_n 0.0046653f $X=7.89 $Y=1.985 $X2=0
+ $Y2=0
cc_361 N_A_514_199#_M1027_g N_VPWR_c_811_n 0.00585385f $X=8.31 $Y=1.985 $X2=0
+ $Y2=0
cc_362 N_A_514_199#_M1035_g N_VPWR_c_811_n 0.00543342f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_363 N_A_514_199#_M1029_d N_VPWR_c_790_n 0.00268223f $X=5.785 $Y=1.485 $X2=0
+ $Y2=0
cc_364 N_A_514_199#_M1018_d N_VPWR_c_790_n 0.00268223f $X=6.625 $Y=1.485 $X2=0
+ $Y2=0
cc_365 N_A_514_199#_M1002_g N_VPWR_c_790_n 0.00792946f $X=2.645 $Y=1.985 $X2=0
+ $Y2=0
cc_366 N_A_514_199#_M1016_g N_VPWR_c_790_n 0.00621619f $X=3.065 $Y=1.985 $X2=0
+ $Y2=0
cc_367 N_A_514_199#_M1008_g N_VPWR_c_790_n 0.010724f $X=7.47 $Y=1.985 $X2=0
+ $Y2=0
cc_368 N_A_514_199#_M1019_g N_VPWR_c_790_n 0.00796766f $X=7.89 $Y=1.985 $X2=0
+ $Y2=0
cc_369 N_A_514_199#_M1027_g N_VPWR_c_790_n 0.0105126f $X=8.31 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_514_199#_M1035_g N_VPWR_c_790_n 0.0104987f $X=8.73 $Y=1.985 $X2=0
+ $Y2=0
cc_371 N_A_514_199#_c_327_n N_VPWR_c_790_n 0.0316145f $X=5.835 $Y=1.94 $X2=0
+ $Y2=0
cc_372 N_A_514_199#_c_411_p N_VPWR_c_790_n 0.00602802f $X=5.92 $Y=2.19 $X2=0
+ $Y2=0
cc_373 N_A_514_199#_c_363_p N_VPWR_c_790_n 0.00935238f $X=6.675 $Y=1.94 $X2=0
+ $Y2=0
cc_374 N_A_514_199#_c_415_p N_VPWR_c_790_n 0.00602802f $X=6.76 $Y=2.19 $X2=0
+ $Y2=0
cc_375 N_A_514_199#_c_348_p N_VPWR_c_790_n 0.00656324f $X=7.225 $Y=1.94 $X2=0
+ $Y2=0
cc_376 N_A_514_199#_c_304_n A_717_297# 0.00308682f $X=3.87 $Y=1.51 $X2=-0.19
+ $Y2=-0.24
cc_377 N_A_514_199#_c_327_n A_890_297# 0.0152665f $X=5.835 $Y=1.94 $X2=-0.19
+ $Y2=-0.24
cc_378 N_A_514_199#_c_289_n N_COUT_c_999_n 0.00654049f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_514_199#_c_290_n N_COUT_c_999_n 5.19831e-19 $X=8.31 $Y=0.995 $X2=0
+ $Y2=0
cc_380 N_A_514_199#_M1019_g N_COUT_c_996_n 0.012932f $X=7.89 $Y=1.985 $X2=0
+ $Y2=0
cc_381 N_A_514_199#_M1027_g N_COUT_c_996_n 0.0156389f $X=8.31 $Y=1.985 $X2=0
+ $Y2=0
cc_382 N_A_514_199#_c_449_p N_COUT_c_996_n 0.0323049f $X=8.06 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_514_199#_c_296_n N_COUT_c_996_n 0.00221825f $X=8.73 $Y=1.16 $X2=0
+ $Y2=0
cc_384 N_A_514_199#_M1008_g N_COUT_c_997_n 7.24989e-19 $X=7.47 $Y=1.985 $X2=0
+ $Y2=0
cc_385 N_A_514_199#_c_293_n N_COUT_c_997_n 0.00519059f $X=7.31 $Y=1.855 $X2=0
+ $Y2=0
cc_386 N_A_514_199#_c_449_p N_COUT_c_997_n 0.013717f $X=8.06 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A_514_199#_c_296_n N_COUT_c_997_n 0.00231083f $X=8.73 $Y=1.16 $X2=0
+ $Y2=0
cc_388 N_A_514_199#_c_289_n N_COUT_c_993_n 0.00850187f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_389 N_A_514_199#_c_290_n N_COUT_c_993_n 0.0133181f $X=8.31 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A_514_199#_c_449_p N_COUT_c_993_n 0.0266982f $X=8.06 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A_514_199#_c_296_n N_COUT_c_993_n 0.00221825f $X=8.73 $Y=1.16 $X2=0
+ $Y2=0
cc_392 N_A_514_199#_c_288_n N_COUT_c_994_n 6.63745e-19 $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_393 N_A_514_199#_c_289_n N_COUT_c_994_n 0.00211835f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_394 N_A_514_199#_c_292_n N_COUT_c_994_n 0.00142929f $X=7.31 $Y=1.075 $X2=0
+ $Y2=0
cc_395 N_A_514_199#_c_449_p N_COUT_c_994_n 0.0197956f $X=8.06 $Y=1.16 $X2=0
+ $Y2=0
cc_396 N_A_514_199#_c_296_n N_COUT_c_994_n 0.0022965f $X=8.73 $Y=1.16 $X2=0
+ $Y2=0
cc_397 N_A_514_199#_c_291_n COUT 0.00549581f $X=8.73 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A_514_199#_c_290_n COUT 0.00243005f $X=8.31 $Y=0.995 $X2=0 $Y2=0
cc_399 N_A_514_199#_M1027_g COUT 0.00243005f $X=8.31 $Y=1.985 $X2=0 $Y2=0
cc_400 N_A_514_199#_c_291_n COUT 0.00884511f $X=8.73 $Y=0.995 $X2=0 $Y2=0
cc_401 N_A_514_199#_M1035_g COUT 0.00460665f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_402 N_A_514_199#_c_449_p COUT 0.0126559f $X=8.06 $Y=1.16 $X2=0 $Y2=0
cc_403 N_A_514_199#_c_296_n COUT 0.0362993f $X=8.73 $Y=1.16 $X2=0 $Y2=0
cc_404 N_A_514_199#_M1035_g COUT 0.0167832f $X=8.73 $Y=1.985 $X2=0 $Y2=0
cc_405 N_A_514_199#_c_345_p N_VGND_M1033_s 0.00811624f $X=7.225 $Y=0.73 $X2=0
+ $Y2=0
cc_406 N_A_514_199#_c_292_n N_VGND_M1033_s 0.00119909f $X=7.31 $Y=1.075 $X2=0
+ $Y2=0
cc_407 N_A_514_199#_c_286_n N_VGND_c_1048_n 0.00728609f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_408 N_A_514_199#_c_287_n N_VGND_c_1049_n 0.001445f $X=3.09 $Y=0.995 $X2=0
+ $Y2=0
cc_409 N_A_514_199#_c_343_p N_VGND_c_1051_n 0.00597571f $X=6.705 $Y=0.38 $X2=0
+ $Y2=0
cc_410 N_A_514_199#_c_288_n N_VGND_c_1052_n 0.00179972f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_A_514_199#_c_345_p N_VGND_c_1052_n 0.0179903f $X=7.225 $Y=0.73 $X2=0
+ $Y2=0
cc_412 N_A_514_199#_c_288_n N_VGND_c_1053_n 0.00585385f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_413 N_A_514_199#_c_289_n N_VGND_c_1053_n 0.00426785f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_414 N_A_514_199#_c_289_n N_VGND_c_1054_n 0.0014456f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_415 N_A_514_199#_c_290_n N_VGND_c_1054_n 0.00160731f $X=8.31 $Y=0.995 $X2=0
+ $Y2=0
cc_416 N_A_514_199#_c_291_n N_VGND_c_1056_n 0.00314466f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_417 N_A_514_199#_c_286_n N_VGND_c_1059_n 0.00368123f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_418 N_A_514_199#_c_287_n N_VGND_c_1059_n 0.00368123f $X=3.09 $Y=0.995 $X2=0
+ $Y2=0
cc_419 N_A_514_199#_c_343_p N_VGND_c_1066_n 0.0310364f $X=6.705 $Y=0.38 $X2=0
+ $Y2=0
cc_420 N_A_514_199#_c_345_p N_VGND_c_1066_n 0.00267483f $X=7.225 $Y=0.73 $X2=0
+ $Y2=0
cc_421 N_A_514_199#_c_290_n N_VGND_c_1067_n 0.00439206f $X=8.31 $Y=0.995 $X2=0
+ $Y2=0
cc_422 N_A_514_199#_c_291_n N_VGND_c_1067_n 0.00543728f $X=8.73 $Y=0.995 $X2=0
+ $Y2=0
cc_423 N_A_514_199#_M1000_d N_VGND_c_1071_n 0.00217615f $X=6.205 $Y=0.235 $X2=0
+ $Y2=0
cc_424 N_A_514_199#_c_286_n N_VGND_c_1071_n 0.00657241f $X=2.67 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_A_514_199#_c_287_n N_VGND_c_1071_n 0.00531362f $X=3.09 $Y=0.995 $X2=0
+ $Y2=0
cc_426 N_A_514_199#_c_288_n N_VGND_c_1071_n 0.010724f $X=7.47 $Y=0.995 $X2=0
+ $Y2=0
cc_427 N_A_514_199#_c_289_n N_VGND_c_1071_n 0.00578036f $X=7.89 $Y=0.995 $X2=0
+ $Y2=0
cc_428 N_A_514_199#_c_290_n N_VGND_c_1071_n 0.00585554f $X=8.31 $Y=0.995 $X2=0
+ $Y2=0
cc_429 N_A_514_199#_c_291_n N_VGND_c_1071_n 0.0105f $X=8.73 $Y=0.995 $X2=0 $Y2=0
cc_430 N_A_514_199#_c_343_p N_VGND_c_1071_n 0.0246498f $X=6.705 $Y=0.38 $X2=0
+ $Y2=0
cc_431 N_A_514_199#_c_345_p N_VGND_c_1071_n 0.00610022f $X=7.225 $Y=0.73 $X2=0
+ $Y2=0
cc_432 N_A_514_199#_c_286_n N_A_467_47#_c_1196_n 0.0079064f $X=2.67 $Y=0.995
+ $X2=0 $Y2=0
cc_433 N_A_514_199#_c_287_n N_A_467_47#_c_1196_n 0.0108472f $X=3.09 $Y=0.995
+ $X2=0 $Y2=0
cc_434 N_A_514_199#_c_303_n N_A_467_47#_c_1196_n 0.00132561f $X=3.005 $Y=1.16
+ $X2=0 $Y2=0
cc_435 N_A_514_199#_c_304_n N_A_467_47#_c_1207_n 0.00324253f $X=3.87 $Y=1.51
+ $X2=0 $Y2=0
cc_436 N_A_514_199#_c_343_p A_1167_47# 0.00235165f $X=6.705 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_437 N_A_514_199#_c_393_p A_1167_47# 0.00197029f $X=6.79 $Y=0.645 $X2=-0.19
+ $Y2=-0.24
cc_438 N_A_514_199#_c_368_p A_1167_47# 0.00361316f $X=6.875 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_439 N_A_c_506_n N_B_c_662_n 0.0240792f $X=3.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_440 N_A_M1026_g N_B_M1007_g 0.0541861f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_441 N_A_c_520_n N_B_M1007_g 0.00227101f $X=4.295 $Y=1.505 $X2=0 $Y2=0
cc_442 N_A_c_530_n N_B_M1007_g 6.6402e-19 $X=4.38 $Y=1.59 $X2=0 $Y2=0
cc_443 N_A_M1028_g N_B_M1032_g 0.02761f $X=5.1 $Y=1.985 $X2=0 $Y2=0
cc_444 N_A_c_520_n N_B_M1032_g 0.00549698f $X=4.295 $Y=1.505 $X2=0 $Y2=0
cc_445 N_A_c_552_n N_B_M1032_g 0.00829481f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_446 N_A_c_530_n N_B_M1032_g 0.00340207f $X=4.38 $Y=1.59 $X2=0 $Y2=0
cc_447 N_A_c_508_n N_B_c_664_n 0.0527918f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_448 N_A_M1029_g N_B_M1003_g 0.0429883f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_449 N_A_c_521_n N_B_M1003_g 0.00299035f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_450 A N_B_M1003_g 0.0122437f $X=6.58 $Y=1.445 $X2=0 $Y2=0
cc_451 N_A_c_509_n N_B_c_665_n 0.0387678f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_452 N_A_M1034_g N_B_M1018_g 0.0412408f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_453 A N_B_M1018_g 0.0144706f $X=6.58 $Y=1.445 $X2=0 $Y2=0
cc_454 N_A_c_575_n N_B_M1018_g 0.00271894f $X=6.695 $Y=1.505 $X2=0 $Y2=0
cc_455 N_A_c_510_n N_B_c_666_n 0.0261808f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_456 N_A_c_511_n N_B_c_666_n 0.0206292f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_457 N_A_c_520_n N_B_c_666_n 0.00373275f $X=4.295 $Y=1.505 $X2=0 $Y2=0
cc_458 N_A_c_552_n N_B_c_667_n 0.0219781f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_459 N_A_c_512_n N_B_c_667_n 0.0141852f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_460 N_A_c_508_n N_B_c_723_n 0.0123223f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_461 N_A_c_521_n N_B_c_723_n 0.0108614f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_462 N_A_c_512_n N_B_c_723_n 0.00243363f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_463 N_A_c_510_n N_B_c_668_n 0.0129498f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_464 N_A_c_520_n N_B_c_668_n 0.00538854f $X=4.295 $Y=1.505 $X2=0 $Y2=0
cc_465 N_A_c_552_n N_B_c_668_n 0.0119252f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_466 N_A_c_512_n N_B_c_668_n 0.00108334f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_467 N_A_c_552_n N_B_c_669_n 0.00624449f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_468 N_A_c_512_n N_B_c_669_n 0.0167941f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_469 N_A_c_507_n N_B_c_670_n 0.0171894f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_470 N_A_c_508_n N_B_c_670_n 0.00150559f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_471 N_A_c_552_n N_B_c_670_n 0.0095326f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_472 N_A_c_521_n N_B_c_670_n 0.0129498f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_473 N_A_c_512_n N_B_c_670_n 0.00827575f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_474 N_A_c_521_n N_B_c_671_n 0.00120585f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_475 N_A_c_512_n N_B_c_671_n 0.0224296f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_476 A N_B_c_671_n 0.00277085f $X=6.58 $Y=1.445 $X2=0 $Y2=0
cc_477 N_A_c_513_n N_B_c_671_n 0.0214707f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_478 N_A_c_514_n N_B_c_671_n 0.0116639f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_c_508_n B 6.23642e-19 $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_480 N_A_c_521_n B 0.0149413f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_481 N_A_c_512_n B 0.00129606f $X=5.71 $Y=1.16 $X2=0 $Y2=0
cc_482 A B 0.0148377f $X=6.58 $Y=1.445 $X2=0 $Y2=0
cc_483 N_A_c_514_n B 0.0173528f $X=6.97 $Y=1.16 $X2=0 $Y2=0
cc_484 N_A_c_552_n N_VPWR_M1028_d 0.00985713f $X=5.625 $Y=1.59 $X2=0 $Y2=0
cc_485 A N_VPWR_M1003_s 0.00431279f $X=6.58 $Y=1.445 $X2=0 $Y2=0
cc_486 N_A_M1026_g N_VPWR_c_795_n 0.00546162f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_487 N_A_M1028_g N_VPWR_c_796_n 0.0110882f $X=5.1 $Y=1.985 $X2=0 $Y2=0
cc_488 N_A_M1029_g N_VPWR_c_796_n 0.00532324f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_489 N_A_M1029_g N_VPWR_c_797_n 0.00433717f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_490 N_A_M1029_g N_VPWR_c_798_n 8.41231e-19 $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_491 N_A_M1034_g N_VPWR_c_798_n 8.11451e-19 $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_492 N_A_M1034_g N_VPWR_c_799_n 0.00433717f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_493 N_A_M1034_g N_VPWR_c_800_n 0.00168836f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_494 N_A_M1026_g N_VPWR_c_809_n 0.00508534f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_495 N_A_M1028_g N_VPWR_c_809_n 0.00433717f $X=5.1 $Y=1.985 $X2=0 $Y2=0
cc_496 N_A_M1026_g N_VPWR_c_790_n 0.00602929f $X=3.51 $Y=1.985 $X2=0 $Y2=0
cc_497 N_A_M1028_g N_VPWR_c_790_n 0.00700833f $X=5.1 $Y=1.985 $X2=0 $Y2=0
cc_498 N_A_M1029_g N_VPWR_c_790_n 0.00640703f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_499 N_A_M1034_g N_VPWR_c_790_n 0.0059964f $X=6.97 $Y=1.985 $X2=0 $Y2=0
cc_500 N_A_c_552_n A_890_297# 0.0122997f $X=5.625 $Y=1.59 $X2=-0.19 $Y2=-0.24
cc_501 N_A_c_506_n N_VGND_c_1049_n 0.00834243f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_502 N_A_c_507_n N_VGND_c_1050_n 0.00164156f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_503 N_A_c_507_n N_VGND_c_1051_n 0.00723946f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_504 N_A_c_508_n N_VGND_c_1051_n 0.00914236f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_505 N_A_c_509_n N_VGND_c_1052_n 0.00323788f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_506 N_A_c_506_n N_VGND_c_1059_n 0.00340533f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_507 N_A_c_507_n N_VGND_c_1063_n 0.00365473f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_508 N_A_c_508_n N_VGND_c_1066_n 0.00341689f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_509 N_A_c_509_n N_VGND_c_1066_n 0.00426565f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_510 N_A_c_506_n N_VGND_c_1071_n 0.00403482f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_511 N_A_c_507_n N_VGND_c_1071_n 0.00597676f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_512 N_A_c_508_n N_VGND_c_1071_n 0.00392002f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_513 N_A_c_509_n N_VGND_c_1071_n 0.00587452f $X=6.97 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A_c_506_n N_A_467_47#_c_1208_n 0.0111056f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A_c_510_n N_A_467_47#_c_1208_n 0.0297332f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_516 N_A_c_511_n N_A_467_47#_c_1208_n 0.00121007f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_517 N_A_c_510_n N_A_467_47#_c_1207_n 0.00360822f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_518 N_A_c_511_n N_A_467_47#_c_1207_n 2.1253e-19 $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_519 N_A_c_510_n N_A_467_47#_c_1197_n 0.0057568f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_520 N_A_c_510_n N_A_467_47#_c_1214_n 0.00914406f $X=4.21 $Y=1.16 $X2=0 $Y2=0
cc_521 N_A_c_507_n N_A_467_47#_c_1198_n 0.00536239f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_522 N_B_M1003_g N_VPWR_c_797_n 0.00346207f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_523 N_B_M1003_g N_VPWR_c_798_n 0.0083298f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_524 N_B_M1018_g N_VPWR_c_798_n 0.00811325f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_525 N_B_M1018_g N_VPWR_c_799_n 0.00346207f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_526 N_B_M1007_g N_VPWR_c_809_n 0.00375986f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_527 N_B_M1032_g N_VPWR_c_809_n 0.00422171f $X=4.375 $Y=1.985 $X2=0 $Y2=0
cc_528 N_B_M1007_g N_VPWR_c_790_n 0.00537192f $X=3.955 $Y=1.985 $X2=0 $Y2=0
cc_529 N_B_M1032_g N_VPWR_c_790_n 0.00647341f $X=4.375 $Y=1.985 $X2=0 $Y2=0
cc_530 N_B_M1003_g N_VPWR_c_790_n 0.00413379f $X=6.13 $Y=1.985 $X2=0 $Y2=0
cc_531 N_B_M1018_g N_VPWR_c_790_n 0.00413379f $X=6.55 $Y=1.985 $X2=0 $Y2=0
cc_532 N_B_c_723_n N_VGND_M1024_d 0.00285509f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_533 N_B_c_670_n N_VGND_M1024_d 0.00245235f $X=5.41 $Y=0.74 $X2=0 $Y2=0
cc_534 N_B_c_662_n N_VGND_c_1049_n 0.00736307f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_535 N_B_c_663_n N_VGND_c_1049_n 7.22994e-19 $X=4.375 $Y=0.995 $X2=0 $Y2=0
cc_536 N_B_c_662_n N_VGND_c_1050_n 7.21572e-19 $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_537 N_B_c_663_n N_VGND_c_1050_n 0.00838542f $X=4.375 $Y=0.995 $X2=0 $Y2=0
cc_538 N_B_c_664_n N_VGND_c_1051_n 0.00188982f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_539 N_B_c_723_n N_VGND_c_1051_n 0.00827684f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_540 N_B_c_670_n N_VGND_c_1051_n 0.0064445f $X=5.41 $Y=0.74 $X2=0 $Y2=0
cc_541 N_B_c_662_n N_VGND_c_1061_n 0.00340533f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_542 N_B_c_663_n N_VGND_c_1061_n 0.00340533f $X=4.375 $Y=0.995 $X2=0 $Y2=0
cc_543 N_B_c_670_n N_VGND_c_1063_n 0.00156102f $X=5.41 $Y=0.74 $X2=0 $Y2=0
cc_544 N_B_c_664_n N_VGND_c_1066_n 0.00415552f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_545 N_B_c_665_n N_VGND_c_1066_n 0.00366111f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_546 N_B_c_723_n N_VGND_c_1066_n 0.00516314f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_547 N_B_c_698_n N_VGND_c_1066_n 0.00154365f $X=6.2 $Y=0.825 $X2=0 $Y2=0
cc_548 N_B_c_662_n N_VGND_c_1071_n 0.00400657f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_549 N_B_c_663_n N_VGND_c_1071_n 0.00400657f $X=4.375 $Y=0.995 $X2=0 $Y2=0
cc_550 N_B_c_664_n N_VGND_c_1071_n 0.0056496f $X=6.13 $Y=0.995 $X2=0 $Y2=0
cc_551 N_B_c_665_n N_VGND_c_1071_n 0.00526833f $X=6.55 $Y=0.995 $X2=0 $Y2=0
cc_552 N_B_c_723_n N_VGND_c_1071_n 0.0103908f $X=6.085 $Y=0.74 $X2=0 $Y2=0
cc_553 N_B_c_670_n N_VGND_c_1071_n 0.00307491f $X=5.41 $Y=0.74 $X2=0 $Y2=0
cc_554 N_B_c_698_n N_VGND_c_1071_n 0.00257233f $X=6.2 $Y=0.825 $X2=0 $Y2=0
cc_555 N_B_c_662_n N_A_467_47#_c_1208_n 0.0114147f $X=3.955 $Y=0.995 $X2=0 $Y2=0
cc_556 N_B_c_663_n N_A_467_47#_c_1197_n 0.0152279f $X=4.375 $Y=0.995 $X2=0 $Y2=0
cc_557 N_B_c_667_n N_A_467_47#_c_1197_n 0.0140675f $X=5.285 $Y=1.08 $X2=0 $Y2=0
cc_558 N_B_c_668_n N_A_467_47#_c_1197_n 0.0119373f $X=4.635 $Y=1.16 $X2=0 $Y2=0
cc_559 N_B_c_669_n N_A_467_47#_c_1197_n 0.0060788f $X=4.635 $Y=1.16 $X2=0 $Y2=0
cc_560 N_B_c_666_n N_A_467_47#_c_1214_n 0.0021626f $X=4.45 $Y=1.16 $X2=0 $Y2=0
cc_561 N_B_c_663_n N_A_467_47#_c_1198_n 0.00169479f $X=4.375 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_B_c_667_n N_A_467_47#_c_1198_n 0.018448f $X=5.285 $Y=1.08 $X2=0 $Y2=0
cc_563 N_B_c_670_n N_A_467_47#_c_1198_n 0.0129973f $X=5.41 $Y=0.74 $X2=0 $Y2=0
cc_564 N_B_c_723_n A_1325_47# 0.00593573f $X=6.085 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_565 N_VPWR_c_790_n N_SUM_M1005_d 0.00218509f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_566 N_VPWR_c_790_n N_SUM_M1022_d 0.00218509f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_567 N_VPWR_c_793_n N_SUM_c_936_n 0.0132514f $X=1.1 $Y=1.68 $X2=0 $Y2=0
cc_568 N_VPWR_c_808_n N_SUM_c_947_n 0.0143494f $X=1.855 $Y=2.72 $X2=0 $Y2=0
cc_569 N_VPWR_c_790_n N_SUM_c_947_n 0.0119017f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_570 N_VPWR_c_804_n SUM 0.0143494f $X=1.015 $Y=2.72 $X2=0 $Y2=0
cc_571 N_VPWR_c_790_n SUM 0.0119017f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_572 N_VPWR_c_790_n A_717_297# 0.00246661f $X=8.97 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_573 N_VPWR_c_790_n A_890_297# 0.00725566f $X=8.97 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_574 N_VPWR_c_790_n N_COUT_M1008_d 0.00572981f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_575 N_VPWR_c_790_n N_COUT_M1027_d 0.00292784f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_576 N_VPWR_c_810_n N_COUT_c_1028_n 0.00862177f $X=7.935 $Y=2.72 $X2=0 $Y2=0
cc_577 N_VPWR_c_790_n N_COUT_c_1028_n 0.00630811f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_578 N_VPWR_M1019_s N_COUT_c_996_n 0.00165831f $X=7.965 $Y=1.485 $X2=0 $Y2=0
cc_579 N_VPWR_c_801_n N_COUT_c_996_n 0.0148589f $X=8.1 $Y=1.92 $X2=0 $Y2=0
cc_580 N_VPWR_c_811_n COUT 0.0123106f $X=8.855 $Y=2.72 $X2=0 $Y2=0
cc_581 N_VPWR_c_790_n COUT 0.0102906f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_582 N_VPWR_c_792_n N_VGND_c_1046_n 0.00695811f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_583 N_VPWR_c_803_n N_VGND_c_1056_n 0.00695811f $X=8.94 $Y=1.66 $X2=0 $Y2=0
cc_584 N_SUM_c_936_n N_VGND_c_1047_n 0.0125734f $X=1.355 $Y=1.2 $X2=0 $Y2=0
cc_585 N_SUM_c_966_n N_VGND_c_1057_n 0.0136871f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_586 N_SUM_c_941_n N_VGND_c_1065_n 0.0136115f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_587 N_SUM_M1014_s N_VGND_c_1071_n 0.00219652f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_588 N_SUM_M1021_s N_VGND_c_1071_n 0.00219652f $X=1.385 $Y=0.235 $X2=0 $Y2=0
cc_589 N_SUM_c_941_n N_VGND_c_1071_n 0.01179f $X=1.52 $Y=0.4 $X2=0 $Y2=0
cc_590 N_SUM_c_966_n N_VGND_c_1071_n 0.0118335f $X=0.68 $Y=0.4 $X2=0 $Y2=0
cc_591 N_COUT_c_993_n N_VGND_M1004_d 0.00162006f $X=8.405 $Y=0.82 $X2=0 $Y2=0
cc_592 N_COUT_c_999_n N_VGND_c_1053_n 0.0108823f $X=7.68 $Y=0.57 $X2=0 $Y2=0
cc_593 N_COUT_c_993_n N_VGND_c_1053_n 0.00193763f $X=8.405 $Y=0.82 $X2=0 $Y2=0
cc_594 N_COUT_c_993_n N_VGND_c_1054_n 0.0122414f $X=8.405 $Y=0.82 $X2=0 $Y2=0
cc_595 N_COUT_c_993_n N_VGND_c_1067_n 0.0021796f $X=8.405 $Y=0.82 $X2=0 $Y2=0
cc_596 COUT N_VGND_c_1067_n 0.0117653f $X=8.42 $Y=0.425 $X2=0 $Y2=0
cc_597 N_COUT_M1001_s N_VGND_c_1071_n 0.00397494f $X=7.545 $Y=0.235 $X2=0 $Y2=0
cc_598 N_COUT_M1010_s N_VGND_c_1071_n 0.0023038f $X=8.385 $Y=0.235 $X2=0 $Y2=0
cc_599 N_COUT_c_999_n N_VGND_c_1071_n 0.00908244f $X=7.68 $Y=0.57 $X2=0 $Y2=0
cc_600 N_COUT_c_993_n N_VGND_c_1071_n 0.00850926f $X=8.405 $Y=0.82 $X2=0 $Y2=0
cc_601 COUT N_VGND_c_1071_n 0.0102437f $X=8.42 $Y=0.425 $X2=0 $Y2=0
cc_602 N_VGND_c_1071_n N_A_467_47#_M1015_d 0.0021262f $X=8.97 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_603 N_VGND_c_1071_n N_A_467_47#_M1017_d 0.00238507f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1071_n N_A_467_47#_M1023_s 0.00258634f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_605 N_VGND_c_1071_n N_A_467_47#_M1024_s 0.0048671f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_1048_n N_A_467_47#_c_1196_n 0.0142345f $X=1.94 $Y=0.38 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1059_n N_A_467_47#_c_1196_n 0.0489351f $X=3.555 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1071_n N_A_467_47#_c_1196_n 0.038975f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_609 N_VGND_M1013_d N_A_467_47#_c_1208_n 0.00419315f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1049_n N_A_467_47#_c_1208_n 0.0170265f $X=3.73 $Y=0.38 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1059_n N_A_467_47#_c_1208_n 0.00237932f $X=3.555 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1061_n N_A_467_47#_c_1208_n 0.00237932f $X=4.42 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1071_n N_A_467_47#_c_1208_n 0.00994979f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_c_1061_n N_A_467_47#_c_1237_n 0.00702781f $X=4.42 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_1071_n N_A_467_47#_c_1237_n 0.00609156f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_M1025_d N_A_467_47#_c_1197_n 0.00474739f $X=4.45 $Y=0.235 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1050_n N_A_467_47#_c_1197_n 0.0196494f $X=4.585 $Y=0.38 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1061_n N_A_467_47#_c_1197_n 0.00237932f $X=4.42 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1063_n N_A_467_47#_c_1197_n 0.00302409f $X=5.385 $Y=0 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1071_n N_A_467_47#_c_1197_n 0.0104658f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_1050_n N_A_467_47#_c_1198_n 0.0173063f $X=4.585 $Y=0.38 $X2=0
+ $Y2=0
cc_622 N_VGND_c_1051_n N_A_467_47#_c_1198_n 0.0145071f $X=5.55 $Y=0.38 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1063_n N_A_467_47#_c_1198_n 0.0186073f $X=5.385 $Y=0 $X2=0 $Y2=0
cc_624 N_VGND_c_1071_n N_A_467_47#_c_1198_n 0.010309f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_1071_n A_1325_47# 0.00263295f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24
cc_626 N_VGND_c_1071_n A_1167_47# 0.00226587f $X=8.97 $Y=0 $X2=-0.19 $Y2=-0.24

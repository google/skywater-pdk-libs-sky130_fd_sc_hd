* File: sky130_fd_sc_hd__and4bb_4.pex.spice
* Created: Tue Sep  1 18:58:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__AND4BB_4%B_N 3 7 9 10 11 16
c34 7 0 1.74445e-19 $X=0.47 $Y=2.275
c35 3 0 1.38832e-19 $X=0.47 $Y=0.445
r36 16 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=1.325
r37 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.515 $Y2=0.995
r38 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r39 10 11 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.53
r40 10 17 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=0.605 $Y=1.19
+ $X2=0.605 $Y2=1.16
r41 9 17 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.605 $Y=0.85
+ $X2=0.605 $Y2=1.16
r42 7 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.47 $Y=2.275
+ $X2=0.47 $Y2=1.325
r43 3 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.47 $Y=0.445
+ $X2=0.47 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%A_174_21# 1 2 3 12 14 16 19 21 23 26 28 30
+ 33 35 37 38 47 49 50 51 52 56 59 60 61 62 71
r144 70 71 59.193 $w=3.42e-07 $l=4.2e-07 $layer=POLY_cond $X=1.785 $Y=1.2
+ $X2=2.205 $Y2=1.2
r145 67 68 59.193 $w=3.42e-07 $l=4.2e-07 $layer=POLY_cond $X=0.945 $Y=1.2
+ $X2=1.365 $Y2=1.2
r146 60 61 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=4.255 $Y=0.385
+ $X2=2.94 $Y2=0.385
r147 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.855 $Y=0.47
+ $X2=2.94 $Y2=0.385
r148 58 59 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.855 $Y=0.47
+ $X2=2.855 $Y2=0.615
r149 54 56 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.975 $Y=1.63
+ $X2=3.985 $Y2=1.63
r150 52 54 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.5 $Y=1.63
+ $X2=2.975 $Y2=1.63
r151 50 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=0.7
+ $X2=2.855 $Y2=0.615
r152 50 51 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.77 $Y=0.7 $X2=2.5
+ $Y2=0.7
r153 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=1.545
+ $X2=2.5 $Y2=1.63
r154 48 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=1.245
+ $X2=2.415 $Y2=1.16
r155 48 49 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.415 $Y=1.245
+ $X2=2.415 $Y2=1.545
r156 47 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=1.075
+ $X2=2.415 $Y2=1.16
r157 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=0.785
+ $X2=2.5 $Y2=0.7
r158 46 47 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.415 $Y=0.785
+ $X2=2.415 $Y2=1.075
r159 45 71 7.04678 $w=3.42e-07 $l=5e-08 $layer=POLY_cond $X=2.255 $Y=1.2
+ $X2=2.205 $Y2=1.2
r160 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=1.16 $X2=2.255 $Y2=1.16
r161 41 70 29.5965 $w=3.42e-07 $l=2.1e-07 $layer=POLY_cond $X=1.575 $Y=1.2
+ $X2=1.785 $Y2=1.2
r162 41 68 29.5965 $w=3.42e-07 $l=2.1e-07 $layer=POLY_cond $X=1.575 $Y=1.2
+ $X2=1.365 $Y2=1.2
r163 40 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.575 $Y=1.16
+ $X2=2.255 $Y2=1.16
r164 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.16 $X2=1.575 $Y2=1.16
r165 38 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.33 $Y=1.16
+ $X2=2.415 $Y2=1.16
r166 38 44 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.33 $Y=1.16
+ $X2=2.255 $Y2=1.16
r167 35 71 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.205 $Y=1.375
+ $X2=2.205 $Y2=1.2
r168 35 37 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.205 $Y=1.375
+ $X2=2.205 $Y2=1.985
r169 31 71 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.205 $Y=1.025
+ $X2=2.205 $Y2=1.2
r170 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.205 $Y=1.025
+ $X2=2.205 $Y2=0.56
r171 28 70 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.785 $Y=1.375
+ $X2=1.785 $Y2=1.2
r172 28 30 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.785 $Y=1.375
+ $X2=1.785 $Y2=1.985
r173 24 70 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.785 $Y=1.025
+ $X2=1.785 $Y2=1.2
r174 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.785 $Y=1.025
+ $X2=1.785 $Y2=0.56
r175 21 68 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.365 $Y=1.375
+ $X2=1.365 $Y2=1.2
r176 21 23 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.365 $Y=1.375
+ $X2=1.365 $Y2=1.985
r177 17 68 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.365 $Y=1.025
+ $X2=1.365 $Y2=1.2
r178 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.365 $Y=1.025
+ $X2=1.365 $Y2=0.56
r179 14 67 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.945 $Y=1.375
+ $X2=0.945 $Y2=1.2
r180 14 16 196.013 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.945 $Y=1.375
+ $X2=0.945 $Y2=1.985
r181 10 67 22.0749 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=1.2
r182 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.945 $Y=1.025
+ $X2=0.945 $Y2=0.56
r183 3 56 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.485 $X2=3.985 $Y2=1.63
r184 2 54 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.485 $X2=2.975 $Y2=1.63
r185 1 60 91 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.235 $X2=4.445 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%D 3 6 8 11 13
c39 6 0 1.1816e-19 $X=2.705 $Y=1.985
r40 11 14 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.16
+ $X2=2.765 $Y2=1.325
r41 11 13 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.16
+ $X2=2.765 $Y2=0.995
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.16 $X2=2.765 $Y2=1.16
r43 8 12 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=2.765 $Y2=1.16
r44 6 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.705 $Y=1.985
+ $X2=2.705 $Y2=1.325
r45 3 13 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.705 $Y=0.56
+ $X2=2.705 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%C 3 6 8 9 13 15
r35 13 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.29 $Y=1.16
+ $X2=3.29 $Y2=1.325
r36 13 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.29 $Y=1.16
+ $X2=3.29 $Y2=0.995
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.335
+ $Y=1.16 $X2=3.335 $Y2=1.16
r38 9 14 1.17198 $w=2.93e-07 $l=3e-08 $layer=LI1_cond $X=3.397 $Y=1.19 $X2=3.397
+ $Y2=1.16
r39 8 14 12.1104 $w=2.93e-07 $l=3.1e-07 $layer=LI1_cond $X=3.397 $Y=0.85
+ $X2=3.397 $Y2=1.16
r40 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.185 $Y=1.985
+ $X2=3.185 $Y2=1.325
r41 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.185 $Y=0.56
+ $X2=3.185 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%A_27_47# 1 2 9 12 15 18 20 22 25 27 30 32
+ 33 37
r91 33 38 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.16
+ $X2=3.815 $Y2=1.325
r92 33 37 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.16
+ $X2=3.815 $Y2=0.995
r93 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.16 $X2=3.815 $Y2=1.16
r94 27 29 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.42
+ $X2=0.215 $Y2=0.585
r95 24 25 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.405 $Y=1.325
+ $X2=4.405 $Y2=1.915
r96 23 32 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.9 $Y=1.24
+ $X2=3.815 $Y2=1.16
r97 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.32 $Y=1.24
+ $X2=4.405 $Y2=1.325
r98 22 23 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.32 $Y=1.24 $X2=3.9
+ $Y2=1.24
r99 21 30 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.215
+ $Y2=2
r100 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.32 $Y=2
+ $X2=4.405 $Y2=1.915
r101 20 21 259.332 $w=1.68e-07 $l=3.975e-06 $layer=LI1_cond $X=4.32 $Y=2
+ $X2=0.345 $Y2=2
r102 16 30 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2
r103 16 18 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2.3
r104 15 30 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.215 $Y2=2
r105 15 29 84.2909 $w=1.73e-07 $l=1.33e-06 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.172 $Y2=0.585
r106 12 38 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.755 $Y=1.985
+ $X2=3.755 $Y2=1.325
r107 9 37 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.755 $Y=0.56
+ $X2=3.755 $Y2=0.995
r108 2 18 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r109 1 27 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%A_832_21# 1 2 7 9 12 15 19 20 21 22 23 24
+ 27 31
r65 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.72 $Y=2.085
+ $X2=5.72 $Y2=2.3
r66 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.72 $Y=0.655
+ $X2=5.72 $Y2=0.42
r67 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.635 $Y=2
+ $X2=5.72 $Y2=2.085
r68 23 24 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.635 $Y=2 $X2=5.12
+ $Y2=2
r69 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.635 $Y=0.74
+ $X2=5.72 $Y2=0.655
r70 21 22 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.635 $Y=0.74
+ $X2=5.12 $Y2=0.74
r71 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.035
+ $Y=1.16 $X2=5.035 $Y2=1.16
r72 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=1.915
+ $X2=5.12 $Y2=2
r73 17 19 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=5.035 $Y=1.915
+ $X2=5.035 $Y2=1.16
r74 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=0.825
+ $X2=5.12 $Y2=0.74
r75 16 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.035 $Y=0.825
+ $X2=5.035 $Y2=1.16
r76 14 20 126.774 $w=3.3e-07 $l=7.25e-07 $layer=POLY_cond $X=4.31 $Y=1.16
+ $X2=5.035 $Y2=1.16
r77 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.31 $Y=1.16
+ $X2=4.235 $Y2=1.16
r78 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=1.16
r79 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=1.985
r80 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=0.995
+ $X2=4.235 $Y2=1.16
r81 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.235 $Y=0.995
+ $X2=4.235 $Y2=0.56
r82 2 31 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=2.065 $X2=5.72 $Y2=2.3
r83 1 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.585
+ $Y=0.235 $X2=5.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%A_N 3 7 9 10 14 15
r24 14 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.57 $Y=1.16
+ $X2=5.57 $Y2=1.325
r25 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.57 $Y=1.16
+ $X2=5.57 $Y2=0.995
r26 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.16 $X2=5.57 $Y2=1.16
r27 9 10 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=5.665 $Y=1.19
+ $X2=5.665 $Y2=1.53
r28 9 15 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=5.665 $Y=1.19
+ $X2=5.665 $Y2=1.16
r29 7 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.51 $Y=2.275
+ $X2=5.51 $Y2=1.325
r30 3 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.51 $Y=0.445
+ $X2=5.51 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%VPWR 1 2 3 4 5 18 22 26 30 34 35 37 38 39
+ 41 46 55 61 62 65 68 71 76 84
r92 82 84 7.9835 $w=5.48e-07 $l=8e-08 $layer=LI1_cond $X=5.29 $Y=2.53 $X2=5.37
+ $Y2=2.53
r93 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r94 80 82 1.84848 $w=5.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.53
+ $X2=5.29 $Y2=2.53
r95 75 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r96 74 78 3.37077 $w=5.48e-07 $l=1.55e-07 $layer=LI1_cond $X=4.37 $Y=2.53
+ $X2=4.525 $Y2=2.53
r97 74 76 6.46121 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=4.37 $Y=2.53 $X2=4.36
+ $Y2=2.53
r98 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r99 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r102 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r103 62 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r104 61 84 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=5.37 $Y2=2.72
r105 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 58 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r108 55 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.495 $Y2=2.72
r109 55 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=2.99 $Y2=2.72
r110 54 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r111 54 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=1.575 $Y2=2.72
r114 51 53 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.72
+ $X2=2.07 $Y2=2.72
r115 50 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r116 50 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r119 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 46 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.575 $Y2=2.72
r121 46 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.15 $Y2=2.72
r122 41 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r123 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 39 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 37 53 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=2.72
+ $X2=2.415 $Y2=2.72
r128 36 57 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=2.99 $Y2=2.72
r129 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=2.72
+ $X2=2.415 $Y2=2.72
r130 35 78 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=4.635 $Y=2.53
+ $X2=4.525 $Y2=2.53
r131 34 80 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.095 $Y=2.53
+ $X2=5.205 $Y2=2.53
r132 34 35 10.0036 $w=5.48e-07 $l=4.6e-07 $layer=LI1_cond $X=5.095 $Y=2.53
+ $X2=4.635 $Y2=2.53
r133 33 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=2.72
+ $X2=3.495 $Y2=2.72
r134 33 76 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.66 $Y=2.72 $X2=4.36
+ $Y2=2.72
r135 28 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.635
+ $X2=3.495 $Y2=2.72
r136 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=2.635
+ $X2=3.495 $Y2=2.34
r137 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.72
r138 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.415 $Y=2.635
+ $X2=2.415 $Y2=2.34
r139 20 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.72
r140 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.575 $Y=2.635
+ $X2=1.575 $Y2=2.34
r141 16 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r142 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.34
r143 5 80 400 $w=1.7e-07 $l=1.2515e-06 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.485 $X2=5.205 $Y2=2.34
r144 5 78 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=1.485 $X2=4.525 $Y2=2.34
r145 4 30 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.485 $X2=3.495 $Y2=2.34
r146 3 26 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.485 $X2=2.415 $Y2=2.34
r147 2 22 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=1.485 $X2=1.575 $Y2=2.34
r148 1 18 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=2.065 $X2=0.68 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%X 1 2 3 4 15 19 21 22 23 24 33 35 41 46
c45 46 0 1.1816e-19 $X=1.995 $Y=1.63
c46 35 0 3.13277e-19 $X=1.155 $Y=0.85
r47 33 41 0.61738 $w=2.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.1 $Y=1.545 $X2=1.1
+ $Y2=1.53
r48 32 35 1.23476 $w=2.78e-07 $l=3e-08 $layer=LI1_cond $X=1.1 $Y=0.82 $X2=1.1
+ $Y2=0.85
r49 24 33 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=1.63 $X2=1.1
+ $Y2=1.545
r50 24 46 37.2497 $w=2.38e-07 $l=7.55e-07 $layer=LI1_cond $X=1.24 $Y=1.63
+ $X2=1.995 $Y2=1.63
r51 24 41 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=1.1 $Y=1.495 $X2=1.1
+ $Y2=1.53
r52 23 24 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.1 $Y=1.19 $X2=1.1
+ $Y2=1.495
r53 22 32 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.735 $X2=1.1
+ $Y2=0.82
r54 22 23 12.8827 $w=2.78e-07 $l=3.13e-07 $layer=LI1_cond $X=1.1 $Y=0.877
+ $X2=1.1 $Y2=1.19
r55 22 35 1.11128 $w=2.78e-07 $l=2.7e-08 $layer=LI1_cond $X=1.1 $Y=0.877 $X2=1.1
+ $Y2=0.85
r56 21 22 35.0328 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=1.91 $Y=0.735
+ $X2=1.24 $Y2=0.735
r57 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.995 $Y=0.65
+ $X2=1.91 $Y2=0.735
r58 17 19 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.995 $Y=0.65
+ $X2=1.995 $Y2=0.42
r59 13 22 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=1.155 $Y=0.65
+ $X2=1.1 $Y2=0.735
r60 13 15 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.155 $Y=0.65
+ $X2=1.155 $Y2=0.42
r61 4 46 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.485 $X2=1.995 $Y2=1.63
r62 3 24 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.485 $X2=1.155 $Y2=1.63
r63 2 19 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=1.995 $Y2=0.42
r64 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HD__AND4BB_4%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 54 55 58 61 64
r96 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r97 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r98 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r99 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r100 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r101 52 65 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=2.53
+ $Y2=0
r102 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r103 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.435
+ $Y2=0
r104 49 51 145.487 $w=1.68e-07 $l=2.23e-06 $layer=LI1_cond $X=2.6 $Y=0 $X2=4.83
+ $Y2=0
r105 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r106 48 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r107 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r108 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.575
+ $Y2=0
r109 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=2.07
+ $Y2=0
r110 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.435
+ $Y2=0
r111 44 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.07
+ $Y2=0
r112 43 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r113 43 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r114 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r115 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.735
+ $Y2=0
r116 40 42 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.15
+ $Y2=0
r117 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.575
+ $Y2=0
r118 39 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.15
+ $Y2=0
r119 34 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.735
+ $Y2=0
r120 34 36 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.23
+ $Y2=0
r121 32 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r122 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r123 30 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.83 $Y2=0
r124 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=5.14
+ $Y2=0
r125 29 54 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.305 $Y=0
+ $X2=5.75 $Y2=0
r126 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.305 $Y=0 $X2=5.14
+ $Y2=0
r127 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.085
+ $X2=5.14 $Y2=0
r128 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.14 $Y=0.085
+ $X2=5.14 $Y2=0.38
r129 21 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0
r130 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=0.085
+ $X2=2.435 $Y2=0.36
r131 17 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0
r132 17 19 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.575 $Y=0.085
+ $X2=1.575 $Y2=0.385
r133 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r134 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.38
r135 4 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.235 $X2=5.14 $Y2=0.38
r136 3 23 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.28
+ $Y=0.235 $X2=2.435 $Y2=0.36
r137 2 19 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.575 $Y2=0.385
r138 1 15 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.735 $Y2=0.38
.ends


* File: sky130_fd_sc_hd__o211ai_2.pxi.spice
* Created: Thu Aug 27 14:34:55 2020
* 
x_PM_SKY130_FD_SC_HD__O211AI_2%C1 N_C1_c_64_n N_C1_M1004_g N_C1_M1002_g
+ N_C1_c_65_n N_C1_M1006_g N_C1_M1009_g C1 N_C1_c_66_n N_C1_c_67_n
+ PM_SKY130_FD_SC_HD__O211AI_2%C1
x_PM_SKY130_FD_SC_HD__O211AI_2%B1 N_B1_c_105_n N_B1_M1001_g N_B1_M1005_g
+ N_B1_c_106_n N_B1_M1013_g N_B1_M1014_g B1 N_B1_c_108_n
+ PM_SKY130_FD_SC_HD__O211AI_2%B1
x_PM_SKY130_FD_SC_HD__O211AI_2%A2 N_A2_c_152_n N_A2_M1003_g N_A2_M1000_g
+ N_A2_c_153_n N_A2_M1010_g N_A2_M1007_g A2 N_A2_c_154_n N_A2_c_155_n
+ PM_SKY130_FD_SC_HD__O211AI_2%A2
x_PM_SKY130_FD_SC_HD__O211AI_2%A1 N_A1_c_195_n N_A1_M1008_g N_A1_M1011_g
+ N_A1_c_196_n N_A1_M1012_g N_A1_M1015_g A1 N_A1_c_197_n A1
+ PM_SKY130_FD_SC_HD__O211AI_2%A1
x_PM_SKY130_FD_SC_HD__O211AI_2%VPWR N_VPWR_M1002_s N_VPWR_M1009_s N_VPWR_M1014_s
+ N_VPWR_M1011_d N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n
+ N_VPWR_c_239_n VPWR N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n
+ N_VPWR_c_243_n N_VPWR_c_234_n N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n
+ PM_SKY130_FD_SC_HD__O211AI_2%VPWR
x_PM_SKY130_FD_SC_HD__O211AI_2%Y N_Y_M1004_s N_Y_M1002_d N_Y_M1005_d N_Y_M1000_s
+ N_Y_c_304_n N_Y_c_305_n N_Y_c_338_n N_Y_c_303_n N_Y_c_306_n N_Y_c_319_n
+ N_Y_c_327_n Y N_Y_c_308_n PM_SKY130_FD_SC_HD__O211AI_2%Y
x_PM_SKY130_FD_SC_HD__O211AI_2%A_487_297# N_A_487_297#_M1000_d
+ N_A_487_297#_M1007_d N_A_487_297#_M1015_s N_A_487_297#_c_355_n
+ N_A_487_297#_c_352_n N_A_487_297#_c_353_n N_A_487_297#_c_354_n
+ PM_SKY130_FD_SC_HD__O211AI_2%A_487_297#
x_PM_SKY130_FD_SC_HD__O211AI_2%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1006_d
+ N_A_27_47#_M1013_d N_A_27_47#_c_378_n N_A_27_47#_c_379_n N_A_27_47#_c_380_n
+ N_A_27_47#_c_399_p PM_SKY130_FD_SC_HD__O211AI_2%A_27_47#
x_PM_SKY130_FD_SC_HD__O211AI_2%A_286_47# N_A_286_47#_M1001_s N_A_286_47#_M1003_s
+ N_A_286_47#_M1008_d N_A_286_47#_c_406_n N_A_286_47#_c_417_n
+ PM_SKY130_FD_SC_HD__O211AI_2%A_286_47#
x_PM_SKY130_FD_SC_HD__O211AI_2%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_M1012_s
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ N_VGND_c_444_n PM_SKY130_FD_SC_HD__O211AI_2%VGND
cc_1 VNB N_C1_c_64_n 0.0215565f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB N_C1_c_65_n 0.0159703f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.995
cc_3 VNB N_C1_c_66_n 0.0161079f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_4 VNB N_C1_c_67_n 0.0555515f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.16
cc_5 VNB N_B1_c_105_n 0.0164337f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_6 VNB N_B1_c_106_n 0.0220812f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.995
cc_7 VNB B1 0.00665371f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_8 VNB N_B1_c_108_n 0.0404119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A2_c_152_n 0.0212151f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_10 VNB N_A2_c_153_n 0.016201f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.995
cc_11 VNB N_A2_c_154_n 0.00893908f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_12 VNB N_A2_c_155_n 0.0381109f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.16
cc_13 VNB N_A1_c_195_n 0.016193f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_14 VNB N_A1_c_196_n 0.0191729f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.995
cc_15 VNB N_A1_c_197_n 0.0366801f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.16
cc_16 VNB A1 0.0282418f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.53
cc_17 VNB N_VPWR_c_234_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_378_n 0.00871655f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_19 VNB N_A_27_47#_c_379_n 0.00176237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_380_n 0.00233548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_286_47#_c_406_n 0.0136538f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=0.56
cc_22 VNB N_VGND_c_435_n 0.00491914f $X=-0.19 $Y=-0.24 $X2=0.925 $Y2=1.985
cc_23 VNB N_VGND_c_436_n 3.0911e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_437_n 0.0122109f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_25 VNB N_VGND_c_438_n 0.0108354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_439_n 0.0573682f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_27 VNB N_VGND_c_440_n 0.0123625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_441_n 0.0128832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_442_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_443_n 0.00436029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_444_n 0.242651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_C1_M1002_g 0.0213135f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_33 VPB N_C1_M1009_g 0.0181347f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_34 VPB N_C1_c_66_n 0.0273104f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_35 VPB N_C1_c_67_n 0.0157052f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.16
cc_36 VPB N_B1_M1005_g 0.0184395f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_37 VPB N_B1_M1014_g 0.0243789f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_38 VPB B1 0.00669577f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_39 VPB N_B1_c_108_n 0.00701377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A2_M1000_g 0.0254715f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_41 VPB N_A2_M1007_g 0.0187919f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_42 VPB N_A2_c_154_n 0.0089665f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_43 VPB N_A2_c_155_n 0.00580464f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.16
cc_44 VPB N_A1_M1011_g 0.0188665f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_45 VPB N_A1_M1015_g 0.0259057f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_46 VPB N_A1_c_197_n 0.00593495f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.16
cc_47 VPB N_VPWR_c_235_n 0.0107363f $X=-0.19 $Y=1.305 $X2=0.925 $Y2=1.985
cc_48 VPB N_VPWR_c_236_n 0.0165287f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_49 VPB N_VPWR_c_237_n 3.20903e-19 $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_50 VPB N_VPWR_c_238_n 0.00951479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_239_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_240_n 0.0154314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_241_n 0.0129398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_242_n 0.0364632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_243_n 0.0172852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_234_n 0.0561598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_245_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_246_n 0.00510842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_247_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_303_n 0.0196855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_487_297#_c_352_n 0.00759381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_487_297#_c_353_n 0.0292274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_487_297#_c_354_n 0.00427601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_C1_c_65_n N_B1_c_105_n 0.0114603f $X=0.925 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_65 N_C1_M1009_g N_B1_M1005_g 0.0270285f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_66 N_C1_c_67_n B1 0.00248457f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_67 N_C1_c_67_n N_B1_c_108_n 0.0225797f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_68 N_C1_c_66_n N_VPWR_M1002_s 0.00779124f $X=0.24 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_69 N_C1_c_66_n N_VPWR_c_235_n 4.72765e-19 $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_70 N_C1_M1002_g N_VPWR_c_236_n 0.00316673f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_71 N_C1_c_66_n N_VPWR_c_236_n 0.0183612f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C1_M1002_g N_VPWR_c_237_n 6.68859e-19 $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_73 N_C1_M1009_g N_VPWR_c_237_n 0.0100534f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_74 N_C1_M1002_g N_VPWR_c_240_n 0.0054895f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_75 N_C1_M1009_g N_VPWR_c_240_n 0.00486043f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_76 N_C1_M1002_g N_VPWR_c_234_n 0.0106777f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_77 N_C1_M1009_g N_VPWR_c_234_n 0.00822531f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_78 N_C1_c_66_n N_VPWR_c_234_n 0.00201903f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C1_M1002_g N_Y_c_304_n 0.0155389f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_80 N_C1_M1009_g N_Y_c_305_n 0.0141904f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_81 N_C1_M1002_g N_Y_c_306_n 0.00284148f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_82 N_C1_M1009_g N_Y_c_306_n 0.00260149f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_83 N_C1_c_64_n N_Y_c_308_n 0.0156771f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_84 N_C1_M1002_g N_Y_c_308_n 0.00483315f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_85 N_C1_c_65_n N_Y_c_308_n 0.00580572f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_86 N_C1_M1009_g N_Y_c_308_n 0.00614436f $X=0.925 $Y=1.985 $X2=0 $Y2=0
cc_87 N_C1_c_66_n N_Y_c_308_n 0.0390015f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C1_c_67_n N_Y_c_308_n 0.0225172f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_89 N_C1_c_64_n N_A_27_47#_c_378_n 0.0121488f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_c_65_n N_A_27_47#_c_378_n 0.0121488f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_91 N_C1_c_66_n N_A_27_47#_c_378_n 0.00871283f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_92 N_C1_c_67_n N_A_27_47#_c_378_n 0.00175409f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_93 N_C1_c_64_n N_VGND_c_439_n 0.00357877f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_94 N_C1_c_65_n N_VGND_c_439_n 0.00357877f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_95 N_C1_c_64_n N_VGND_c_444_n 0.00622994f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_96 N_C1_c_65_n N_VGND_c_444_n 0.00530427f $X=0.925 $Y=0.995 $X2=0 $Y2=0
cc_97 B1 N_A2_c_154_n 0.0130184f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_98 N_B1_c_108_n N_A2_c_154_n 0.00174873f $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B1_M1005_g N_VPWR_c_237_n 0.00989496f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_100 N_B1_M1014_g N_VPWR_c_237_n 6.00419e-19 $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_101 N_B1_M1005_g N_VPWR_c_238_n 6.00419e-19 $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_102 N_B1_M1014_g N_VPWR_c_238_n 0.0109942f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_103 N_B1_M1005_g N_VPWR_c_241_n 0.00486043f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_104 N_B1_M1014_g N_VPWR_c_241_n 0.00486043f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_105 N_B1_M1005_g N_VPWR_c_234_n 0.00822531f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_106 N_B1_M1014_g N_VPWR_c_234_n 0.00822531f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_107 N_B1_M1005_g N_Y_c_305_n 0.0136034f $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_108 B1 N_Y_c_305_n 0.0274584f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B1_c_108_n N_Y_c_305_n 3.22594e-19 $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B1_M1014_g N_Y_c_303_n 0.0156905f $X=1.785 $Y=1.985 $X2=0 $Y2=0
cc_111 B1 N_Y_c_303_n 0.013958f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_112 B1 N_Y_c_319_n 0.0149215f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_113 N_B1_c_108_n N_Y_c_319_n 7.10237e-19 $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_105_n N_Y_c_308_n 5.69371e-19 $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B1_M1005_g N_Y_c_308_n 8.83454e-19 $X=1.355 $Y=1.985 $X2=0 $Y2=0
cc_116 B1 N_Y_c_308_n 0.0242465f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_117 N_B1_c_108_n N_Y_c_308_n 6.5392e-19 $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_118 B1 N_A_27_47#_c_379_n 0.015337f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_119 N_B1_c_108_n N_A_27_47#_c_379_n 6.09178e-19 $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_c_105_n N_A_27_47#_c_380_n 0.0104786f $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_106_n N_A_27_47#_c_380_n 0.00873911f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_122 B1 N_A_27_47#_c_380_n 0.00367704f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B1_c_105_n N_A_286_47#_c_406_n 0.0028282f $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B1_c_106_n N_A_286_47#_c_406_n 0.01238f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_125 B1 N_A_286_47#_c_406_n 0.0243676f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B1_c_108_n N_A_286_47#_c_406_n 0.00238284f $X=1.785 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B1_c_106_n N_VGND_c_435_n 0.00219146f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_c_105_n N_VGND_c_439_n 0.00357877f $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_c_106_n N_VGND_c_439_n 0.00357877f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_105_n N_VGND_c_444_n 0.00530427f $X=1.355 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_106_n N_VGND_c_444_n 0.00657863f $X=1.785 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A2_c_153_n N_A1_c_195_n 0.0265841f $X=3.205 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A2_M1007_g N_A1_M1011_g 0.0235424f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_134 N_A2_c_154_n N_A1_M1011_g 7.45547e-19 $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A2_c_154_n N_A1_c_197_n 0.00178044f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A2_c_155_n N_A1_c_197_n 0.0206299f $X=3.205 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A2_c_154_n A1 0.019437f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A2_c_155_n A1 6.58457e-19 $X=3.205 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A2_M1000_g N_VPWR_c_238_n 0.00546767f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A2_M1007_g N_VPWR_c_239_n 0.00107483f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_141 N_A2_M1000_g N_VPWR_c_242_n 0.00357877f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A2_M1007_g N_VPWR_c_242_n 0.00357877f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_143 N_A2_M1000_g N_VPWR_c_234_n 0.00657863f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_144 N_A2_M1007_g N_VPWR_c_234_n 0.00530427f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A2_M1000_g N_Y_c_303_n 0.0111217f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A2_c_154_n N_Y_c_303_n 0.0305971f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A2_M1000_g N_Y_c_327_n 0.0142626f $X=2.775 $Y=1.985 $X2=0 $Y2=0
cc_148 N_A2_M1007_g N_Y_c_327_n 0.00657002f $X=3.205 $Y=1.985 $X2=0 $Y2=0
cc_149 N_A2_c_154_n N_Y_c_327_n 0.0211595f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_155_n N_Y_c_327_n 7.11446e-19 $X=3.205 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_M1000_g N_A_487_297#_c_355_n 0.00926773f $X=2.775 $Y=1.985 $X2=0
+ $Y2=0
cc_152 N_A2_M1007_g N_A_487_297#_c_355_n 0.0114566f $X=3.205 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A2_c_152_n N_A_286_47#_c_406_n 0.0135285f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A2_c_153_n N_A_286_47#_c_406_n 0.0109444f $X=3.205 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_154_n N_A_286_47#_c_406_n 0.0509494f $X=3.17 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A2_c_155_n N_A_286_47#_c_406_n 0.00238284f $X=3.205 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_152_n N_VGND_c_435_n 0.00873326f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A2_c_153_n N_VGND_c_435_n 0.00104385f $X=3.205 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_152_n N_VGND_c_436_n 0.00104385f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_153_n N_VGND_c_436_n 0.00763402f $X=3.205 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_152_n N_VGND_c_440_n 0.00353537f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_153_n N_VGND_c_440_n 0.00353537f $X=3.205 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_152_n N_VGND_c_444_n 0.00415708f $X=2.775 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_153_n N_VGND_c_444_n 0.00415708f $X=3.205 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_M1011_g N_VPWR_c_239_n 0.0115361f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_166 N_A1_M1015_g N_VPWR_c_239_n 0.0122606f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A1_M1011_g N_VPWR_c_242_n 0.00486043f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_168 N_A1_M1015_g N_VPWR_c_243_n 0.00486043f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_169 N_A1_M1011_g N_VPWR_c_234_n 0.00825064f $X=3.635 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A1_M1015_g N_VPWR_c_234_n 0.00920993f $X=4.065 $Y=1.985 $X2=0 $Y2=0
cc_171 N_A1_M1011_g N_A_487_297#_c_352_n 0.0135976f $X=3.635 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A1_M1015_g N_A_487_297#_c_352_n 0.0160316f $X=4.065 $Y=1.985 $X2=0
+ $Y2=0
cc_173 N_A1_c_197_n N_A_487_297#_c_352_n 0.00222995f $X=4.065 $Y=1.16 $X2=0
+ $Y2=0
cc_174 A1 N_A_487_297#_c_352_n 0.0491777f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_175 N_A1_c_195_n N_A_286_47#_c_406_n 0.0109387f $X=3.635 $Y=0.995 $X2=0 $Y2=0
cc_176 A1 N_A_286_47#_c_406_n 0.0111255f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_177 N_A1_c_197_n N_A_286_47#_c_417_n 0.00241809f $X=4.065 $Y=1.16 $X2=0 $Y2=0
cc_178 A1 N_A_286_47#_c_417_n 0.0106143f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_179 A1 N_VGND_M1012_s 0.0039464f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_180 N_A1_c_195_n N_VGND_c_436_n 0.00763402f $X=3.635 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_196_n N_VGND_c_436_n 0.00104385f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_195_n N_VGND_c_438_n 0.00104385f $X=3.635 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_196_n N_VGND_c_438_n 0.00884918f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_184 A1 N_VGND_c_438_n 0.0129587f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_185 N_A1_c_195_n N_VGND_c_441_n 0.00353537f $X=3.635 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A1_c_196_n N_VGND_c_441_n 0.00486043f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_195_n N_VGND_c_444_n 0.00415708f $X=3.635 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_196_n N_VGND_c_444_n 0.00830219f $X=4.065 $Y=0.995 $X2=0 $Y2=0
cc_189 A1 N_VGND_c_444_n 0.00210615f $X=4.37 $Y=0.85 $X2=0 $Y2=0
cc_190 N_VPWR_c_234_n N_Y_M1002_d 0.00379452f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_234_n N_Y_M1005_d 0.00535672f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_234_n N_Y_M1000_s 0.00224864f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_240_n N_Y_c_304_n 0.0156896f $X=0.975 $Y=2.72 $X2=0 $Y2=0
cc_194 N_VPWR_c_234_n N_Y_c_304_n 0.00975383f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_M1009_s N_Y_c_305_n 0.00367486f $X=1 $Y=1.485 $X2=0 $Y2=0
cc_196 N_VPWR_c_237_n N_Y_c_305_n 0.0148206f $X=1.14 $Y=2 $X2=0 $Y2=0
cc_197 N_VPWR_c_241_n N_Y_c_338_n 0.0124538f $X=1.835 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_234_n N_Y_c_338_n 0.00724021f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_M1014_s N_Y_c_303_n 0.0111237f $X=1.86 $Y=1.485 $X2=0 $Y2=0
cc_200 N_VPWR_c_238_n N_Y_c_303_n 0.0191431f $X=2 $Y=2 $X2=0 $Y2=0
cc_201 N_VPWR_c_238_n N_Y_c_327_n 0.00521952f $X=2 $Y=2 $X2=0 $Y2=0
cc_202 N_VPWR_c_234_n N_A_487_297#_M1000_d 0.00212619f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_203 N_VPWR_c_234_n N_A_487_297#_M1007_d 0.00375984f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_234_n N_A_487_297#_M1015_s 0.00369639f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_242_n N_A_487_297#_c_355_n 0.0486451f $X=3.685 $Y=2.72 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_234_n N_A_487_297#_c_355_n 0.0307636f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VPWR_M1011_d N_A_487_297#_c_352_n 0.00351725f $X=3.71 $Y=1.485 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_239_n N_A_487_297#_c_352_n 0.0170777f $X=3.85 $Y=1.95 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_243_n N_A_487_297#_c_353_n 0.0178131f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_234_n N_A_487_297#_c_353_n 0.00993603f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_238_n N_A_487_297#_c_354_n 0.0241716f $X=2 $Y=2 $X2=0 $Y2=0
cc_212 N_VPWR_c_242_n N_A_487_297#_c_354_n 0.0170482f $X=3.685 $Y=2.72 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_234_n N_A_487_297#_c_354_n 0.00978235f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_Y_c_303_n N_A_487_297#_M1000_d 0.0063757f $X=2.825 $Y=1.625 $X2=-0.19
+ $Y2=1.305
cc_215 N_Y_M1000_s N_A_487_297#_c_355_n 0.0033237f $X=2.85 $Y=1.485 $X2=0 $Y2=0
cc_216 N_Y_c_303_n N_A_487_297#_c_355_n 0.0030313f $X=2.825 $Y=1.625 $X2=0 $Y2=0
cc_217 N_Y_c_327_n N_A_487_297#_c_355_n 0.0158133f $X=2.99 $Y=1.7 $X2=0 $Y2=0
cc_218 N_Y_c_303_n N_A_487_297#_c_354_n 0.0104783f $X=2.825 $Y=1.625 $X2=0 $Y2=0
cc_219 N_Y_M1004_s N_A_27_47#_c_378_n 0.00344076f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_220 N_Y_c_308_n N_A_27_47#_c_378_n 0.0126991f $X=0.71 $Y=0.76 $X2=0 $Y2=0
cc_221 N_Y_c_308_n N_A_27_47#_c_379_n 0.00840798f $X=0.71 $Y=0.76 $X2=0 $Y2=0
cc_222 N_Y_M1004_s N_VGND_c_444_n 0.00224864f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_380_n N_A_286_47#_M1001_s 0.00323923f $X=2 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_27_47#_M1013_d N_A_286_47#_c_406_n 0.0124861f $X=1.86 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_380_n N_A_286_47#_c_406_n 0.0410385f $X=2 $Y=0.36 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_380_n N_VGND_c_435_n 0.0135209f $X=2 $Y=0.36 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_378_n N_VGND_c_439_n 0.0539155f $X=1.045 $Y=0.35 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_380_n N_VGND_c_439_n 0.0529196f $X=2 $Y=0.36 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_399_p N_VGND_c_439_n 0.0124663f $X=1.14 $Y=0.36 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1004_d N_VGND_c_444_n 0.00229841f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_M1006_d N_VGND_c_444_n 0.00223239f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_232 N_A_27_47#_M1013_d N_VGND_c_444_n 0.00229841f $X=1.86 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_378_n N_VGND_c_444_n 0.0339576f $X=1.045 $Y=0.35 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_380_n N_VGND_c_444_n 0.033285f $X=2 $Y=0.36 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_399_p N_VGND_c_444_n 0.00730424f $X=1.14 $Y=0.36 $X2=0 $Y2=0
cc_236 N_A_286_47#_c_406_n N_VGND_M1003_d 0.00645735f $X=3.755 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_237 N_A_286_47#_c_406_n N_VGND_M1010_d 0.00828556f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_286_47#_c_406_n N_VGND_c_435_n 0.0188779f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_239 N_A_286_47#_c_406_n N_VGND_c_436_n 0.0146754f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_286_47#_c_406_n N_VGND_c_439_n 0.00425741f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_286_47#_c_406_n N_VGND_c_440_n 0.00817434f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_286_47#_c_406_n N_VGND_c_441_n 0.00249635f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_286_47#_c_417_n N_VGND_c_441_n 0.00435302f $X=3.85 $Y=0.68 $X2=0
+ $Y2=0
cc_244 N_A_286_47#_M1001_s N_VGND_c_444_n 0.00224864f $X=1.43 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_286_47#_M1003_s N_VGND_c_444_n 0.00326987f $X=2.85 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_286_47#_M1008_d N_VGND_c_444_n 0.00437709f $X=3.71 $Y=0.235 $X2=0
+ $Y2=0
cc_247 N_A_286_47#_c_406_n N_VGND_c_444_n 0.0293518f $X=3.755 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_286_47#_c_417_n N_VGND_c_444_n 0.00598996f $X=3.85 $Y=0.68 $X2=0
+ $Y2=0

* File: sky130_fd_sc_hd__dlrbn_1.pex.spice
* Created: Thu Aug 27 14:16:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DLRBN_1%GATE_N 4 5 7 8 10 13 17 19 20 24 26
c43 19 0 5.39299e-20 $X=0.23 $Y=1.19
c44 13 0 2.71124e-20 $X=0.47 $Y=0.805
r45 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r46 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r47 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r48 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r49 15 17 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=1.665
+ $X2=0.47 $Y2=1.665
r50 11 13 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.47 $Y2=0.805
r51 8 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=1.74 $X2=0.47
+ $Y2=1.665
r52 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.47 $Y=1.74
+ $X2=0.47 $Y2=2.135
r53 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.805
r54 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r55 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r56 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r57 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r58 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_27_47# 1 2 9 13 17 20 24 28 29 30 38 42 45
+ 47 52 54 56 57 60 63 64 68 71 75 79
c168 20 0 1.41946e-19 $X=3.335 $Y=2.275
c169 13 0 2.6965e-20 $X=0.89 $Y=2.135
c170 9 0 2.6965e-20 $X=0.89 $Y=0.445
r171 64 79 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=3.095 $Y2=1.415
r172 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.015 $Y=1.53
+ $X2=3.015 $Y2=1.53
r173 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.695 $Y=1.53
+ $X2=0.695 $Y2=1.53
r174 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.84 $Y=1.53
+ $X2=0.695 $Y2=1.53
r175 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=3.015 $Y2=1.53
r176 56 57 2.51237 $w=1.4e-07 $l=2.03e-06 $layer=MET1_cond $X=2.87 $Y=1.53
+ $X2=0.84 $Y2=1.53
r177 52 71 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=0.87
+ $X2=2.8 $Y2=0.705
r178 51 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.8 $Y=0.87
+ $X2=3.01 $Y2=0.87
r179 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.8
+ $Y=0.87 $X2=2.8 $Y2=0.87
r180 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=1.795
+ $X2=0.695 $Y2=1.53
r181 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.695 $Y=1.4
+ $X2=0.695 $Y2=1.53
r182 46 68 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=0.755 $Y=1.235
+ $X2=0.89 $Y2=1.235
r183 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.4
r184 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.235
+ $X2=0.725 $Y2=1.07
r185 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.235 $X2=0.755 $Y2=1.235
r186 39 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=3.18 $Y=1.74
+ $X2=3.335 $Y2=1.74
r187 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.74 $X2=3.18 $Y2=1.74
r188 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.53
r189 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=1.585
+ $X2=3.095 $Y2=1.74
r190 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=0.87
r191 34 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.01 $Y=1.035
+ $X2=3.01 $Y2=1.415
r192 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.695 $Y=0.805
+ $X2=0.695 $Y2=1.07
r193 31 42 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.215 $Y2=1.88
r194 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.695 $Y2=1.795
r195 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=1.88
+ $X2=0.345 $Y2=1.88
r196 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.695 $Y2=0.805
r197 28 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.345 $Y2=0.72
r198 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.345 $Y2=0.72
r199 22 24 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.215 $Y=0.635
+ $X2=0.215 $Y2=0.51
r200 18 75 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=1.74
r201 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.335 $Y=1.875
+ $X2=3.335 $Y2=2.275
r202 17 71 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.415
+ $X2=2.79 $Y2=0.705
r203 11 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=1.235
r204 11 13 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.89 $Y=1.37
+ $X2=0.89 $Y2=2.135
r205 7 68 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.89 $Y=1.1
+ $X2=0.89 $Y2=1.235
r206 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.89 $Y=1.1 $X2=0.89
+ $Y2=0.445
r207 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r208 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%D 3 7 9 13 15
c40 13 0 1.12109e-19 $X=1.625 $Y=1.04
r41 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.625 $Y=1.04
+ $X2=1.83 $Y2=1.04
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.04 $X2=1.625 $Y2=1.04
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.625 $Y=1.19
+ $X2=1.625 $Y2=1.04
r44 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.205
+ $X2=1.83 $Y2=1.04
r45 5 7 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.83 $Y=1.205 $X2=1.83
+ $Y2=2.165
r46 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=0.875
+ $X2=1.83 $Y2=1.04
r47 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.83 $Y=0.875 $X2=1.83
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_299_47# 1 2 9 12 16 18 20 21 22 23 25 32
+ 34
c83 32 0 1.12109e-19 $X=2.255 $Y=0.93
c84 18 0 7.13094e-20 $X=1.97 $Y=0.7
r85 32 35 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=1.095
r86 32 34 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.93
+ $X2=2.255 $Y2=0.765
r87 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r88 25 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.51
+ $X2=1.62 $Y2=0.7
r89 22 31 8.96794 $w=3.07e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.155 $Y2=0.93
r90 22 23 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.055 $Y=1.095
+ $X2=2.055 $Y2=1.495
r91 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=2.055 $Y2=1.495
r92 20 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.97 $Y=1.58
+ $X2=1.785 $Y2=1.58
r93 19 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.7
+ $X2=1.62 $Y2=0.7
r94 18 31 9.14007 $w=3.07e-07 $l=3.0895e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=2.155 $Y2=0.93
r95 18 19 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.97 $Y=0.7
+ $X2=1.705 $Y2=0.7
r96 14 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.785 $Y2=1.58
r97 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.99
r98 12 35 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.25 $Y=2.165
+ $X2=2.25 $Y2=1.095
r99 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.765
r100 2 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.845 $X2=1.62 $Y2=1.99
r101 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_193_47# 1 2 9 11 12 15 19 22 24 26 27 30
+ 33 37 38
c112 38 0 1.41946e-19 $X=2.67 $Y=1.52
r113 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.52 $X2=2.67 $Y2=1.52
r114 34 38 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.612 $Y=1.87
+ $X2=2.612 $Y2=1.52
r115 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=1.87
+ $X2=2.555 $Y2=1.87
r116 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.155 $Y=1.87
+ $X2=1.155 $Y2=1.87
r117 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.3 $Y=1.87
+ $X2=1.155 $Y2=1.87
r118 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=2.555 $Y2=1.87
r119 26 27 1.37376 $w=1.4e-07 $l=1.11e-06 $layer=MET1_cond $X=2.41 $Y=1.87
+ $X2=1.3 $Y2=1.87
r120 24 30 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.87
r121 24 25 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.127 $Y=1.797
+ $X2=1.127 $Y2=1.685
r122 22 25 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.1 $Y=0.51
+ $X2=1.1 $Y2=1.685
r123 18 37 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=2.67 $Y=1.55 $X2=2.67
+ $Y2=1.52
r124 18 19 41.7507 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=2.67 $Y=1.55
+ $X2=2.67 $Y2=1.685
r125 17 37 27.7717 $w=2.7e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.395
+ $X2=2.67 $Y2=1.52
r126 13 15 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.22 $Y=1.245
+ $X2=3.22 $Y2=0.415
r127 12 17 79.8255 $w=7.8e-08 $l=1.68375e-07 $layer=POLY_cond $X=2.805 $Y=1.32
+ $X2=2.67 $Y2=1.395
r128 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=3.22 $Y2=1.245
r129 11 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.145 $Y=1.32
+ $X2=2.805 $Y2=1.32
r130 9 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.73 $Y=2.275
+ $X2=2.73 $Y2=1.685
r131 2 30 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.965
+ $Y=1.815 $X2=1.1 $Y2=1.96
r132 1 22 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_724_21# 1 2 9 13 15 17 20 22 23 24 25 26
+ 28 29 31 35 37 40 42 45 46 49 51 56 59
c128 9 0 1.07053e-19 $X=3.695 $Y=0.445
r129 57 66 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.79 $Y=1.16
+ $X2=5.935 $Y2=1.16
r130 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.79
+ $Y=1.16 $X2=5.79 $Y2=1.16
r131 54 56 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=5.75 $Y=1.535
+ $X2=5.75 $Y2=1.16
r132 53 56 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.75 $Y=0.825
+ $X2=5.75 $Y2=1.16
r133 52 59 4.04103 $w=2.8e-07 $l=1.27574e-07 $layer=LI1_cond $X=4.97 $Y=1.65
+ $X2=4.865 $Y2=1.7
r134 51 54 6.8319 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=5.625 $Y=1.65
+ $X2=5.75 $Y2=1.535
r135 51 52 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.625 $Y=1.65
+ $X2=4.97 $Y2=1.65
r136 47 59 2.39622 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=1.865
+ $X2=4.865 $Y2=1.7
r137 47 49 21.3896 $w=2.08e-07 $l=4.05e-07 $layer=LI1_cond $X=4.865 $Y=1.865
+ $X2=4.865 $Y2=2.27
r138 45 53 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.625 $Y=0.74
+ $X2=5.75 $Y2=0.825
r139 45 46 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=5.625 $Y=0.74
+ $X2=4.54 $Y2=0.74
r140 42 46 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.39 $Y=0.655
+ $X2=4.54 $Y2=0.74
r141 42 44 3.86333 $w=3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.39 $Y=0.655 $X2=4.39
+ $Y2=0.56
r142 40 60 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.925 $Y=1.7
+ $X2=3.695 $Y2=1.7
r143 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.925
+ $Y=1.7 $X2=3.925 $Y2=1.7
r144 37 59 4.04103 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=4.76 $Y=1.7
+ $X2=4.865 $Y2=1.7
r145 37 39 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=4.76 $Y=1.7
+ $X2=3.925 $Y2=1.7
r146 33 35 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=6.745 $Y=1.695
+ $X2=6.875 $Y2=1.695
r147 29 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.875 $Y=1.77
+ $X2=6.875 $Y2=1.695
r148 29 31 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.875 $Y=1.77
+ $X2=6.875 $Y2=2.165
r149 26 28 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.875 $Y=0.73
+ $X2=6.875 $Y2=0.445
r150 25 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.745 $Y=1.62
+ $X2=6.745 $Y2=1.695
r151 24 25 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=6.745 $Y=1.325
+ $X2=6.745 $Y2=1.62
r152 23 66 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=1.16
+ $X2=5.935 $Y2=1.16
r153 22 24 45.3305 $w=1.82e-07 $l=1.94808e-07 $layer=POLY_cond $X=6.81 $Y=1.16
+ $X2=6.745 $Y2=1.325
r154 22 26 115.512 $w=1.82e-07 $l=4.61357e-07 $layer=POLY_cond $X=6.81 $Y=1.16
+ $X2=6.875 $Y2=0.73
r155 22 23 115.408 $w=3.3e-07 $l=6.6e-07 $layer=POLY_cond $X=6.67 $Y=1.16
+ $X2=6.01 $Y2=1.16
r156 18 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=1.325
+ $X2=5.935 $Y2=1.16
r157 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.935 $Y=1.325
+ $X2=5.935 $Y2=1.985
r158 15 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=0.995
+ $X2=5.935 $Y2=1.16
r159 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.935 $Y=0.995
+ $X2=5.935 $Y2=0.56
r160 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=1.7
r161 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.695 $Y=1.865
+ $X2=3.695 $Y2=2.275
r162 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=1.7
r163 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.695 $Y=1.535
+ $X2=3.695 $Y2=0.445
r164 2 59 600 $w=1.7e-07 $l=3.46627e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.885 $Y2=1.755
r165 2 49 600 $w=1.7e-07 $l=8.68101e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.485 $X2=4.885 $Y2=2.27
r166 1 44 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.235 $X2=4.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_561_413# 1 2 7 9 12 14 15 16 20 25 26 27
+ 30
c82 30 0 1.20256e-19 $X=4.135 $Y=1.16
c83 26 0 1.65126e-19 $X=3.565 $Y=1.325
r84 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.135
+ $Y=1.16 $X2=4.135 $Y2=1.16
r85 28 30 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.65 $Y=1.16
+ $X2=4.135 $Y2=1.16
r86 26 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.49 $Y2=1.16
r87 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.565 $Y=1.325
+ $X2=3.565 $Y2=2.255
r88 25 28 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.415 $Y=0.995
+ $X2=3.49 $Y2=1.16
r89 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.415 $Y=0.535
+ $X2=3.415 $Y2=0.995
r90 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.565 $Y2=2.255
r91 20 22 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.48 $Y=2.34
+ $X2=3.065 $Y2=2.34
r92 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.415 $Y2=0.535
r93 16 18 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.45
+ $X2=3.005 $Y2=0.45
r94 14 31 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.135 $Y2=1.16
r95 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.635 $Y2=1.16
r96 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.16
r97 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.635 $Y=1.325
+ $X2=4.635 $Y2=1.985
r98 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.635 $Y=0.995
+ $X2=4.635 $Y2=0.56
r100 2 22 600 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.065 $X2=3.065 $Y2=2.34
r101 1 18 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.235 $X2=3.005 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%RESET_B 3 6 8 9 13 15 22
c36 13 0 1.20256e-19 $X=5.055 $Y=1.16
c37 9 0 1.07053e-19 $X=5.25 $Y=1.105
r38 14 22 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.055 $Y=1.16
+ $X2=5.295 $Y2=1.16
r39 13 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.16
+ $X2=5.055 $Y2=1.325
r40 13 15 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.16
+ $X2=5.055 $Y2=0.995
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.16 $X2=5.055 $Y2=1.16
r42 9 22 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=5.335 $Y=1.16 $X2=5.295
+ $Y2=1.16
r43 8 14 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.875 $Y=1.16
+ $X2=5.055 $Y2=1.16
r44 6 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.095 $Y=1.985
+ $X2=5.095 $Y2=1.325
r45 3 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.095 $Y=0.56
+ $X2=5.095 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%A_1308_47# 1 2 9 12 16 20 24 25 27 29
r47 25 30 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.285 $Y=1.16
+ $X2=7.285 $Y2=1.325
r48 25 29 46.1296 $w=3.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.285 $Y=1.16
+ $X2=7.285 $Y2=0.995
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.305
+ $Y=1.16 $X2=7.305 $Y2=1.16
r50 22 27 0.221902 $w=3.3e-07 $l=1.27475e-07 $layer=LI1_cond $X=6.83 $Y=1.16
+ $X2=6.705 $Y2=1.155
r51 22 24 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=6.83 $Y=1.16
+ $X2=7.305 $Y2=1.16
r52 18 27 7.38875 $w=2.1e-07 $l=1.7e-07 $layer=LI1_cond $X=6.705 $Y=1.325
+ $X2=6.705 $Y2=1.155
r53 18 20 38.7221 $w=2.48e-07 $l=8.4e-07 $layer=LI1_cond $X=6.705 $Y=1.325
+ $X2=6.705 $Y2=2.165
r54 14 27 7.38875 $w=2.1e-07 $l=1.88944e-07 $layer=LI1_cond $X=6.665 $Y=0.985
+ $X2=6.705 $Y2=1.155
r55 14 16 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.665 $Y=0.985
+ $X2=6.665 $Y2=0.51
r56 12 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.35 $Y=1.985
+ $X2=7.35 $Y2=1.325
r57 9 29 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.35 $Y=0.56 $X2=7.35
+ $Y2=0.995
r58 2 20 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.845 $X2=6.665 $Y2=2.165
r59 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.54
+ $Y=0.235 $X2=6.665 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 46 51
+ 59 60 64 71 72 75 78 85 92
r113 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r114 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 85 88 11.3143 $w=7.38e-07 $l=7e-07 $layer=LI1_cond $X=5.52 $Y=2.02 $X2=5.52
+ $Y2=2.72
r116 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r117 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r118 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 72 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r120 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r121 69 92 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.305 $Y=2.72
+ $X2=7.157 $Y2=2.72
r122 69 71 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.305 $Y=2.72
+ $X2=7.59 $Y2=2.72
r123 68 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r124 68 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r125 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r126 65 88 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=2.72
+ $X2=5.52 $Y2=2.72
r127 65 67 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.89 $Y=2.72
+ $X2=6.67 $Y2=2.72
r128 64 92 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=7.157 $Y2=2.72
r129 64 67 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.01 $Y=2.72
+ $X2=6.67 $Y2=2.72
r130 63 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r131 63 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r133 60 82 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.59 $Y=2.72
+ $X2=4.37 $Y2=2.72
r134 60 62 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.59 $Y=2.72
+ $X2=4.83 $Y2=2.72
r135 59 88 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=2.72
+ $X2=5.52 $Y2=2.72
r136 59 62 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.15 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 58 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r140 55 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 54 57 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r142 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r143 52 78 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.112 $Y2=2.72
r144 52 54 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r145 51 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.82 $Y=2.72
+ $X2=3.45 $Y2=2.72
r146 50 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 50 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r149 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=0.68 $Y2=2.72
r150 47 49 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 46 78 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=2.112 $Y2=2.72
r152 46 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.61 $Y2=2.72
r153 41 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.68 $Y2=2.72
r154 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r155 39 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r156 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r157 35 92 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.157 $Y=2.635
+ $X2=7.157 $Y2=2.72
r158 35 37 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=7.157 $Y=2.635
+ $X2=7.157 $Y2=2
r159 33 82 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.425 $Y=2.34
+ $X2=4.425 $Y2=2.635
r160 27 82 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=4.37 $Y2=2.72
r161 27 51 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=2.72
+ $X2=3.82 $Y2=2.72
r162 27 29 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.955 $Y=2.635
+ $X2=3.955 $Y2=2.3
r163 23 78 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2.72
r164 23 25 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.112 $Y=2.635
+ $X2=2.112 $Y2=2
r165 19 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.72
r166 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.68 $Y=2.635
+ $X2=0.68 $Y2=2.22
r167 6 37 300 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_PDIFF $count=2 $X=6.95
+ $Y=1.845 $X2=7.14 $Y2=2
r168 5 85 150 $w=1.7e-07 $l=7.77785e-07 $layer=licon1_PDIFF $count=4 $X=5.17
+ $Y=1.485 $X2=5.725 $Y2=2.02
r169 4 33 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.485 $X2=4.425 $Y2=2.34
r170 3 29 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=2.065 $X2=3.905 $Y2=2.3
r171 2 25 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.845 $X2=2.04 $Y2=2
r172 1 21 600 $w=1.7e-07 $l=4.67654e-07 $layer=licon1_PDIFF $count=1 $X=0.545
+ $Y=1.815 $X2=0.68 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%Q 1 2 7 8 9 10 11 12
r18 12 32 9.00346 $w=3.18e-07 $l=2.5e-07 $layer=LI1_cond $X=6.22 $Y=2.21
+ $X2=6.22 $Y2=1.96
r19 11 32 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=6.22 $Y=1.87 $X2=6.22
+ $Y2=1.96
r20 10 11 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=6.22 $Y=1.53
+ $X2=6.22 $Y2=1.87
r21 9 10 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=6.22 $Y=1.19 $X2=6.22
+ $Y2=1.53
r22 8 9 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=6.22 $Y=0.85 $X2=6.22
+ $Y2=1.19
r23 7 8 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=6.22 $Y=0.51 $X2=6.22
+ $Y2=0.85
r24 2 32 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=6.01
+ $Y=1.485 $X2=6.145 $Y2=1.96
r25 1 7 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=6.01
+ $Y=0.235 $X2=6.145 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%Q_N 1 2 7 8 9 34
r13 16 34 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=7.605 $Y=1.915
+ $X2=7.605 $Y2=1.87
r14 8 34 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=7.605 $Y=1.85
+ $X2=7.605 $Y2=1.87
r15 8 9 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=7.605 $Y=1.935
+ $X2=7.605 $Y2=2.21
r16 8 16 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=7.605 $Y=1.935
+ $X2=7.605 $Y2=1.915
r17 7 8 46.3094 $w=1.73e-07 $l=1.19e-06 $layer=LI1_cond $X=7.647 $Y=0.595
+ $X2=7.647 $Y2=1.785
r18 2 8 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=7.425
+ $Y=1.485 $X2=7.56 $Y2=1.96
r19 1 7 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.235 $X2=7.56 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HD__DLRBN_1%VGND 1 2 3 4 5 18 22 26 30 32 34 39 44 57 64
+ 65 68 71 74 79 85 87
c115 65 0 2.71124e-20 $X=7.59 $Y=0
c116 2 0 7.13094e-20 $X=1.905 $Y=0.235
r117 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r118 83 85 9.12166 $w=5.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.75 $Y=0.2
+ $X2=5.875 $Y2=0.2
r119 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r120 81 83 0.839353 $w=5.68e-07 $l=4e-08 $layer=LI1_cond $X=5.71 $Y=0.2 $X2=5.75
+ $Y2=0.2
r121 78 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r122 77 81 8.81321 $w=5.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.71 $Y2=0.2
r123 77 79 9.75117 $w=5.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.29 $Y=0.2
+ $X2=5.135 $Y2=0.2
r124 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r125 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r126 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r127 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r128 65 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=7.13
+ $Y2=0
r129 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r130 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.14
+ $Y2=0
r131 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.305 $Y=0
+ $X2=7.59 $Y2=0
r132 61 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r133 61 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=5.75
+ $Y2=0
r134 60 85 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=5.875 $Y2=0
r135 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r136 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=7.14
+ $Y2=0
r137 57 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=6.67 $Y2=0
r138 56 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r139 56 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r140 55 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=5.135 $Y2=0
r141 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r142 53 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.905
+ $Y2=0
r143 53 55 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.83
+ $Y2=0
r144 51 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r145 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r146 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r147 48 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r148 47 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r149 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r150 45 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.04
+ $Y2=0
r151 45 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0
+ $X2=2.53 $Y2=0
r152 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.905
+ $Y2=0
r153 44 50 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.45
+ $Y2=0
r154 43 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r155 43 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r156 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r157 40 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.68
+ $Y2=0
r158 40 42 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=1.61 $Y2=0
r159 39 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.04
+ $Y2=0
r160 39 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.61 $Y2=0
r161 34 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.68
+ $Y2=0
r162 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r163 32 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r164 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r165 28 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0
r166 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.14 $Y=0.085
+ $X2=7.14 $Y2=0.38
r167 24 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0
r168 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.905 $Y=0.085
+ $X2=3.905 $Y2=0.445
r169 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0
r170 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.04 $Y=0.085
+ $X2=2.04 $Y2=0.36
r171 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0
r172 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.68 $Y=0.085
+ $X2=0.68 $Y2=0.38
r173 5 30 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.235 $X2=7.14 $Y2=0.38
r174 4 81 91 $w=1.7e-07 $l=5.9925e-07 $layer=licon1_NDIFF $count=2 $X=5.17
+ $Y=0.235 $X2=5.71 $Y2=0.36
r175 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.77
+ $Y=0.235 $X2=3.905 $Y2=0.445
r176 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.04 $Y2=0.36
r177 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.38
.ends


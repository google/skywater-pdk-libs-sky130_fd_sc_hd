* File: sky130_fd_sc_hd__lpflow_clkbufkapwr_4.spice.SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4.pxi
* Created: Thu Aug 27 14:23:34 2020
* 
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A N_A_M1003_g N_A_M1006_g A A
+ N_A_c_51_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A_27_47# N_A_27_47#_M1003_s
+ N_A_27_47#_M1006_s N_A_27_47#_M1002_g N_A_27_47#_M1000_g N_A_27_47#_M1007_g
+ N_A_27_47#_M1001_g N_A_27_47#_M1008_g N_A_27_47#_M1004_g N_A_27_47#_M1009_g
+ N_A_27_47#_M1005_g N_A_27_47#_c_94_n N_A_27_47#_c_102_n N_A_27_47#_c_114_n
+ N_A_27_47#_c_103_n N_A_27_47#_c_119_n N_A_27_47#_c_147_p N_A_27_47#_c_95_n
+ N_A_27_47#_c_104_n N_A_27_47#_c_96_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%A_27_47#
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%KAPWR N_KAPWR_M1006_d N_KAPWR_M1007_s
+ N_KAPWR_M1009_s N_KAPWR_c_200_n N_KAPWR_c_201_n N_KAPWR_c_210_n
+ N_KAPWR_c_212_n N_KAPWR_c_215_n N_KAPWR_c_218_n KAPWR N_KAPWR_c_203_n
+ N_KAPWR_c_238_p KAPWR PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%X N_X_M1000_d N_X_M1004_d N_X_M1002_d
+ N_X_M1008_d N_X_c_256_n N_X_c_269_n N_X_c_257_n N_X_c_258_n N_X_c_279_n
+ N_X_c_283_n N_X_c_259_n N_X_c_313_n X X X N_X_c_262_n
+ PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%X
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VGND N_VGND_M1003_d N_VGND_M1001_s
+ N_VGND_M1005_s N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n
+ VGND N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VGND
x_PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VPWR VPWR N_VPWR_c_387_n
+ N_VPWR_c_386_n PM_SKY130_FD_SC_HD__LPFLOW_CLKBUFKAPWR_4%VPWR
cc_1 VNB N_A_M1003_g 0.0322943f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.445
cc_2 VNB A 0.00620969f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_3 VNB N_A_c_51_n 0.0251851f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_A_27_47#_M1002_g 4.17371e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_5 VNB N_A_27_47#_M1000_g 0.0295782f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_6 VNB N_A_27_47#_M1007_g 4.55724e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_7 VNB N_A_27_47#_M1001_g 0.0276999f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_8 VNB N_A_27_47#_M1008_g 4.56723e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1004_g 0.0276748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1009_g 5.58244e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1005_g 0.0366072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_94_n 0.0330143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_95_n 0.0131987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_96_n 0.0706034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_X_c_256_n 6.31183e-19 $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_16 VNB N_X_c_257_n 0.00518223f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_17 VNB N_X_c_258_n 0.00217909f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.19
cc_18 VNB N_X_c_259_n 0.00204615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB X 0.0337654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_341_n 0.00475331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_342_n 0.00404131f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_22 VNB N_VGND_c_343_n 0.0120207f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.85
cc_23 VNB N_VGND_c_344_n 0.00474766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_345_n 0.0164986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_346_n 0.0175222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_347_n 0.0158977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_348_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_349_n 0.0048778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_350_n 0.161822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_386_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.765
cc_31 VPB N_A_M1006_g 0.0229606f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.985
cc_32 VPB A 0.00221579f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_33 VPB N_A_c_51_n 0.00537042f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_34 VPB N_A_27_47#_M1002_g 0.0198993f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_35 VPB N_A_27_47#_M1007_g 0.0197727f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_36 VPB N_A_27_47#_M1008_g 0.0197632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_M1009_g 0.0240996f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_94_n 0.00904608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_102_n 0.0261567f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_103_n 0.00175845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_104_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_KAPWR_c_200_n 0.00994025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_KAPWR_c_201_n 0.00876329f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.85
cc_44 VPB X 0.0058073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_X_c_262_n 0.012335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_387_n 0.0747018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_386_n 0.0423834f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.765
cc_48 N_A_M1006_g N_A_27_47#_M1002_g 0.0228414f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_A_27_47#_M1000_g 0.0183348f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_50 A N_A_27_47#_M1000_g 0.0050309f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_51 N_A_c_51_n N_A_27_47#_M1000_g 0.00287228f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_A_27_47#_c_94_n 0.0101619f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_53 N_A_M1006_g N_A_27_47#_c_94_n 0.0059274f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_94_n 0.0429918f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_55 N_A_c_51_n N_A_27_47#_c_94_n 0.00797697f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_M1006_g N_A_27_47#_c_102_n 0.004518f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_57 N_A_M1006_g N_A_27_47#_c_114_n 0.0104162f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_58 A N_A_27_47#_c_114_n 0.0251553f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_59 N_A_c_51_n N_A_27_47#_c_114_n 5.45329e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_M1006_g N_A_27_47#_c_103_n 9.07197e-19 $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_61 A N_A_27_47#_c_103_n 0.00600199f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_62 A N_A_27_47#_c_119_n 0.0143279f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_63 A N_A_27_47#_c_96_n 0.00251756f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_c_51_n N_A_27_47#_c_96_n 0.0154138f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_KAPWR_c_201_n 0.00240782f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_66 N_A_M1006_g N_KAPWR_c_203_n 0.0064863f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_X_c_256_n 7.63641e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_X_c_258_n 2.1267e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_X_c_258_n 0.00990658f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_VGND_c_341_n 0.00318753f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_71 A N_VGND_c_341_n 0.0152693f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_72 N_A_c_51_n N_VGND_c_341_n 3.07485e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_M1003_g N_VGND_c_345_n 0.00466641f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 A N_VGND_c_345_n 0.00176987f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_VGND_c_350_n 0.00775648f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_76 A N_VGND_c_350_n 0.00378105f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_VPWR_c_387_n 0.0054895f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_78 N_A_M1006_g N_VPWR_c_386_n 0.00619867f $X=0.475 $Y=1.985 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_114_n N_KAPWR_M1006_d 0.00577523f $X=0.945 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_47#_M1008_g N_KAPWR_c_200_n 0.00211474f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_81 N_A_27_47#_M1009_g N_KAPWR_c_200_n 0.00341645f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_82 N_A_27_47#_M1006_s N_KAPWR_c_201_n 7.18041e-19 $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_83 N_A_27_47#_c_102_n N_KAPWR_c_201_n 0.0285517f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_114_n N_KAPWR_c_201_n 0.00509698f $X=0.945 $Y=1.58 $X2=0
+ $Y2=0
cc_85 N_A_27_47#_c_102_n N_KAPWR_c_210_n 4.3931e-19 $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_114_n N_KAPWR_c_210_n 0.00127334f $X=0.945 $Y=1.58 $X2=0
+ $Y2=0
cc_87 N_A_27_47#_M1002_g N_KAPWR_c_212_n 2.13337e-19 $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_88 N_A_27_47#_M1007_g N_KAPWR_c_212_n 0.00301408f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_89 N_A_27_47#_M1008_g N_KAPWR_c_212_n 0.00301408f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_M1002_g N_KAPWR_c_215_n 0.00279183f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_M1007_g N_KAPWR_c_215_n 0.00185592f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_c_114_n N_KAPWR_c_215_n 0.00568827f $X=0.945 $Y=1.58 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_M1007_g N_KAPWR_c_218_n 8.6046e-19 $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_M1008_g N_KAPWR_c_218_n 9.69549e-19 $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_102_n N_KAPWR_c_203_n 0.0262387f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_114_n N_KAPWR_c_203_n 0.0184355f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_114_n N_X_M1002_d 0.00266014f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1000_g N_X_c_256_n 0.00655439f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1001_g N_X_c_256_n 0.00115565f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_27_47#_M1002_g N_X_c_269_n 0.00437181f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_27_47#_M1007_g N_X_c_269_n 7.04672e-19 $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_27_47#_M1001_g N_X_c_257_n 0.0122792f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_27_47#_M1004_g N_X_c_257_n 0.0122792f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_147_p N_X_c_257_n 0.054594f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_96_n N_X_c_257_n 0.0023301f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_106 N_A_27_47#_M1000_g N_X_c_258_n 0.00456754f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_119_n N_X_c_258_n 0.00901782f $X=1.115 $Y=1.16 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_147_p N_X_c_258_n 0.0150434f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_96_n N_X_c_258_n 0.00240878f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_110 N_A_27_47#_M1007_g N_X_c_279_n 0.00696893f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_27_47#_M1008_g N_X_c_279_n 0.012546f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_147_p N_X_c_279_n 0.0131166f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_96_n N_X_c_279_n 0.00181808f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_114 N_A_27_47#_M1002_g N_X_c_283_n 0.00447897f $X=0.955 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_27_47#_M1007_g N_X_c_283_n 0.00830056f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_114_n N_X_c_283_n 0.00275116f $X=0.945 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_147_p N_X_c_283_n 0.007234f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_96_n N_X_c_283_n 0.00180683f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1004_g N_X_c_259_n 0.00114296f $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1005_g N_X_c_259_n 0.00216977f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1008_g X 6.2445e-19 $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1004_g X 6.0408e-19 $X=1.82 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_27_47#_M1009_g X 0.00525161f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_124 N_A_27_47#_M1005_g X 0.018959f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_27_47#_c_147_p X 0.0136122f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_96_n X 0.0174538f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1008_g N_X_c_262_n 0.00226561f $X=1.815 $Y=1.985 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1009_g N_X_c_262_n 0.012256f $X=2.245 $Y=1.985 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_147_p N_X_c_262_n 0.0128752f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_96_n N_X_c_262_n 0.00233619f $X=2.245 $Y=1.157 $X2=0 $Y2=0
cc_131 N_A_27_47#_M1000_g N_VGND_c_341_n 0.00157173f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_M1001_g N_VGND_c_342_n 0.00166998f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_M1004_g N_VGND_c_342_n 0.00159632f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_M1005_g N_VGND_c_344_n 0.00341661f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_95_n N_VGND_c_345_n 0.0186529f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_136 N_A_27_47#_M1000_g N_VGND_c_346_n 0.0055185f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1001_g N_VGND_c_346_n 0.00439206f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_M1004_g N_VGND_c_347_n 0.00439206f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_M1005_g N_VGND_c_347_n 0.00439206f $X=2.25 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1003_s N_VGND_c_350_n 0.00262044f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_M1000_g N_VGND_c_350_n 0.00995296f $X=0.96 $Y=0.445 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1001_g N_VGND_c_350_n 0.00590932f $X=1.39 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1004_g N_VGND_c_350_n 0.00592186f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1005_g N_VGND_c_350_n 0.0068734f $X=2.25 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_95_n N_VGND_c_350_n 0.0113402f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_146 N_A_27_47#_M1002_g N_VPWR_c_387_n 0.00579312f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_M1007_g N_VPWR_c_387_n 0.00426947f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_M1008_g N_VPWR_c_387_n 0.00428402f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_M1009_g N_VPWR_c_387_n 0.00585385f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_c_102_n N_VPWR_c_387_n 0.0185301f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_151 N_A_27_47#_M1006_s N_VPWR_c_386_n 0.00127304f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_M1002_g N_VPWR_c_386_n 0.00535792f $X=0.955 $Y=1.985 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_M1007_g N_VPWR_c_386_n 0.00491693f $X=1.385 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_M1008_g N_VPWR_c_386_n 0.00488573f $X=1.815 $Y=1.985 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_M1009_g N_VPWR_c_386_n 0.00625765f $X=2.245 $Y=1.985 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_102_n N_VPWR_c_386_n 0.0024874f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_157 N_KAPWR_c_215_n N_X_M1002_d 5.48427e-19 $X=1.435 $Y=2.21 $X2=0 $Y2=0
cc_158 N_KAPWR_c_200_n N_X_M1008_d 5.62186e-19 $X=2.315 $Y=2.24 $X2=0 $Y2=0
cc_159 N_KAPWR_c_210_n N_X_c_269_n 4.19008e-19 $X=0.84 $Y=2.21 $X2=0 $Y2=0
cc_160 N_KAPWR_c_212_n N_X_c_269_n 0.0147812f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_161 N_KAPWR_c_215_n N_X_c_269_n 0.0198417f $X=1.435 $Y=2.21 $X2=0 $Y2=0
cc_162 N_KAPWR_c_218_n N_X_c_269_n 0.00191784f $X=1.725 $Y=2.21 $X2=0 $Y2=0
cc_163 N_KAPWR_c_203_n N_X_c_269_n 0.0189713f $X=0.69 $Y=2 $X2=0 $Y2=0
cc_164 N_KAPWR_M1007_s N_X_c_279_n 0.00433084f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_165 N_KAPWR_c_200_n N_X_c_279_n 0.004286f $X=2.315 $Y=2.24 $X2=0 $Y2=0
cc_166 N_KAPWR_c_212_n N_X_c_279_n 0.0153341f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_167 N_KAPWR_c_215_n N_X_c_279_n 0.00124502f $X=1.435 $Y=2.21 $X2=0 $Y2=0
cc_168 N_KAPWR_c_218_n N_X_c_279_n 0.00862108f $X=1.725 $Y=2.21 $X2=0 $Y2=0
cc_169 N_KAPWR_c_215_n N_X_c_283_n 0.00382166f $X=1.435 $Y=2.21 $X2=0 $Y2=0
cc_170 N_KAPWR_c_200_n N_X_c_313_n 0.0180484f $X=2.315 $Y=2.24 $X2=0 $Y2=0
cc_171 N_KAPWR_c_212_n N_X_c_313_n 0.0147764f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_172 N_KAPWR_c_218_n N_X_c_313_n 0.00202021f $X=1.725 $Y=2.21 $X2=0 $Y2=0
cc_173 N_KAPWR_c_238_p N_X_c_313_n 0.00822148f $X=2.46 $Y=1.93 $X2=0 $Y2=0
cc_174 N_KAPWR_M1009_s N_X_c_262_n 0.00323085f $X=2.32 $Y=1.485 $X2=0 $Y2=0
cc_175 N_KAPWR_c_200_n N_X_c_262_n 0.00733832f $X=2.315 $Y=2.24 $X2=0 $Y2=0
cc_176 N_KAPWR_c_238_p N_X_c_262_n 0.0182224f $X=2.46 $Y=1.93 $X2=0 $Y2=0
cc_177 N_KAPWR_c_200_n N_VPWR_c_387_n 0.00207699f $X=2.315 $Y=2.24 $X2=0 $Y2=0
cc_178 N_KAPWR_c_201_n N_VPWR_c_387_n 0.00135384f $X=0.55 $Y=2.21 $X2=0 $Y2=0
cc_179 N_KAPWR_c_212_n N_VPWR_c_387_n 0.0181657f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_180 N_KAPWR_c_215_n N_VPWR_c_387_n 0.00151667f $X=1.435 $Y=2.21 $X2=0 $Y2=0
cc_181 N_KAPWR_c_218_n N_VPWR_c_387_n 2.22823e-19 $X=1.725 $Y=2.21 $X2=0 $Y2=0
cc_182 N_KAPWR_c_203_n N_VPWR_c_387_n 0.0198218f $X=0.69 $Y=2 $X2=0 $Y2=0
cc_183 N_KAPWR_c_238_p N_VPWR_c_387_n 0.0185087f $X=2.46 $Y=1.93 $X2=0 $Y2=0
cc_184 N_KAPWR_M1006_d N_VPWR_c_386_n 0.00143931f $X=0.55 $Y=1.485 $X2=0 $Y2=0
cc_185 N_KAPWR_M1007_s N_VPWR_c_386_n 0.00113449f $X=1.46 $Y=1.485 $X2=0 $Y2=0
cc_186 N_KAPWR_M1009_s N_VPWR_c_386_n 0.00130485f $X=2.32 $Y=1.485 $X2=0 $Y2=0
cc_187 N_KAPWR_c_201_n N_VPWR_c_386_n 0.268806f $X=0.55 $Y=2.21 $X2=0 $Y2=0
cc_188 N_KAPWR_c_212_n N_VPWR_c_386_n 0.00273177f $X=1.58 $Y=2.225 $X2=0 $Y2=0
cc_189 N_KAPWR_c_203_n N_VPWR_c_386_n 0.0029759f $X=0.69 $Y=2 $X2=0 $Y2=0
cc_190 N_KAPWR_c_238_p N_VPWR_c_386_n 0.00263498f $X=2.46 $Y=1.93 $X2=0 $Y2=0
cc_191 N_X_c_257_n N_VGND_c_342_n 0.0162872f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_192 X N_VGND_c_343_n 6.74578e-19 $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_193 X N_VGND_c_344_n 0.0201078f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_194 N_X_c_256_n N_VGND_c_346_n 0.010662f $X=1.175 $Y=0.51 $X2=0 $Y2=0
cc_195 N_X_c_257_n N_VGND_c_346_n 0.00224999f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_196 N_X_c_257_n N_VGND_c_347_n 0.00461204f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_197 N_X_c_259_n N_VGND_c_347_n 0.0092385f $X=2.035 $Y=0.51 $X2=0 $Y2=0
cc_198 N_X_M1000_d N_VGND_c_350_n 0.0023797f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_199 N_X_M1004_d N_VGND_c_350_n 0.00244557f $X=1.895 $Y=0.235 $X2=0 $Y2=0
cc_200 N_X_c_256_n N_VGND_c_350_n 0.0105577f $X=1.175 $Y=0.51 $X2=0 $Y2=0
cc_201 N_X_c_257_n N_VGND_c_350_n 0.0121304f $X=1.905 $Y=0.82 $X2=0 $Y2=0
cc_202 N_X_c_259_n N_VGND_c_350_n 0.00930021f $X=2.035 $Y=0.51 $X2=0 $Y2=0
cc_203 X N_VGND_c_350_n 0.00223695f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_204 N_X_c_269_n N_VPWR_c_387_n 0.0143059f $X=1.17 $Y=2.165 $X2=0 $Y2=0
cc_205 N_X_c_279_n N_VPWR_c_387_n 0.00200542f $X=1.905 $Y=1.857 $X2=0 $Y2=0
cc_206 N_X_c_283_n N_VPWR_c_387_n 0.00128772f $X=1.39 $Y=1.857 $X2=0 $Y2=0
cc_207 N_X_c_313_n N_VPWR_c_387_n 0.0138731f $X=2.03 $Y=1.96 $X2=0 $Y2=0
cc_208 N_X_M1002_d N_VPWR_c_386_n 0.00121005f $X=1.03 $Y=1.485 $X2=0 $Y2=0
cc_209 N_X_M1008_d N_VPWR_c_386_n 0.00122755f $X=1.89 $Y=1.485 $X2=0 $Y2=0
cc_210 N_X_c_269_n N_VPWR_c_386_n 0.0021899f $X=1.17 $Y=2.165 $X2=0 $Y2=0
cc_211 N_X_c_313_n N_VPWR_c_386_n 0.00211614f $X=2.03 $Y=1.96 $X2=0 $Y2=0

* File: sky130_fd_sc_hd__decap_8.spice.pex
* Created: Thu Aug 27 14:13:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HD__DECAP_8%VGND 1 9 10 11 12 21 33 36
r22 35 36 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r23 33 35 0.445255 $w=8.22e-07 $l=3e-08 $layer=LI1_cond $X=3.42 $Y=0.385
+ $X2=3.45 $Y2=0.385
r24 30 36 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=3.45
+ $Y2=0
r25 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r26 23 26 0.262178 $w=1.396e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r27 20 29 7.51576 $w=1.396e-06 $l=8.6e-07 $layer=LI1_cond $X=1.55 $Y=0.645
+ $X2=0.69 $Y2=0.645
r28 19 21 8.47369 $w=1.49e-06 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.87
+ $X2=1.715 $Y2=1.87
r29 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.29 $X2=1.55 $Y2=1.29
r30 16 29 1.1361 $w=1.396e-06 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.69 $Y2=0.645
r31 16 26 2.62178 $w=1.396e-06 $l=3e-07 $layer=LI1_cond $X=0.56 $Y=0.645
+ $X2=0.26 $Y2=0.645
r32 15 19 32.8283 $w=1.49e-06 $l=9.9e-07 $layer=POLY_cond $X=0.56 $Y=1.87
+ $X2=1.55 $Y2=1.87
r33 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.56
+ $Y=1.29 $X2=0.56 $Y2=1.29
r34 12 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r35 12 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r36 11 20 2.92381 $w=1.396e-06 $l=3.40147e-07 $layer=LI1_cond $X=1.735 $Y=0.385
+ $X2=1.55 $Y2=0.645
r37 10 33 4.05283 $w=9.4e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=0.385
+ $X2=3.42 $Y2=0.385
r38 10 11 18.0404 $w=9.38e-07 $l=1.39e-06 $layer=LI1_cond $X=3.125 $Y=0.385
+ $X2=1.735 $Y2=0.385
r39 9 21 5.33186 $w=1.13e-06 $l=1.25e-07 $layer=POLY_cond $X=1.84 $Y=2.05
+ $X2=1.715 $Y2=2.05
r40 1 33 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=3.285 $Y=0.235
+ $X2=3.42 $Y2=0.475
r41 1 26 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HD__DECAP_8%VPWR 1 9 10 11 12 17 19 30 33
r23 32 33 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r24 30 32 0.215041 $w=1.702e-06 $l=3e-08 $layer=LI1_cond $X=3.42 $Y=1.915
+ $X2=3.45 $Y2=1.915
r25 23 26 0.323894 $w=1.13e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=2.175
+ $X2=0.26 $Y2=2.175
r26 20 30 2.15041 $w=1.702e-06 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.915
+ $X2=3.42 $Y2=1.915
r27 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.11 $X2=3.12 $Y2=1.11
r28 16 20 7.38308 $w=1.702e-06 $l=1.03e-06 $layer=LI1_cond $X=2.09 $Y=1.915
+ $X2=3.12 $Y2=1.915
r29 15 19 45.2647 $w=1.17e-06 $l=1.03e-06 $layer=POLY_cond $X=2.09 $Y=0.69
+ $X2=3.12 $Y2=0.69
r30 15 17 12.167 $w=1.17e-06 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=0.69
+ $X2=1.925 $Y2=0.69
r31 15 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.09
+ $Y=1.11 $X2=2.09 $Y2=1.11
r32 12 33 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r33 12 23 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r34 11 26 4.56277 $w=1.26e-06 $l=4.55e-07 $layer=LI1_cond $X=0.715 $Y=2.175
+ $X2=0.26 $Y2=2.175
r35 10 16 2.17397 $w=1.702e-06 $l=3.40147e-07 $layer=LI1_cond $X=1.905 $Y=2.175
+ $X2=2.09 $Y2=1.915
r36 10 11 11.5222 $w=1.258e-06 $l=1.19e-06 $layer=LI1_cond $X=1.905 $Y=2.175
+ $X2=0.715 $Y2=2.175
r37 9 17 5.05802 $w=8.1e-07 $l=8.5e-08 $layer=POLY_cond $X=1.84 $Y=0.51
+ $X2=1.925 $Y2=0.51
r38 1 30 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.615 $X2=3.42 $Y2=1.83
r39 1 26 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends


* File: sky130_fd_sc_hd__o2bb2a_2.pxi.spice
* Created: Thu Aug 27 14:38:20 2020
* 
x_PM_SKY130_FD_SC_HD__O2BB2A_2%A_84_21# N_A_84_21#_M1013_s N_A_84_21#_M1009_d
+ N_A_84_21#_c_79_n N_A_84_21#_M1000_g N_A_84_21#_M1002_g N_A_84_21#_c_80_n
+ N_A_84_21#_M1004_g N_A_84_21#_M1010_g N_A_84_21#_c_81_n N_A_84_21#_c_82_n
+ N_A_84_21#_c_91_n N_A_84_21#_c_92_n N_A_84_21#_c_143_p N_A_84_21#_c_93_n
+ N_A_84_21#_c_83_n N_A_84_21#_c_84_n N_A_84_21#_c_85_n N_A_84_21#_c_86_n
+ N_A_84_21#_c_110_p PM_SKY130_FD_SC_HD__O2BB2A_2%A_84_21#
x_PM_SKY130_FD_SC_HD__O2BB2A_2%A1_N N_A1_N_M1003_g N_A1_N_M1001_g A1_N
+ N_A1_N_c_195_n PM_SKY130_FD_SC_HD__O2BB2A_2%A1_N
x_PM_SKY130_FD_SC_HD__O2BB2A_2%A2_N N_A2_N_M1007_g N_A2_N_M1006_g N_A2_N_c_232_n
+ N_A2_N_c_233_n A2_N N_A2_N_c_235_n PM_SKY130_FD_SC_HD__O2BB2A_2%A2_N
x_PM_SKY130_FD_SC_HD__O2BB2A_2%A_295_369# N_A_295_369#_M1007_d
+ N_A_295_369#_M1001_d N_A_295_369#_M1009_g N_A_295_369#_M1013_g
+ N_A_295_369#_c_280_n N_A_295_369#_c_281_n N_A_295_369#_c_282_n
+ N_A_295_369#_c_276_n N_A_295_369#_c_283_n N_A_295_369#_c_277_n
+ PM_SKY130_FD_SC_HD__O2BB2A_2%A_295_369#
x_PM_SKY130_FD_SC_HD__O2BB2A_2%B2 N_B2_M1005_g N_B2_M1012_g N_B2_c_343_n
+ N_B2_c_344_n B2 PM_SKY130_FD_SC_HD__O2BB2A_2%B2
x_PM_SKY130_FD_SC_HD__O2BB2A_2%B1 N_B1_M1008_g N_B1_M1011_g B1 B1 N_B1_c_394_n
+ PM_SKY130_FD_SC_HD__O2BB2A_2%B1
x_PM_SKY130_FD_SC_HD__O2BB2A_2%VPWR N_VPWR_M1002_s N_VPWR_M1010_s N_VPWR_M1006_d
+ N_VPWR_M1011_d N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ N_VPWR_c_424_n VPWR N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n
+ N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_419_n VPWR
+ PM_SKY130_FD_SC_HD__O2BB2A_2%VPWR
x_PM_SKY130_FD_SC_HD__O2BB2A_2%X N_X_M1000_s N_X_M1002_d N_X_c_482_n N_X_c_484_n
+ N_X_c_487_n N_X_c_480_n X N_X_c_497_n PM_SKY130_FD_SC_HD__O2BB2A_2%X
x_PM_SKY130_FD_SC_HD__O2BB2A_2%VGND N_VGND_M1000_d N_VGND_M1004_d N_VGND_M1005_d
+ N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n VGND
+ N_VGND_c_515_n N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n
+ N_VGND_c_520_n VGND PM_SKY130_FD_SC_HD__O2BB2A_2%VGND
x_PM_SKY130_FD_SC_HD__O2BB2A_2%A_581_47# N_A_581_47#_M1013_d N_A_581_47#_M1008_d
+ N_A_581_47#_c_573_n N_A_581_47#_c_574_n N_A_581_47#_c_575_n
+ N_A_581_47#_c_576_n PM_SKY130_FD_SC_HD__O2BB2A_2%A_581_47#
cc_1 VNB N_A_84_21#_c_79_n 0.0208627f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.995
cc_2 VNB N_A_84_21#_c_80_n 0.0167644f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.995
cc_3 VNB N_A_84_21#_c_81_n 0.00209149f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.16
cc_4 VNB N_A_84_21#_c_82_n 0.0502309f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.16
cc_5 VNB N_A_84_21#_c_83_n 0.00151591f $X=-0.19 $Y=-0.24 $X2=2.62 $Y2=0.485
cc_6 VNB N_A_84_21#_c_84_n 0.00319233f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=1.075
cc_7 VNB N_A_84_21#_c_85_n 0.00159184f $X=-0.19 $Y=-0.24 $X2=2.705 $Y2=1.245
cc_8 VNB N_A_84_21#_c_86_n 5.1593e-19 $X=-0.19 $Y=-0.24 $X2=2.907 $Y2=1.495
cc_9 VNB N_A1_N_M1003_g 0.0304792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A1_N 0.00882155f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_11 VNB N_A1_N_c_195_n 0.0219031f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_A2_N_M1006_g 0.0118112f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_N_c_232_n 0.0072395f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_14 VNB N_A2_N_c_233_n 0.0335408f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_15 VNB A2_N 0.00143774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_N_c_235_n 0.0203224f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_17 VNB N_A_295_369#_M1013_g 0.0518037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_295_369#_c_276_n 0.00379932f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.445
cc_19 VNB N_A_295_369#_c_277_n 0.0146576f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=0.69
cc_20 VNB N_B2_M1005_g 0.0262372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B2_c_343_n 0.00537183f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_22 VNB N_B2_c_344_n 0.0190068f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_23 VNB N_B1_M1008_g 0.0353013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB B1 0.00879609f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_25 VNB N_B1_c_394_n 0.03661f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_26 VNB N_VPWR_c_419_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_480_n 0.00103298f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_28 VNB N_VGND_c_511_n 0.0106114f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_29 VNB N_VGND_c_512_n 0.0341371f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_30 VNB N_VGND_c_513_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_31 VNB N_VGND_c_514_n 0.00468754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_515_n 0.0188517f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.16
cc_33 VNB N_VGND_c_516_n 0.0578945f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.97
cc_34 VNB N_VGND_c_517_n 0.0177197f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.53
cc_35 VNB N_VGND_c_518_n 0.226346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_519_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.657 $Y2=0.69
cc_37 VNB N_VGND_c_520_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=2.907 $Y2=1.97
cc_38 VNB N_A_581_47#_c_573_n 4.9051e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=0.56
cc_39 VNB N_A_581_47#_c_574_n 0.0168418f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_40 VNB N_A_581_47#_c_575_n 0.00324178f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_41 VNB N_A_581_47#_c_576_n 0.0161609f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=0.56
cc_42 VPB N_A_84_21#_M1002_g 0.0233526f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_43 VPB N_A_84_21#_M1010_g 0.0182799f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.985
cc_44 VPB N_A_84_21#_c_81_n 0.00141115f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_45 VPB N_A_84_21#_c_82_n 0.00822284f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_46 VPB N_A_84_21#_c_91_n 0.00184058f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.885
cc_47 VPB N_A_84_21#_c_92_n 0.00634457f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.97
cc_48 VPB N_A_84_21#_c_93_n 0.00654296f $X=-0.19 $Y=1.305 $X2=1.185 $Y2=1.53
cc_49 VPB N_A_84_21#_c_86_n 4.37229e-19 $X=-0.19 $Y=1.305 $X2=2.907 $Y2=1.495
cc_50 VPB N_A1_N_M1001_g 0.0414746f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_51 VPB N_A1_N_c_195_n 0.00437623f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_52 VPB N_A2_N_M1006_g 0.0429188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_295_369#_M1009_g 0.0207759f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.56
cc_54 VPB N_A_295_369#_M1013_g 0.00303362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_295_369#_c_280_n 0.0502441f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_56 VPB N_A_295_369#_c_281_n 0.0122806f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_57 VPB N_A_295_369#_c_282_n 0.00950066f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.325
cc_58 VPB N_A_295_369#_c_283_n 0.00803733f $X=-0.19 $Y=1.305 $X2=2.63 $Y2=1.97
cc_59 VPB N_A_295_369#_c_277_n 8.54583e-19 $X=-0.19 $Y=1.305 $X2=2.695 $Y2=0.69
cc_60 VPB N_B2_M1012_g 0.0364124f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_61 VPB N_B2_c_343_n 0.00156391f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.56
cc_62 VPB N_B2_c_344_n 0.0048081f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_63 VPB B2 0.00908182f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.995
cc_64 VPB N_B1_M1011_g 0.0483158f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.995
cc_65 VPB B1 0.0161504f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=0.56
cc_66 VPB N_B1_c_394_n 0.00982204f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_67 VPB N_VPWR_c_420_n 0.0105855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_421_n 0.0490186f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_69 VPB N_VPWR_c_422_n 0.00272569f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.445
cc_70 VPB N_VPWR_c_423_n 0.0101104f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.16
cc_71 VPB N_VPWR_c_424_n 0.0307945f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_425_n 0.015316f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.97
cc_73 VPB N_VPWR_c_426_n 0.0240162f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_427_n 0.0303387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_428_n 0.00507288f $X=-0.19 $Y=1.305 $X2=2.907 $Y2=2
cc_76 VPB N_VPWR_c_429_n 0.0138739f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_77 VPB N_VPWR_c_419_n 0.0438146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_X_c_480_n 9.41025e-19 $X=-0.19 $Y=1.305 $X2=0.915 $Y2=0.56
cc_79 N_A_84_21#_c_80_n N_A1_N_M1003_g 0.0187727f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_84_21#_M1010_g N_A1_N_M1001_g 0.0348015f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_81 N_A_84_21#_c_81_n N_A1_N_M1001_g 0.00222807f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_84_21#_c_91_n N_A1_N_M1001_g 0.00415725f $X=1.185 $Y=1.885 $X2=0 $Y2=0
cc_83 N_A_84_21#_c_92_n N_A1_N_M1001_g 0.0138792f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_84 N_A_84_21#_c_93_n N_A1_N_M1001_g 0.002419f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_85 N_A_84_21#_c_81_n A1_N 0.0154755f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_82_n A1_N 0.00140069f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_92_n A1_N 0.00353597f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_93_n A1_N 0.00419335f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_89 N_A_84_21#_c_81_n N_A1_N_c_195_n 0.00102065f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_82_n N_A1_N_c_195_n 0.0223879f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_92_n N_A2_N_M1006_g 0.0171337f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_92_n N_A_295_369#_M1001_d 0.00853544f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_93 N_A_84_21#_c_92_n N_A_295_369#_M1009_g 0.0147182f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_94 N_A_84_21#_c_110_p N_A_295_369#_M1009_g 0.0115099f $X=3.02 $Y=2 $X2=0
+ $Y2=0
cc_95 N_A_84_21#_c_83_n N_A_295_369#_M1013_g 0.00467857f $X=2.62 $Y=0.485 $X2=0
+ $Y2=0
cc_96 N_A_84_21#_c_84_n N_A_295_369#_M1013_g 0.0105368f $X=2.705 $Y=1.075 $X2=0
+ $Y2=0
cc_97 N_A_84_21#_c_85_n N_A_295_369#_M1013_g 0.00576018f $X=2.705 $Y=1.245 $X2=0
+ $Y2=0
cc_98 N_A_84_21#_c_86_n N_A_295_369#_M1013_g 0.00326592f $X=2.907 $Y=1.495 $X2=0
+ $Y2=0
cc_99 N_A_84_21#_c_92_n N_A_295_369#_c_280_n 0.0140966f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_100 N_A_84_21#_c_83_n N_A_295_369#_c_280_n 0.00182253f $X=2.62 $Y=0.485 $X2=0
+ $Y2=0
cc_101 N_A_84_21#_c_85_n N_A_295_369#_c_280_n 6.14215e-19 $X=2.705 $Y=1.245
+ $X2=0 $Y2=0
cc_102 N_A_84_21#_c_86_n N_A_295_369#_c_280_n 0.00572493f $X=2.907 $Y=1.495
+ $X2=0 $Y2=0
cc_103 N_A_84_21#_c_92_n N_A_295_369#_c_281_n 0.011155f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_104 N_A_84_21#_c_86_n N_A_295_369#_c_281_n 0.00343895f $X=2.907 $Y=1.495
+ $X2=0 $Y2=0
cc_105 N_A_84_21#_c_91_n N_A_295_369#_c_282_n 0.00791067f $X=1.185 $Y=1.885
+ $X2=0 $Y2=0
cc_106 N_A_84_21#_c_92_n N_A_295_369#_c_282_n 0.0492496f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_107 N_A_84_21#_c_93_n N_A_295_369#_c_282_n 0.0100855f $X=1.185 $Y=1.53 $X2=0
+ $Y2=0
cc_108 N_A_84_21#_c_83_n N_A_295_369#_c_276_n 0.0140331f $X=2.62 $Y=0.485 $X2=0
+ $Y2=0
cc_109 N_A_84_21#_c_92_n N_A_295_369#_c_283_n 0.0214628f $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_110 N_A_84_21#_c_86_n N_A_295_369#_c_283_n 0.0269621f $X=2.907 $Y=1.495 $X2=0
+ $Y2=0
cc_111 N_A_84_21#_c_83_n N_A_295_369#_c_277_n 0.00951375f $X=2.62 $Y=0.485 $X2=0
+ $Y2=0
cc_112 N_A_84_21#_c_84_n N_A_295_369#_c_277_n 0.0324162f $X=2.705 $Y=1.075 $X2=0
+ $Y2=0
cc_113 N_A_84_21#_c_86_n N_A_295_369#_c_277_n 0.0060268f $X=2.907 $Y=1.495 $X2=0
+ $Y2=0
cc_114 N_A_84_21#_c_83_n N_B2_M1005_g 2.90542e-19 $X=2.62 $Y=0.485 $X2=0 $Y2=0
cc_115 N_A_84_21#_c_84_n N_B2_M1005_g 4.42792e-19 $X=2.705 $Y=1.075 $X2=0 $Y2=0
cc_116 N_A_84_21#_c_92_n N_B2_M1012_g 0.00929249f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_117 N_A_84_21#_c_86_n N_B2_M1012_g 5.23107e-19 $X=2.907 $Y=1.495 $X2=0 $Y2=0
cc_118 N_A_84_21#_c_110_p N_B2_M1012_g 0.0034236f $X=3.02 $Y=2 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_92_n N_B2_c_343_n 0.0182474f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_120 N_A_84_21#_c_85_n N_B2_c_343_n 0.0197242f $X=2.705 $Y=1.245 $X2=0 $Y2=0
cc_121 N_A_84_21#_c_92_n N_B2_c_344_n 0.00139774f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_122 N_A_84_21#_c_84_n N_B2_c_344_n 4.2387e-19 $X=2.705 $Y=1.075 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_85_n N_B2_c_344_n 2.01387e-19 $X=2.705 $Y=1.245 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_92_n B2 0.0498524f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_86_n B2 0.00491462f $X=2.907 $Y=1.495 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_91_n N_VPWR_M1010_s 0.00409302f $X=1.185 $Y=1.885 $X2=0
+ $Y2=0
cc_127 N_A_84_21#_c_143_p N_VPWR_M1010_s 0.00409058f $X=1.27 $Y=1.97 $X2=0 $Y2=0
cc_128 N_A_84_21#_c_93_n N_VPWR_M1010_s 0.00204498f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_92_n N_VPWR_M1006_d 0.0182075f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_130 N_A_84_21#_M1002_g N_VPWR_c_421_n 0.00475737f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_A_84_21#_M1002_g N_VPWR_c_422_n 4.81859e-19 $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_84_21#_M1010_g N_VPWR_c_422_n 0.00747419f $X=0.915 $Y=1.985 $X2=0
+ $Y2=0
cc_133 N_A_84_21#_c_143_p N_VPWR_c_422_n 0.0131715f $X=1.27 $Y=1.97 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_93_n N_VPWR_c_422_n 0.00236443f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_135 N_A_84_21#_M1002_g N_VPWR_c_425_n 0.00533769f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_136 N_A_84_21#_M1010_g N_VPWR_c_425_n 0.0046653f $X=0.915 $Y=1.985 $X2=0
+ $Y2=0
cc_137 N_A_84_21#_c_92_n N_VPWR_c_426_n 0.0124071f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_138 N_A_84_21#_c_92_n N_VPWR_c_427_n 0.00410636f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_139 N_A_84_21#_c_110_p N_VPWR_c_427_n 0.0161955f $X=3.02 $Y=2 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_92_n N_VPWR_c_429_n 0.0295056f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_110_p N_VPWR_c_429_n 0.0105582f $X=3.02 $Y=2 $X2=0 $Y2=0
cc_142 N_A_84_21#_M1009_d N_VPWR_c_419_n 0.00233757f $X=2.885 $Y=1.845 $X2=0
+ $Y2=0
cc_143 N_A_84_21#_M1002_g N_VPWR_c_419_n 0.0103065f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_144 N_A_84_21#_M1010_g N_VPWR_c_419_n 0.00789179f $X=0.915 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_84_21#_c_92_n N_VPWR_c_419_n 0.031758f $X=2.63 $Y=1.97 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_143_p N_VPWR_c_419_n 7.95799e-19 $X=1.27 $Y=1.97 $X2=0 $Y2=0
cc_147 N_A_84_21#_c_110_p N_VPWR_c_419_n 0.0127238f $X=3.02 $Y=2 $X2=0 $Y2=0
cc_148 N_A_84_21#_c_79_n N_X_c_482_n 0.00483966f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_80_n N_X_c_482_n 0.00470742f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_84_21#_c_79_n N_X_c_484_n 0.00189307f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_84_21#_c_80_n N_X_c_484_n 0.00393368f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_82_n N_X_c_484_n 0.00194336f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_84_21#_M1002_g N_X_c_487_n 0.00143964f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_154 N_A_84_21#_c_82_n N_X_c_487_n 0.00144574f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_79_n N_X_c_480_n 0.00514632f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_84_21#_M1002_g N_X_c_480_n 0.01081f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_80_n N_X_c_480_n 0.00342125f $X=0.915 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_84_21#_M1010_g N_X_c_480_n 0.003123f $X=0.915 $Y=1.985 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_81_n N_X_c_480_n 0.0309161f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_84_21#_c_82_n N_X_c_480_n 0.024289f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_84_21#_c_91_n N_X_c_480_n 0.00699907f $X=1.185 $Y=1.885 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_93_n N_X_c_480_n 0.0126944f $X=1.185 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A_84_21#_M1002_g N_X_c_497_n 0.00642666f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_79_n N_VGND_c_512_n 0.00501374f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_84_21#_c_80_n N_VGND_c_513_n 0.00505437f $X=0.915 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_84_21#_c_82_n N_VGND_c_513_n 0.00118907f $X=0.96 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_84_21#_c_79_n N_VGND_c_515_n 0.00533769f $X=0.495 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_84_21#_c_80_n N_VGND_c_515_n 0.00541359f $X=0.915 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_84_21#_c_83_n N_VGND_c_516_n 0.010457f $X=2.62 $Y=0.485 $X2=0 $Y2=0
cc_170 N_A_84_21#_M1013_s N_VGND_c_518_n 0.00356607f $X=2.495 $Y=0.235 $X2=0
+ $Y2=0
cc_171 N_A_84_21#_c_79_n N_VGND_c_518_n 0.0103065f $X=0.495 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_80_n N_VGND_c_518_n 0.00981417f $X=0.915 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_84_21#_c_83_n N_VGND_c_518_n 0.00887248f $X=2.62 $Y=0.485 $X2=0 $Y2=0
cc_174 N_A_84_21#_c_83_n N_A_581_47#_c_573_n 0.0167089f $X=2.62 $Y=0.485 $X2=0
+ $Y2=0
cc_175 N_A_84_21#_c_92_n N_A_581_47#_c_575_n 5.82402e-19 $X=2.63 $Y=1.97 $X2=0
+ $Y2=0
cc_176 N_A_84_21#_c_84_n N_A_581_47#_c_575_n 0.0142077f $X=2.705 $Y=1.075 $X2=0
+ $Y2=0
cc_177 N_A1_N_M1001_g N_A2_N_M1006_g 0.0403258f $X=1.4 $Y=2.165 $X2=0 $Y2=0
cc_178 A1_N N_A2_N_M1006_g 0.00181076f $X=1.515 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A1_N_c_195_n N_A2_N_M1006_g 0.00881312f $X=1.44 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A1_N_M1003_g N_A2_N_c_232_n 0.00427327f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_181 A1_N N_A2_N_c_232_n 0.0158717f $X=1.515 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A1_N_c_195_n N_A2_N_c_232_n 0.00203454f $X=1.44 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A1_N_c_195_n N_A2_N_c_233_n 0.00687752f $X=1.44 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A1_N_M1003_g A2_N 0.00205785f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A1_N_M1003_g N_A2_N_c_235_n 0.031774f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A1_N_M1001_g N_A_295_369#_c_282_n 0.00676621f $X=1.4 $Y=2.165 $X2=0
+ $Y2=0
cc_187 A1_N N_A_295_369#_c_282_n 0.0150276f $X=1.515 $Y=1.105 $X2=0 $Y2=0
cc_188 N_A1_N_c_195_n N_A_295_369#_c_282_n 0.00231747f $X=1.44 $Y=1.16 $X2=0
+ $Y2=0
cc_189 A1_N N_A_295_369#_c_277_n 0.00659601f $X=1.515 $Y=1.105 $X2=0 $Y2=0
cc_190 N_A1_N_M1001_g N_VPWR_c_422_n 0.00433972f $X=1.4 $Y=2.165 $X2=0 $Y2=0
cc_191 N_A1_N_M1001_g N_VPWR_c_426_n 0.00429465f $X=1.4 $Y=2.165 $X2=0 $Y2=0
cc_192 N_A1_N_M1001_g N_VPWR_c_419_n 0.0063007f $X=1.4 $Y=2.165 $X2=0 $Y2=0
cc_193 N_A1_N_M1003_g N_X_c_482_n 3.76466e-19 $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A1_N_M1003_g N_VGND_c_513_n 0.00767959f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_195 A1_N N_VGND_c_513_n 9.9771e-19 $X=1.515 $Y=1.105 $X2=0 $Y2=0
cc_196 N_A1_N_M1003_g N_VGND_c_516_n 0.00585385f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A1_N_M1003_g N_VGND_c_518_n 0.0110899f $X=1.395 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A2_N_M1006_g N_A_295_369#_M1009_g 0.011473f $X=1.95 $Y=2.165 $X2=0
+ $Y2=0
cc_199 N_A2_N_c_233_n N_A_295_369#_M1013_g 0.00328794f $X=1.94 $Y=0.935 $X2=0
+ $Y2=0
cc_200 N_A2_N_M1006_g N_A_295_369#_c_280_n 0.0200293f $X=1.95 $Y=2.165 $X2=0
+ $Y2=0
cc_201 N_A2_N_M1006_g N_A_295_369#_c_282_n 0.0133765f $X=1.95 $Y=2.165 $X2=0
+ $Y2=0
cc_202 N_A2_N_c_232_n N_A_295_369#_c_282_n 0.0116307f $X=1.625 $Y=0.905 $X2=0
+ $Y2=0
cc_203 N_A2_N_c_233_n N_A_295_369#_c_282_n 0.00329605f $X=1.94 $Y=0.935 $X2=0
+ $Y2=0
cc_204 N_A2_N_c_232_n N_A_295_369#_c_276_n 0.00673523f $X=1.625 $Y=0.905 $X2=0
+ $Y2=0
cc_205 N_A2_N_c_233_n N_A_295_369#_c_276_n 0.00226202f $X=1.94 $Y=0.935 $X2=0
+ $Y2=0
cc_206 N_A2_N_c_235_n N_A_295_369#_c_276_n 0.00259127f $X=1.93 $Y=0.77 $X2=0
+ $Y2=0
cc_207 N_A2_N_M1006_g N_A_295_369#_c_283_n 2.10865e-19 $X=1.95 $Y=2.165 $X2=0
+ $Y2=0
cc_208 N_A2_N_M1006_g N_A_295_369#_c_277_n 0.00975624f $X=1.95 $Y=2.165 $X2=0
+ $Y2=0
cc_209 N_A2_N_c_232_n N_A_295_369#_c_277_n 0.0273904f $X=1.625 $Y=0.905 $X2=0
+ $Y2=0
cc_210 N_A2_N_c_233_n N_A_295_369#_c_277_n 0.00373932f $X=1.94 $Y=0.935 $X2=0
+ $Y2=0
cc_211 A2_N N_A_295_369#_c_277_n 0.00470786f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_212 N_A2_N_c_235_n N_A_295_369#_c_277_n 0.00217843f $X=1.93 $Y=0.77 $X2=0
+ $Y2=0
cc_213 N_A2_N_M1006_g N_VPWR_c_426_n 0.00429465f $X=1.95 $Y=2.165 $X2=0 $Y2=0
cc_214 N_A2_N_M1006_g N_VPWR_c_429_n 0.0103051f $X=1.95 $Y=2.165 $X2=0 $Y2=0
cc_215 N_A2_N_M1006_g N_VPWR_c_419_n 0.00708152f $X=1.95 $Y=2.165 $X2=0 $Y2=0
cc_216 N_A2_N_c_232_n N_X_c_484_n 0.00222162f $X=1.625 $Y=0.905 $X2=0 $Y2=0
cc_217 N_A2_N_c_232_n N_VGND_c_513_n 8.49459e-19 $X=1.625 $Y=0.905 $X2=0 $Y2=0
cc_218 A2_N N_VGND_c_513_n 0.0110811f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_219 N_A2_N_c_232_n N_VGND_c_516_n 0.00236127f $X=1.625 $Y=0.905 $X2=0 $Y2=0
cc_220 A2_N N_VGND_c_516_n 0.00799532f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_221 N_A2_N_c_235_n N_VGND_c_516_n 0.0042834f $X=1.93 $Y=0.77 $X2=0 $Y2=0
cc_222 N_A2_N_c_232_n N_VGND_c_518_n 0.00411405f $X=1.625 $Y=0.905 $X2=0 $Y2=0
cc_223 A2_N N_VGND_c_518_n 0.00776053f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_224 N_A2_N_c_235_n N_VGND_c_518_n 0.0074896f $X=1.93 $Y=0.77 $X2=0 $Y2=0
cc_225 A2_N A_294_47# 0.00485199f $X=1.515 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_226 N_A_295_369#_M1013_g N_B2_M1005_g 0.0242003f $X=2.83 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_295_369#_M1009_g N_B2_M1012_g 0.0131603f $X=2.81 $Y=2.165 $X2=0 $Y2=0
cc_228 N_A_295_369#_M1013_g N_B2_M1012_g 0.0169755f $X=2.83 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A_295_369#_M1013_g N_B2_c_343_n 0.00167467f $X=2.83 $Y=0.445 $X2=0
+ $Y2=0
cc_230 N_A_295_369#_M1013_g N_B2_c_344_n 0.0197362f $X=2.83 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_295_369#_M1009_g N_VPWR_c_427_n 0.00409647f $X=2.81 $Y=2.165 $X2=0
+ $Y2=0
cc_232 N_A_295_369#_M1009_g N_VPWR_c_429_n 0.00653875f $X=2.81 $Y=2.165 $X2=0
+ $Y2=0
cc_233 N_A_295_369#_M1001_d N_VPWR_c_419_n 0.00484561f $X=1.475 $Y=1.845 $X2=0
+ $Y2=0
cc_234 N_A_295_369#_M1009_g N_VPWR_c_419_n 0.00655805f $X=2.81 $Y=2.165 $X2=0
+ $Y2=0
cc_235 N_A_295_369#_M1013_g N_VGND_c_516_n 0.00551068f $X=2.83 $Y=0.445 $X2=0
+ $Y2=0
cc_236 N_A_295_369#_c_276_n N_VGND_c_516_n 0.0152503f $X=2.195 $Y=0.48 $X2=0
+ $Y2=0
cc_237 N_A_295_369#_M1007_d N_VGND_c_518_n 0.00228556f $X=1.935 $Y=0.235 $X2=0
+ $Y2=0
cc_238 N_A_295_369#_M1013_g N_VGND_c_518_n 0.0113344f $X=2.83 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_295_369#_c_276_n N_VGND_c_518_n 0.0157351f $X=2.195 $Y=0.48 $X2=0
+ $Y2=0
cc_240 N_A_295_369#_M1013_g N_A_581_47#_c_573_n 4.98506e-19 $X=2.83 $Y=0.445
+ $X2=0 $Y2=0
cc_241 N_A_295_369#_M1013_g N_A_581_47#_c_575_n 0.00146399f $X=2.83 $Y=0.445
+ $X2=0 $Y2=0
cc_242 N_B2_M1005_g N_B1_M1008_g 0.0258966f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_243 N_B2_M1012_g N_B1_M1011_g 0.0501288f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_244 B2 N_B1_M1011_g 0.0104584f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_245 N_B2_c_343_n B1 0.0203467f $X=3.355 $Y=1.2 $X2=0 $Y2=0
cc_246 N_B2_c_344_n B1 2.04424e-19 $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_247 B2 B1 0.0235332f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_248 N_B2_c_343_n N_B1_c_394_n 0.00190925f $X=3.355 $Y=1.2 $X2=0 $Y2=0
cc_249 N_B2_c_344_n N_B1_c_394_n 0.0217078f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_250 N_B2_M1012_g N_VPWR_c_424_n 0.00150124f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_251 B2 N_VPWR_c_424_n 0.0388882f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_252 N_B2_M1012_g N_VPWR_c_427_n 0.00572216f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_253 B2 N_VPWR_c_427_n 0.00868579f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_254 N_B2_M1012_g N_VPWR_c_419_n 0.0105447f $X=3.25 $Y=2.165 $X2=0 $Y2=0
cc_255 B2 N_VPWR_c_419_n 0.00634211f $X=3.355 $Y=1.445 $X2=0 $Y2=0
cc_256 B2 A_665_369# 0.0111542f $X=3.355 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_257 N_B2_M1005_g N_VGND_c_514_n 0.00268723f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_258 N_B2_M1005_g N_VGND_c_516_n 0.00434819f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_259 N_B2_M1005_g N_VGND_c_518_n 0.00592382f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_260 N_B2_M1005_g N_A_581_47#_c_573_n 0.00569407f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_261 N_B2_M1005_g N_A_581_47#_c_574_n 0.00977346f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_262 N_B2_c_343_n N_A_581_47#_c_574_n 0.026246f $X=3.355 $Y=1.2 $X2=0 $Y2=0
cc_263 N_B2_c_344_n N_A_581_47#_c_574_n 0.00148047f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B2_M1005_g N_A_581_47#_c_575_n 0.0018717f $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_265 N_B2_c_343_n N_A_581_47#_c_575_n 0.0181026f $X=3.355 $Y=1.2 $X2=0 $Y2=0
cc_266 N_B2_c_344_n N_A_581_47#_c_575_n 0.0015306f $X=3.25 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B2_M1005_g N_A_581_47#_c_576_n 5.07436e-19 $X=3.25 $Y=0.445 $X2=0 $Y2=0
cc_268 N_B1_M1011_g N_VPWR_c_424_n 0.0136165f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_269 B1 N_VPWR_c_424_n 0.028818f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_270 N_B1_c_394_n N_VPWR_c_424_n 0.00111969f $X=3.865 $Y=1.16 $X2=0 $Y2=0
cc_271 N_B1_M1011_g N_VPWR_c_427_n 0.00525069f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_272 N_B1_M1011_g N_VPWR_c_419_n 0.00891732f $X=3.67 $Y=2.165 $X2=0 $Y2=0
cc_273 N_B1_M1008_g N_VGND_c_514_n 0.00268723f $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_274 N_B1_M1008_g N_VGND_c_517_n 0.00425893f $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_275 N_B1_M1008_g N_VGND_c_518_n 0.00677018f $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_276 N_B1_M1008_g N_A_581_47#_c_573_n 4.95296e-19 $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_277 N_B1_M1008_g N_A_581_47#_c_574_n 0.0164689f $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_278 B1 N_A_581_47#_c_574_n 0.0295892f $X=3.815 $Y=1.105 $X2=0 $Y2=0
cc_279 N_B1_c_394_n N_A_581_47#_c_574_n 0.0071376f $X=3.865 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B1_M1008_g N_A_581_47#_c_576_n 0.00766804f $X=3.67 $Y=0.445 $X2=0 $Y2=0
cc_281 N_VPWR_c_419_n N_X_M1002_d 0.0038878f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_421_n N_X_c_480_n 0.0401048f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_283 N_VPWR_c_425_n N_X_c_497_n 0.0154848f $X=0.96 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_419_n N_X_c_497_n 0.00951427f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_419_n A_665_369# 0.00572363f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_286 N_VPWR_c_421_n N_VGND_c_512_n 0.0111763f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_287 N_X_c_482_n N_VGND_c_512_n 0.0252065f $X=0.705 $Y=0.37 $X2=0 $Y2=0
cc_288 N_X_c_482_n N_VGND_c_513_n 0.0328814f $X=0.705 $Y=0.37 $X2=0 $Y2=0
cc_289 N_X_c_482_n N_VGND_c_515_n 0.0191504f $X=0.705 $Y=0.37 $X2=0 $Y2=0
cc_290 N_X_M1000_s N_VGND_c_518_n 0.00215201f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_291 N_X_c_482_n N_VGND_c_518_n 0.0123629f $X=0.705 $Y=0.37 $X2=0 $Y2=0
cc_292 N_VGND_c_518_n A_294_47# 0.00449915f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_293 N_VGND_c_518_n N_A_581_47#_M1013_d 0.00398008f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_294 N_VGND_c_518_n N_A_581_47#_M1008_d 0.00214228f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_c_516_n N_A_581_47#_c_573_n 0.00966659f $X=3.375 $Y=0 $X2=0 $Y2=0
cc_296 N_VGND_c_518_n N_A_581_47#_c_573_n 0.00839587f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_297 N_VGND_c_514_n N_A_581_47#_c_574_n 0.0128746f $X=3.46 $Y=0.39 $X2=0 $Y2=0
cc_298 N_VGND_c_516_n N_A_581_47#_c_574_n 0.00263328f $X=3.375 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_517_n N_A_581_47#_c_574_n 0.00236451f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_300 N_VGND_c_518_n N_A_581_47#_c_574_n 0.0087883f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_301 N_VGND_c_517_n N_A_581_47#_c_576_n 0.014713f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_302 N_VGND_c_518_n N_A_581_47#_c_576_n 0.0119488f $X=3.91 $Y=0 $X2=0 $Y2=0

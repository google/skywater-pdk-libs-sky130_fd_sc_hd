* File: sky130_fd_sc_hd__o22a_1.spice.SKY130_FD_SC_HD__O22A_1.pxi
* Created: Thu Aug 27 14:37:30 2020
* 
x_PM_SKY130_FD_SC_HD__O22A_1%A_78_199# N_A_78_199#_M1004_d N_A_78_199#_M1002_d
+ N_A_78_199#_c_53_n N_A_78_199#_M1008_g N_A_78_199#_M1003_g N_A_78_199#_c_54_n
+ N_A_78_199#_c_55_n N_A_78_199#_c_94_p N_A_78_199#_c_62_p N_A_78_199#_c_96_p
+ N_A_78_199#_c_63_p N_A_78_199#_c_64_p N_A_78_199#_c_56_n N_A_78_199#_c_57_n
+ PM_SKY130_FD_SC_HD__O22A_1%A_78_199#
x_PM_SKY130_FD_SC_HD__O22A_1%B1 N_B1_M1006_g N_B1_c_125_n N_B1_M1004_g B1
+ N_B1_c_127_n PM_SKY130_FD_SC_HD__O22A_1%B1
x_PM_SKY130_FD_SC_HD__O22A_1%B2 N_B2_M1002_g N_B2_c_158_n N_B2_M1001_g B2
+ N_B2_c_159_n N_B2_c_160_n B2 PM_SKY130_FD_SC_HD__O22A_1%B2
x_PM_SKY130_FD_SC_HD__O22A_1%A2 N_A2_M1000_g N_A2_M1007_g N_A2_c_194_n
+ N_A2_c_195_n A2 N_A2_c_196_n PM_SKY130_FD_SC_HD__O22A_1%A2
x_PM_SKY130_FD_SC_HD__O22A_1%A1 N_A1_M1005_g N_A1_M1009_g A1 N_A1_c_238_n
+ N_A1_c_239_n PM_SKY130_FD_SC_HD__O22A_1%A1
x_PM_SKY130_FD_SC_HD__O22A_1%X N_X_M1008_s N_X_M1003_s X N_X_c_262_n
+ PM_SKY130_FD_SC_HD__O22A_1%X
x_PM_SKY130_FD_SC_HD__O22A_1%VPWR N_VPWR_M1003_d N_VPWR_M1009_d N_VPWR_c_276_n
+ N_VPWR_c_277_n VPWR N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n
+ N_VPWR_c_275_n PM_SKY130_FD_SC_HD__O22A_1%VPWR
x_PM_SKY130_FD_SC_HD__O22A_1%VGND N_VGND_M1008_d N_VGND_M1000_d N_VGND_c_320_n
+ N_VGND_c_321_n N_VGND_c_322_n VGND N_VGND_c_323_n N_VGND_c_324_n
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n PM_SKY130_FD_SC_HD__O22A_1%VGND
x_PM_SKY130_FD_SC_HD__O22A_1%A_215_47# N_A_215_47#_M1004_s N_A_215_47#_M1001_d
+ N_A_215_47#_M1005_d N_A_215_47#_c_369_n N_A_215_47#_c_382_n
+ N_A_215_47#_c_376_n N_A_215_47#_c_370_n N_A_215_47#_c_371_n
+ PM_SKY130_FD_SC_HD__O22A_1%A_215_47#
cc_1 VNB N_A_78_199#_c_53_n 0.0230649f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_78_199#_c_54_n 0.00137788f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_3 VNB N_A_78_199#_c_55_n 0.034971f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.16
cc_4 VNB N_A_78_199#_c_56_n 0.00255278f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.73
cc_5 VNB N_A_78_199#_c_57_n 0.00940817f $X=-0.19 $Y=-0.24 $X2=1.42 $Y2=0.77
cc_6 VNB N_B1_c_125_n 0.0200849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB B1 0.00189861f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB N_B1_c_127_n 0.03071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B2_c_158_n 0.0171375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B2_c_159_n 0.0195481f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_11 VNB N_B2_c_160_n 0.00465685f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_12 VNB N_A2_c_194_n 0.00334867f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_13 VNB N_A2_c_195_n 0.020301f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_14 VNB N_A2_c_196_n 0.0172054f $X=-0.19 $Y=-0.24 $X2=0.672 $Y2=1.495
cc_15 VNB A1 0.0114652f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_A1_c_238_n 0.0309602f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_17 VNB N_A1_c_239_n 0.0222254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_262_n 0.0423323f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_19 VNB N_VPWR_c_275_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_320_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_VGND_c_321_n 0.0411704f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.985
cc_22 VNB N_VGND_c_322_n 0.00463598f $X=-0.19 $Y=-0.24 $X2=0.672 $Y2=1.495
cc_23 VNB N_VGND_c_323_n 0.0187447f $X=-0.19 $Y=-0.24 $X2=1.42 $Y2=0.805
cc_24 VNB N_VGND_c_324_n 0.0173701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_325_n 0.183722f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.77
cc_26 VNB N_VGND_c_326_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_327_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.16
cc_28 VNB N_A_215_47#_c_369_n 0.00241395f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.325
cc_29 VNB N_A_215_47#_c_370_n 0.00773281f $X=-0.19 $Y=-0.24 $X2=0.672 $Y2=1.16
cc_30 VNB N_A_215_47#_c_371_n 0.016608f $X=-0.19 $Y=-0.24 $X2=0.81 $Y2=0.805
cc_31 VPB N_A_78_199#_M1003_g 0.0256068f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_32 VPB N_A_78_199#_c_54_n 0.00217762f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_33 VPB N_A_78_199#_c_55_n 0.0104282f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.16
cc_34 VPB N_B1_M1006_g 0.022011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB B1 0.00315795f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_36 VPB N_B1_c_127_n 0.0100029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B2_M1002_g 0.0206829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_B2_c_159_n 0.00393786f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_39 VPB N_B2_c_160_n 0.00201087f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_40 VPB N_A2_M1007_g 0.0184111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A2_c_194_n 0.0115851f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_42 VPB N_A2_c_195_n 0.00497124f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_43 VPB N_A1_M1009_g 0.0242019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A1_c_238_n 0.00655583f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_45 VPB N_X_c_262_n 0.0473378f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.325
cc_46 VPB N_VPWR_c_276_n 0.0099172f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_47 VPB N_VPWR_c_277_n 0.0452565f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_48 VPB N_VPWR_c_278_n 0.0161648f $X=-0.19 $Y=1.305 $X2=0.672 $Y2=1.495
cc_49 VPB N_VPWR_c_279_n 0.0393907f $X=-0.19 $Y=1.305 $X2=0.81 $Y2=0.805
cc_50 VPB N_VPWR_c_280_n 0.0153853f $X=-0.19 $Y=1.305 $X2=1.42 $Y2=0.77
cc_51 VPB N_VPWR_c_275_n 0.0430347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A_78_199#_c_54_n N_B1_M1006_g 0.0043364f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_78_199#_c_62_p N_B1_M1006_g 0.0195776f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_54 N_A_78_199#_c_63_p N_B1_M1006_g 5.92605e-19 $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_55 N_A_78_199#_c_64_p N_B1_M1006_g 0.0023078f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_56 N_A_78_199#_c_54_n N_B1_c_125_n 0.00247681f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_78_199#_c_56_n N_B1_c_125_n 0.0069705f $X=1.62 $Y=0.73 $X2=0 $Y2=0
cc_58 N_A_78_199#_c_57_n N_B1_c_125_n 0.00931075f $X=1.42 $Y=0.77 $X2=0 $Y2=0
cc_59 N_A_78_199#_c_54_n B1 0.0196416f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_78_199#_c_55_n B1 0.00151421f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_78_199#_c_62_p B1 0.0240683f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_62 N_A_78_199#_c_57_n B1 0.0253303f $X=1.42 $Y=0.77 $X2=0 $Y2=0
cc_63 N_A_78_199#_c_54_n N_B1_c_127_n 8.39646e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_78_199#_c_55_n N_B1_c_127_n 0.0216064f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_78_199#_c_62_p N_B1_c_127_n 0.00183798f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_66 N_A_78_199#_c_57_n N_B1_c_127_n 0.00746472f $X=1.42 $Y=0.77 $X2=0 $Y2=0
cc_67 N_A_78_199#_c_62_p N_B2_M1002_g 0.00514666f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_68 N_A_78_199#_c_63_p N_B2_M1002_g 0.00619177f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_69 N_A_78_199#_c_64_p N_B2_M1002_g 0.014681f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_70 N_A_78_199#_c_56_n N_B2_c_158_n 0.00385556f $X=1.62 $Y=0.73 $X2=0 $Y2=0
cc_71 N_A_78_199#_c_63_p N_B2_c_159_n 0.00285844f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_72 N_A_78_199#_c_56_n N_B2_c_159_n 0.00173935f $X=1.62 $Y=0.73 $X2=0 $Y2=0
cc_73 N_A_78_199#_c_62_p N_B2_c_160_n 0.0134392f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_74 N_A_78_199#_c_63_p N_B2_c_160_n 0.018278f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_75 N_A_78_199#_c_56_n N_B2_c_160_n 0.0190747f $X=1.62 $Y=0.73 $X2=0 $Y2=0
cc_76 N_A_78_199#_c_63_p N_A2_M1007_g 0.00245076f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_77 N_A_78_199#_c_64_p N_A2_M1007_g 0.0072191f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_78 N_A_78_199#_c_63_p N_A2_c_194_n 0.00995938f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_79 N_A_78_199#_c_63_p A2 0.00957118f $X=1.927 $Y=1.805 $X2=0 $Y2=0
cc_80 N_A_78_199#_c_64_p A2 0.0276688f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_81 N_A_78_199#_c_53_n N_X_c_262_n 0.00506422f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_78_199#_M1003_g N_X_c_262_n 0.00356334f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_83 N_A_78_199#_c_54_n N_X_c_262_n 0.0456507f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_78_199#_c_55_n N_X_c_262_n 0.00942681f $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_78_199#_c_94_p N_X_c_262_n 0.00794912f $X=0.81 $Y=0.805 $X2=0 $Y2=0
cc_86 N_A_78_199#_c_62_p N_VPWR_M1003_d 0.0137578f $X=1.735 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_78_199#_c_96_p N_VPWR_M1003_d 0.00278894f $X=0.81 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_78_199#_M1003_g N_VPWR_c_278_n 0.00546359f $X=0.49 $Y=1.985 $X2=0
+ $Y2=0
cc_89 N_A_78_199#_c_64_p N_VPWR_c_279_n 0.0246809f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_90 N_A_78_199#_M1003_g N_VPWR_c_280_n 0.0128077f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_78_199#_c_55_n N_VPWR_c_280_n 8.32196e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_78_199#_c_62_p N_VPWR_c_280_n 0.0387238f $X=1.735 $Y=1.6 $X2=0 $Y2=0
cc_93 N_A_78_199#_c_96_p N_VPWR_c_280_n 0.0176249f $X=0.81 $Y=1.6 $X2=0 $Y2=0
cc_94 N_A_78_199#_c_64_p N_VPWR_c_280_n 0.0240363f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_95 N_A_78_199#_M1002_d N_VPWR_c_275_n 0.0105888f $X=1.845 $Y=1.485 $X2=0
+ $Y2=0
cc_96 N_A_78_199#_M1003_g N_VPWR_c_275_n 0.0100933f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_78_199#_c_64_p N_VPWR_c_275_n 0.0141791f $X=1.98 $Y=1.96 $X2=0 $Y2=0
cc_98 N_A_78_199#_c_62_p A_292_297# 0.00613803f $X=1.735 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_78_199#_c_94_p N_VGND_M1008_d 0.00298767f $X=0.81 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_78_199#_c_53_n N_VGND_c_320_n 0.00438629f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_101 N_A_78_199#_c_55_n N_VGND_c_320_n 7.01852e-19 $X=0.69 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_78_199#_c_94_p N_VGND_c_320_n 0.0139733f $X=0.81 $Y=0.805 $X2=0 $Y2=0
cc_103 N_A_78_199#_c_94_p N_VGND_c_321_n 7.3395e-19 $X=0.81 $Y=0.805 $X2=0 $Y2=0
cc_104 N_A_78_199#_c_57_n N_VGND_c_321_n 0.00350332f $X=1.42 $Y=0.77 $X2=0 $Y2=0
cc_105 N_A_78_199#_c_53_n N_VGND_c_323_n 0.00575449f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_78_199#_c_94_p N_VGND_c_323_n 5.41497e-19 $X=0.81 $Y=0.805 $X2=0
+ $Y2=0
cc_107 N_A_78_199#_M1004_d N_VGND_c_325_n 0.00219239f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_108 N_A_78_199#_c_53_n N_VGND_c_325_n 0.0126455f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_78_199#_c_94_p N_VGND_c_325_n 0.00367143f $X=0.81 $Y=0.805 $X2=0
+ $Y2=0
cc_110 N_A_78_199#_c_57_n N_VGND_c_325_n 0.00687275f $X=1.42 $Y=0.77 $X2=0 $Y2=0
cc_111 N_A_78_199#_c_57_n N_A_215_47#_M1004_s 0.0031941f $X=1.42 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_112 N_A_78_199#_M1004_d N_A_215_47#_c_369_n 0.00323205f $X=1.485 $Y=0.235
+ $X2=0 $Y2=0
cc_113 N_A_78_199#_c_56_n N_A_215_47#_c_369_n 0.0173867f $X=1.62 $Y=0.73 $X2=0
+ $Y2=0
cc_114 N_A_78_199#_c_57_n N_A_215_47#_c_369_n 0.0167975f $X=1.42 $Y=0.77 $X2=0
+ $Y2=0
cc_115 N_A_78_199#_c_63_p N_A_215_47#_c_376_n 0.00492167f $X=1.927 $Y=1.805
+ $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_B2_M1002_g 0.034551f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_117 N_B1_c_125_n N_B2_c_158_n 0.0270099f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_127_n N_B2_c_159_n 0.0560029f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_119 B1 N_B2_c_160_n 0.0183737f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_c_127_n N_B2_c_160_n 0.00203072f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B1_M1006_g N_VPWR_c_279_n 0.00468308f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_122 N_B1_M1006_g N_VPWR_c_280_n 0.0162479f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_123 N_B1_M1006_g N_VPWR_c_275_n 0.00790314f $X=1.385 $Y=1.985 $X2=0 $Y2=0
cc_124 N_B1_c_125_n N_VGND_c_320_n 0.00241512f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_125 N_B1_c_125_n N_VGND_c_321_n 0.00366111f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_125_n N_VGND_c_325_n 0.0065944f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_125_n N_A_215_47#_c_369_n 0.00833791f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B2_M1002_g N_A2_M1007_g 0.01569f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_129 N_B2_M1002_g N_A2_c_194_n 8.99376e-19 $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_130 N_B2_c_159_n N_A2_c_194_n 7.56644e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_131 N_B2_c_160_n N_A2_c_194_n 0.021387f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B2_c_159_n N_A2_c_195_n 0.0219996f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B2_c_160_n N_A2_c_195_n 8.4425e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B2_c_158_n N_A2_c_196_n 0.0188951f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B2_M1002_g N_VPWR_c_279_n 0.0041991f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_136 N_B2_M1002_g N_VPWR_c_280_n 0.00284876f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_137 N_B2_M1002_g N_VPWR_c_275_n 0.00711876f $X=1.77 $Y=1.985 $X2=0 $Y2=0
cc_138 N_B2_c_158_n N_VGND_c_321_n 0.00366111f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B2_c_158_n N_VGND_c_325_n 0.00552681f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B2_c_158_n N_A_215_47#_c_369_n 0.0122623f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B2_c_160_n N_A_215_47#_c_369_n 0.00359996f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B2_c_159_n N_A_215_47#_c_376_n 2.22869e-19 $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_143 N_B2_c_160_n N_A_215_47#_c_376_n 0.00257395f $X=1.83 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A2_M1007_g N_A1_M1009_g 0.0493022f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_145 N_A2_c_194_n N_A1_M1009_g 9.18971e-19 $X=2.545 $Y=1.615 $X2=0 $Y2=0
cc_146 N_A2_c_194_n A1 0.0167247f $X=2.545 $Y=1.615 $X2=0 $Y2=0
cc_147 N_A2_c_195_n A1 6.48781e-19 $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_194_n N_A1_c_238_n 0.0042179f $X=2.545 $Y=1.615 $X2=0 $Y2=0
cc_149 N_A2_c_195_n N_A1_c_238_n 0.0493022f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A2_c_196_n N_A1_c_239_n 0.0274982f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_M1007_g N_VPWR_c_277_n 0.00216944f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_152 N_A2_c_194_n N_VPWR_c_277_n 0.00721642f $X=2.545 $Y=1.615 $X2=0 $Y2=0
cc_153 N_A2_M1007_g N_VPWR_c_279_n 0.00558092f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_154 A2 N_VPWR_c_279_n 0.00797507f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_155 N_A2_M1007_g N_VPWR_c_275_n 0.0104368f $X=2.39 $Y=1.985 $X2=0 $Y2=0
cc_156 A2 N_VPWR_c_275_n 0.00730368f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_157 A2 A_493_297# 0.00106578f $X=2.445 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_158 N_A2_c_196_n N_VGND_c_321_n 0.00420155f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_196_n N_VGND_c_322_n 0.00268723f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_196_n N_VGND_c_325_n 0.00590766f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_196_n N_A_215_47#_c_382_n 0.00218599f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_194_n N_A_215_47#_c_376_n 0.00596145f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_163 N_A2_c_195_n N_A_215_47#_c_376_n 0.00177877f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A2_c_196_n N_A_215_47#_c_376_n 0.0043816f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_194_n N_A_215_47#_c_370_n 0.016507f $X=2.545 $Y=1.615 $X2=0 $Y2=0
cc_166 N_A2_c_195_n N_A_215_47#_c_370_n 0.00152287f $X=2.33 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A2_c_196_n N_A_215_47#_c_370_n 0.00852077f $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_196_n N_A_215_47#_c_371_n 5.05864e-19 $X=2.32 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_M1009_g N_VPWR_c_277_n 0.0159507f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_170 A1 N_VPWR_c_277_n 0.025263f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_171 N_A1_c_238_n N_VPWR_c_277_n 0.00467935f $X=2.835 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_M1009_g N_VPWR_c_279_n 0.00544582f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_173 N_A1_M1009_g N_VPWR_c_275_n 0.00906165f $X=2.75 $Y=1.985 $X2=0 $Y2=0
cc_174 N_A1_c_239_n N_VGND_c_322_n 0.00268723f $X=2.845 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A1_c_239_n N_VGND_c_324_n 0.00421028f $X=2.845 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A1_c_239_n N_VGND_c_325_n 0.00663995f $X=2.845 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A1_c_239_n N_A_215_47#_c_376_n 4.48251e-19 $X=2.845 $Y=0.995 $X2=0
+ $Y2=0
cc_178 A1 N_A_215_47#_c_370_n 0.0281676f $X=2.905 $Y=1.105 $X2=0 $Y2=0
cc_179 N_A1_c_238_n N_A_215_47#_c_370_n 0.00452653f $X=2.835 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A1_c_239_n N_A_215_47#_c_370_n 0.00944054f $X=2.845 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A1_c_239_n N_A_215_47#_c_371_n 0.00576778f $X=2.845 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_X_c_262_n N_VPWR_c_278_n 0.0194075f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_183 N_X_M1003_s N_VPWR_c_275_n 0.00399293f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_184 N_X_c_262_n N_VPWR_c_275_n 0.0107063f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_185 N_X_c_262_n N_VGND_c_323_n 0.0109446f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_186 N_X_M1008_s N_VGND_c_325_n 0.00328323f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_187 N_X_c_262_n N_VGND_c_325_n 0.0100809f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_188 N_VPWR_c_275_n A_292_297# 0.0100452f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_189 N_VPWR_c_275_n A_493_297# 0.00279219f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_190 N_VGND_c_325_n N_A_215_47#_M1004_s 0.00211652f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_191 N_VGND_c_325_n N_A_215_47#_M1001_d 0.00283285f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_325_n N_A_215_47#_M1005_d 0.00210425f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_320_n N_A_215_47#_c_369_n 0.0106215f $X=0.68 $Y=0.38 $X2=0 $Y2=0
cc_194 N_VGND_c_321_n N_A_215_47#_c_369_n 0.0413054f $X=2.455 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_325_n N_A_215_47#_c_369_n 0.0320106f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_321_n N_A_215_47#_c_382_n 0.0164414f $X=2.455 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_325_n N_A_215_47#_c_382_n 0.0121819f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_M1000_d N_A_215_47#_c_370_n 0.00436355f $X=2.405 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_VGND_c_321_n N_A_215_47#_c_370_n 0.00211912f $X=2.455 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_c_322_n N_A_215_47#_c_370_n 0.012114f $X=2.54 $Y=0.36 $X2=0 $Y2=0
cc_201 N_VGND_c_324_n N_A_215_47#_c_370_n 0.00211912f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_325_n N_A_215_47#_c_370_n 0.00857469f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_324_n N_A_215_47#_c_371_n 0.01858f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_325_n N_A_215_47#_c_371_n 0.0125989f $X=2.99 $Y=0 $X2=0 $Y2=0

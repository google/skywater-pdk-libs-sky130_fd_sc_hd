* File: sky130_fd_sc_hd__a32o_1.spice
* Created: Thu Aug 27 14:05:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hd__a32o_1.spice.pex"
.subckt sky130_fd_sc_hd__a32o_1  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_93_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.167375 AS=0.2145 PD=1.165 PS=1.96 NRD=0.912 NRS=11.988 M=1 R=4.33333
+ SA=75000.3 SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1008 A_256_47# N_A3_M1008_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65 AD=0.0975
+ AS=0.167375 PD=0.95 PS=1.165 NRD=17.532 NRS=42.456 M=1 R=4.33333 SA=75000.9
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1009 A_346_47# N_A2_M1009_g A_256_47# VNB NSHORT L=0.15 W=0.65 AD=0.14625
+ AS=0.0975 PD=1.1 PS=0.95 NRD=31.38 NRS=17.532 M=1 R=4.33333 SA=75001.4
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1000 N_A_93_21#_M1000_d N_A1_M1000_g A_346_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.143 AS=0.14625 PD=1.09 PS=1.1 NRD=13.836 NRS=31.38 M=1 R=4.33333 SA=75002
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 A_584_47# N_B1_M1002_g N_A_93_21#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.143 PD=0.86 PS=1.09 NRD=9.228 NRS=15.684 M=1 R=4.33333
+ SA=75002.6 SB=75000.5 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B2_M1003_g A_584_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.06825 PD=1.83 PS=0.86 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.9 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_93_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1
+ AD=0.2425 AS=0.33 PD=1.485 PS=2.66 NRD=16.7253 NRS=12.7853 M=1 R=6.66667
+ SA=75000.3 SB=75002.9 A=0.15 P=2.3 MULT=1
MM1011 N_A_250_297#_M1011_d N_A3_M1011_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1
+ AD=0.165 AS=0.2425 PD=1.33 PS=1.485 NRD=4.9053 NRS=23.6203 M=1 R=6.66667
+ SA=75000.9 SB=75002.2 A=0.15 P=2.3 MULT=1
MM1007 N_VPWR_M1007_d N_A2_M1007_g N_A_250_297#_M1011_d VPB PHIGHVT L=0.15 W=1
+ AD=0.225 AS=0.165 PD=1.45 PS=1.33 NRD=16.7253 NRS=4.9053 M=1 R=6.66667
+ SA=75001.4 SB=75001.7 A=0.15 P=2.3 MULT=1
MM1010 N_A_250_297#_M1010_d N_A1_M1010_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1
+ AD=0.185 AS=0.225 PD=1.37 PS=1.45 NRD=7.8603 NRS=16.7253 M=1 R=6.66667
+ SA=75002 SB=75001.1 A=0.15 P=2.3 MULT=1
MM1006 N_A_93_21#_M1006_d N_B1_M1006_g N_A_250_297#_M1010_d VPB PHIGHVT L=0.15
+ W=1 AD=0.14 AS=0.185 PD=1.28 PS=1.37 NRD=0 NRS=9.8303 M=1 R=6.66667 SA=75002.5
+ SB=75000.6 A=0.15 P=2.3 MULT=1
MM1001 N_A_250_297#_M1001_d N_B2_M1001_g N_A_93_21#_M1006_d VPB PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=6.66667 SA=75002.9
+ SB=75000.2 A=0.15 P=2.3 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hd__a32o_1.spice.SKY130_FD_SC_HD__A32O_1.pxi"
*
.ends
*
*

* File: sky130_fd_sc_hd__and2b_1.pxi.spice
* Created: Tue Sep  1 18:57:09 2020
* 
x_PM_SKY130_FD_SC_HD__AND2B_1%A_N N_A_N_M1007_g N_A_N_M1003_g A_N A_N A_N
+ N_A_N_c_57_n PM_SKY130_FD_SC_HD__AND2B_1%A_N
x_PM_SKY130_FD_SC_HD__AND2B_1%A_27_413# N_A_27_413#_M1007_d N_A_27_413#_M1003_s
+ N_A_27_413#_M1004_g N_A_27_413#_M1001_g N_A_27_413#_c_93_n N_A_27_413#_c_94_n
+ N_A_27_413#_c_95_n N_A_27_413#_c_87_n N_A_27_413#_c_88_n N_A_27_413#_c_89_n
+ N_A_27_413#_c_90_n N_A_27_413#_c_91_n PM_SKY130_FD_SC_HD__AND2B_1%A_27_413#
x_PM_SKY130_FD_SC_HD__AND2B_1%B N_B_c_149_n N_B_M1000_g N_B_M1002_g B B
+ PM_SKY130_FD_SC_HD__AND2B_1%B
x_PM_SKY130_FD_SC_HD__AND2B_1%A_207_413# N_A_207_413#_M1001_s
+ N_A_207_413#_M1004_d N_A_207_413#_M1005_g N_A_207_413#_M1006_g
+ N_A_207_413#_c_187_n N_A_207_413#_c_181_n N_A_207_413#_c_182_n
+ N_A_207_413#_c_183_n N_A_207_413#_c_184_n N_A_207_413#_c_204_n
+ N_A_207_413#_c_185_n PM_SKY130_FD_SC_HD__AND2B_1%A_207_413#
x_PM_SKY130_FD_SC_HD__AND2B_1%VPWR N_VPWR_M1003_d N_VPWR_M1000_d N_VPWR_c_240_n
+ VPWR N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_239_n N_VPWR_c_244_n
+ N_VPWR_c_245_n N_VPWR_c_246_n PM_SKY130_FD_SC_HD__AND2B_1%VPWR
x_PM_SKY130_FD_SC_HD__AND2B_1%X N_X_M1005_d N_X_M1006_d N_X_c_278_n N_X_c_275_n
+ N_X_c_276_n X X X PM_SKY130_FD_SC_HD__AND2B_1%X
x_PM_SKY130_FD_SC_HD__AND2B_1%VGND N_VGND_M1007_s N_VGND_M1002_d N_VGND_c_293_n
+ N_VGND_c_294_n N_VGND_c_295_n VGND N_VGND_c_296_n N_VGND_c_297_n
+ N_VGND_c_298_n N_VGND_c_299_n PM_SKY130_FD_SC_HD__AND2B_1%VGND
cc_1 VNB N_A_N_M1007_g 0.0393258f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB A_N 0.0222233f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_A_N_c_57_n 0.0327074f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_4 VNB N_A_27_413#_M1004_g 0.0103574f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB N_A_27_413#_M1001_g 0.0214621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_413#_c_87_n 0.00391333f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_413#_c_88_n 0.00358141f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.19
cc_8 VNB N_A_27_413#_c_89_n 0.00438079f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.53
cc_9 VNB N_A_27_413#_c_90_n 0.00645363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_91_n 0.052475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_149_n 0.0175653f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_12 VNB N_B_M1002_g 0.0368067f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_13 VNB N_A_207_413#_c_181_n 0.00503027f $X=-0.19 $Y=-0.24 $X2=0.37 $Y2=1.325
cc_14 VNB N_A_207_413#_c_182_n 0.0147971f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=0.85
cc_15 VNB N_A_207_413#_c_183_n 0.00422495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_207_413#_c_184_n 0.0238813f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_17 VNB N_A_207_413#_c_185_n 0.0190083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_239_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.53
cc_19 VNB N_X_c_275_n 0.0236658f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_20 VNB N_X_c_276_n 0.00442969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB X 0.0149399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_293_n 0.0102466f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=2.275
cc_23 VNB N_VGND_c_294_n 0.0183467f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_24 VNB N_VGND_c_295_n 4.89851e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_296_n 0.0380941f $X=-0.19 $Y=-0.24 $X2=0.36 $Y2=1.16
cc_26 VNB N_VGND_c_297_n 0.0152458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_298_n 0.165382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_299_n 0.00523338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_N_M1003_g 0.0633079f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=2.275
cc_30 VPB A_N 0.0149437f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_31 VPB N_A_N_c_57_n 0.00746041f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_32 VPB N_A_27_413#_M1004_g 0.0504244f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_33 VPB N_A_27_413#_c_93_n 0.00221098f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_34 VPB N_A_27_413#_c_94_n 0.00839139f $X=-0.19 $Y=1.305 $X2=0.37 $Y2=1.325
cc_35 VPB N_A_27_413#_c_95_n 0.0109439f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=0.85
cc_36 VPB N_A_27_413#_c_88_n 0.00931385f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.19
cc_37 VPB N_B_c_149_n 0.0661509f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_38 VPB N_B_M1000_g 0.0257968f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.445
cc_39 VPB B 0.00634275f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_40 VPB N_A_207_413#_M1006_g 0.0254547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_207_413#_c_187_n 0.00613575f $X=-0.19 $Y=1.305 $X2=0.36 $Y2=1.16
cc_42 VPB N_A_207_413#_c_182_n 0.00730743f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=0.85
cc_43 VPB N_A_207_413#_c_183_n 0.00243367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_207_413#_c_184_n 0.00571563f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_45 VPB N_VPWR_c_240_n 0.00222879f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_46 VPB N_VPWR_c_241_n 0.015299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_242_n 0.0185743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_239_n 0.0457452f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.53
cc_49 VPB N_VPWR_c_244_n 0.00507571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_245_n 0.0177746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_246_n 0.0202241f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_278_n 0.00577345f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_53 VPB N_X_c_275_n 0.0120803f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_54 VPB X 0.0242568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_A_N_c_57_n N_A_27_413#_M1004_g 0.0239506f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_N_M1003_g N_A_27_413#_c_93_n 0.00187427f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_57 N_A_N_M1003_g N_A_27_413#_c_94_n 0.0188736f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_58 A_N N_A_27_413#_c_94_n 0.00808417f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_59 A_N N_A_27_413#_c_95_n 0.0158932f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_60 N_A_N_c_57_n N_A_27_413#_c_95_n 6.27406e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_N_M1007_g N_A_27_413#_c_87_n 0.00517713f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_62 A_N N_A_27_413#_c_87_n 0.00304427f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 A_N N_A_27_413#_c_88_n 0.0366831f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_N_c_57_n N_A_27_413#_c_88_n 0.00824519f $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_N_M1007_g N_A_27_413#_c_90_n 0.00287322f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_66 A_N N_A_27_413#_c_90_n 0.0268997f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A_N_M1007_g N_A_27_413#_c_91_n 0.0239506f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_68 A_N N_A_27_413#_c_91_n 3.71011e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_69 N_A_N_M1003_g N_A_207_413#_c_187_n 5.08711e-19 $X=0.47 $Y=2.275 $X2=0
+ $Y2=0
cc_70 N_A_N_M1003_g N_VPWR_c_240_n 0.0100411f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_71 N_A_N_M1003_g N_VPWR_c_241_n 0.00347311f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_72 N_A_N_M1003_g N_VPWR_c_239_n 0.00511644f $X=0.47 $Y=2.275 $X2=0 $Y2=0
cc_73 N_A_N_M1007_g N_VGND_c_294_n 0.0119879f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_74 A_N N_VGND_c_294_n 0.0213825f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_N_c_57_n N_VGND_c_294_n 8.25827e-19 $X=0.36 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_N_M1007_g N_VGND_c_296_n 0.0046653f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_N_M1007_g N_VGND_c_298_n 0.00872928f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_78 A_N N_VGND_c_298_n 0.00181266f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_27_413#_M1004_g N_B_c_149_n 0.0398731f $X=0.96 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_413#_c_91_n N_B_c_149_n 0.00440824f $X=1.065 $Y=0.97 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_27_413#_M1004_g N_B_M1002_g 2.81756e-19 $X=0.96 $Y=2.275 $X2=0 $Y2=0
cc_82 N_A_27_413#_M1001_g N_B_M1002_g 0.0439798f $X=1.41 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_27_413#_c_91_n N_B_M1002_g 0.00326355f $X=1.065 $Y=0.97 $X2=0 $Y2=0
cc_84 N_A_27_413#_M1004_g N_A_207_413#_c_187_n 0.0169169f $X=0.96 $Y=2.275 $X2=0
+ $Y2=0
cc_85 N_A_27_413#_c_93_n N_A_207_413#_c_187_n 0.00264049f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_86 N_A_27_413#_c_94_n N_A_207_413#_c_187_n 0.0191891f $X=0.615 $Y=1.9 $X2=0
+ $Y2=0
cc_87 N_A_27_413#_c_88_n N_A_207_413#_c_187_n 0.0235485f $X=0.732 $Y=1.785 $X2=0
+ $Y2=0
cc_88 N_A_27_413#_M1001_g N_A_207_413#_c_181_n 0.0054182f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_89 N_A_27_413#_c_89_n N_A_207_413#_c_181_n 0.0064045f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_90 N_A_27_413#_c_90_n N_A_207_413#_c_181_n 0.0103445f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_91 N_A_27_413#_c_91_n N_A_207_413#_c_181_n 0.00460502f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_92 N_A_27_413#_M1004_g N_A_207_413#_c_182_n 0.00622899f $X=0.96 $Y=2.275
+ $X2=0 $Y2=0
cc_93 N_A_27_413#_c_88_n N_A_207_413#_c_182_n 0.0211138f $X=0.732 $Y=1.785 $X2=0
+ $Y2=0
cc_94 N_A_27_413#_c_90_n N_A_207_413#_c_182_n 0.0274125f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_95 N_A_27_413#_c_91_n N_A_207_413#_c_182_n 0.0143099f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_M1001_g N_A_207_413#_c_204_n 0.00541516f $X=1.41 $Y=0.445
+ $X2=0 $Y2=0
cc_97 N_A_27_413#_c_89_n N_A_207_413#_c_204_n 0.018232f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_c_90_n N_A_207_413#_c_204_n 0.00236721f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_99 N_A_27_413#_c_91_n N_A_207_413#_c_204_n 0.00638575f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_100 N_A_27_413#_M1004_g N_VPWR_c_240_n 0.00319712f $X=0.96 $Y=2.275 $X2=0
+ $Y2=0
cc_101 N_A_27_413#_c_94_n N_VPWR_c_240_n 0.0245249f $X=0.615 $Y=1.9 $X2=0 $Y2=0
cc_102 N_A_27_413#_c_93_n N_VPWR_c_241_n 0.0102625f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_103 N_A_27_413#_c_94_n N_VPWR_c_241_n 0.0025049f $X=0.615 $Y=1.9 $X2=0 $Y2=0
cc_104 N_A_27_413#_M1003_s N_VPWR_c_239_n 0.00375546f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_105 N_A_27_413#_M1004_g N_VPWR_c_239_n 0.0104232f $X=0.96 $Y=2.275 $X2=0
+ $Y2=0
cc_106 N_A_27_413#_c_93_n N_VPWR_c_239_n 0.00640243f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_107 N_A_27_413#_c_94_n N_VPWR_c_239_n 0.00558823f $X=0.615 $Y=1.9 $X2=0 $Y2=0
cc_108 N_A_27_413#_M1004_g N_VPWR_c_245_n 0.00564994f $X=0.96 $Y=2.275 $X2=0
+ $Y2=0
cc_109 N_A_27_413#_M1001_g N_VGND_c_295_n 0.00185979f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_110 N_A_27_413#_M1001_g N_VGND_c_296_n 0.00388886f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_111 N_A_27_413#_c_89_n N_VGND_c_296_n 0.0140003f $X=0.68 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_27_413#_M1007_d N_VGND_c_298_n 0.00388065f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_113 N_A_27_413#_M1001_g N_VGND_c_298_n 0.00673847f $X=1.41 $Y=0.445 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_c_89_n N_VGND_c_298_n 0.00898311f $X=0.68 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_c_90_n N_VGND_c_298_n 0.00980064f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_116 N_A_27_413#_c_91_n N_VGND_c_298_n 0.00574233f $X=1.065 $Y=0.97 $X2=0
+ $Y2=0
cc_117 N_B_c_149_n N_A_207_413#_M1006_g 0.016411f $X=1.4 $Y=1.895 $X2=0 $Y2=0
cc_118 N_B_c_149_n N_A_207_413#_c_187_n 0.0107208f $X=1.4 $Y=1.895 $X2=0 $Y2=0
cc_119 B N_A_207_413#_c_187_n 0.025312f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_120 N_B_M1002_g N_A_207_413#_c_181_n 0.00551534f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B_c_149_n N_A_207_413#_c_182_n 0.0355669f $X=1.4 $Y=1.895 $X2=0 $Y2=0
cc_122 N_B_M1002_g N_A_207_413#_c_182_n 0.0156002f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_123 B N_A_207_413#_c_182_n 0.0317237f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_124 B N_A_207_413#_c_183_n 0.0147586f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_125 N_B_M1002_g N_A_207_413#_c_184_n 0.0219814f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_126 B N_A_207_413#_c_184_n 0.00180735f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_127 N_B_M1002_g N_A_207_413#_c_185_n 0.0247851f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_128 B N_VPWR_M1000_d 0.00763102f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_129 N_B_M1000_g N_VPWR_c_239_n 0.0119149f $X=1.4 $Y=2.275 $X2=0 $Y2=0
cc_130 B N_VPWR_c_239_n 0.00319716f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_131 N_B_M1000_g N_VPWR_c_245_n 0.00585385f $X=1.4 $Y=2.275 $X2=0 $Y2=0
cc_132 N_B_c_149_n N_VPWR_c_246_n 0.00202247f $X=1.4 $Y=1.895 $X2=0 $Y2=0
cc_133 N_B_M1000_g N_VPWR_c_246_n 0.00360298f $X=1.4 $Y=2.275 $X2=0 $Y2=0
cc_134 B N_VPWR_c_246_n 0.0447684f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_135 N_B_c_149_n N_X_c_278_n 5.09616e-19 $X=1.4 $Y=1.895 $X2=0 $Y2=0
cc_136 N_B_M1002_g N_VGND_c_295_n 0.015832f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B_M1002_g N_VGND_c_296_n 0.00486043f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B_M1002_g N_VGND_c_298_n 0.00822386f $X=1.8 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_207_413#_M1006_g N_VPWR_c_242_n 0.00566002f $X=2.29 $Y=1.985 $X2=0
+ $Y2=0
cc_140 N_A_207_413#_M1004_d N_VPWR_c_239_n 0.00308576f $X=1.035 $Y=2.065 $X2=0
+ $Y2=0
cc_141 N_A_207_413#_M1006_g N_VPWR_c_239_n 0.01253f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_142 N_A_207_413#_c_187_n N_VPWR_c_239_n 0.0105781f $X=1.18 $Y=2.225 $X2=0
+ $Y2=0
cc_143 N_A_207_413#_c_187_n N_VPWR_c_245_n 0.0129171f $X=1.18 $Y=2.225 $X2=0
+ $Y2=0
cc_144 N_A_207_413#_M1006_g N_VPWR_c_246_n 0.011029f $X=2.29 $Y=1.985 $X2=0
+ $Y2=0
cc_145 N_A_207_413#_M1006_g N_X_c_278_n 0.00402782f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_146 N_A_207_413#_c_182_n N_X_c_275_n 0.00521577f $X=1.88 $Y=1.135 $X2=0 $Y2=0
cc_147 N_A_207_413#_c_183_n N_X_c_275_n 0.029567f $X=2.22 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_207_413#_c_185_n N_X_c_275_n 0.0224779f $X=2.225 $Y=0.985 $X2=0 $Y2=0
cc_149 N_A_207_413#_M1006_g X 0.0132976f $X=2.29 $Y=1.985 $X2=0 $Y2=0
cc_150 N_A_207_413#_c_182_n N_VGND_c_295_n 0.00120465f $X=1.88 $Y=1.135 $X2=0
+ $Y2=0
cc_151 N_A_207_413#_c_183_n N_VGND_c_295_n 0.0153821f $X=2.22 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_207_413#_c_184_n N_VGND_c_295_n 6.3588e-19 $X=2.22 $Y=1.16 $X2=0
+ $Y2=0
cc_153 N_A_207_413#_c_185_n N_VGND_c_295_n 0.0106687f $X=2.225 $Y=0.985 $X2=0
+ $Y2=0
cc_154 N_A_207_413#_c_204_n N_VGND_c_296_n 0.0160751f $X=1.2 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_207_413#_c_185_n N_VGND_c_297_n 0.0046653f $X=2.225 $Y=0.985 $X2=0
+ $Y2=0
cc_156 N_A_207_413#_M1001_s N_VGND_c_298_n 0.00239557f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_157 N_A_207_413#_c_204_n N_VGND_c_298_n 0.0127737f $X=1.2 $Y=0.445 $X2=0
+ $Y2=0
cc_158 N_A_207_413#_c_185_n N_VGND_c_298_n 0.00895857f $X=2.225 $Y=0.985 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_239_n N_X_M1006_d 0.00220323f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_242_n X 0.0117541f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_239_n X 0.0109747f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_162 X N_VGND_c_297_n 0.0164883f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_163 N_X_M1005_d N_VGND_c_298_n 0.00387172f $X=2.365 $Y=0.235 $X2=0 $Y2=0
cc_164 X N_VGND_c_298_n 0.00914879f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_165 N_VGND_c_298_n A_297_47# 0.0100898f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24

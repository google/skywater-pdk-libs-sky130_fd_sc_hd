* File: sky130_fd_sc_hd__nor2b_4.spice.SKY130_FD_SC_HD__NOR2B_4.pxi
* Created: Thu Aug 27 14:31:52 2020
* 
x_PM_SKY130_FD_SC_HD__NOR2B_4%A N_A_c_86_n N_A_M1002_g N_A_M1001_g N_A_c_87_n
+ N_A_M1004_g N_A_M1012_g N_A_c_88_n N_A_M1008_g N_A_M1014_g N_A_c_89_n
+ N_A_M1009_g N_A_M1017_g A N_A_c_90_n N_A_c_91_n PM_SKY130_FD_SC_HD__NOR2B_4%A
x_PM_SKY130_FD_SC_HD__NOR2B_4%A_419_21# N_A_419_21#_M1003_s N_A_419_21#_M1011_s
+ N_A_419_21#_c_165_n N_A_419_21#_M1005_g N_A_419_21#_M1000_g
+ N_A_419_21#_c_166_n N_A_419_21#_M1010_g N_A_419_21#_M1006_g
+ N_A_419_21#_c_167_n N_A_419_21#_M1013_g N_A_419_21#_M1007_g
+ N_A_419_21#_c_168_n N_A_419_21#_M1016_g N_A_419_21#_M1015_g
+ N_A_419_21#_c_213_p N_A_419_21#_c_169_n N_A_419_21#_c_170_n
+ N_A_419_21#_c_171_n N_A_419_21#_c_180_n N_A_419_21#_c_172_n
+ N_A_419_21#_c_173_n N_A_419_21#_c_181_n N_A_419_21#_c_182_n
+ N_A_419_21#_c_174_n PM_SKY130_FD_SC_HD__NOR2B_4%A_419_21#
x_PM_SKY130_FD_SC_HD__NOR2B_4%B_N N_B_N_c_280_n N_B_N_M1003_g N_B_N_M1011_g B_N
+ N_B_N_c_282_n B_N PM_SKY130_FD_SC_HD__NOR2B_4%B_N
x_PM_SKY130_FD_SC_HD__NOR2B_4%A_27_297# N_A_27_297#_M1001_s N_A_27_297#_M1012_s
+ N_A_27_297#_M1017_s N_A_27_297#_M1006_d N_A_27_297#_M1015_d
+ N_A_27_297#_c_307_n N_A_27_297#_c_308_n N_A_27_297#_c_309_n
+ N_A_27_297#_c_355_p N_A_27_297#_c_310_n N_A_27_297#_c_311_n
+ N_A_27_297#_c_326_n N_A_27_297#_c_333_n N_A_27_297#_c_335_n
+ N_A_27_297#_c_339_n N_A_27_297#_c_312_n N_A_27_297#_c_313_n
+ N_A_27_297#_c_314_n N_A_27_297#_c_348_n PM_SKY130_FD_SC_HD__NOR2B_4%A_27_297#
x_PM_SKY130_FD_SC_HD__NOR2B_4%VPWR N_VPWR_M1001_d N_VPWR_M1014_d N_VPWR_M1011_d
+ N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n VPWR
+ N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_394_n
+ N_VPWR_c_385_n PM_SKY130_FD_SC_HD__NOR2B_4%VPWR
x_PM_SKY130_FD_SC_HD__NOR2B_4%Y N_Y_M1002_d N_Y_M1008_d N_Y_M1005_s N_Y_M1013_s
+ N_Y_M1000_s N_Y_M1007_s N_Y_c_462_n N_Y_c_451_n N_Y_c_452_n N_Y_c_473_n
+ N_Y_c_453_n N_Y_c_478_n N_Y_c_454_n N_Y_c_520_n N_Y_c_455_n N_Y_c_503_n
+ N_Y_c_459_n N_Y_c_521_n N_Y_c_456_n N_Y_c_457_n N_Y_c_460_n N_Y_c_461_n Y
+ PM_SKY130_FD_SC_HD__NOR2B_4%Y
x_PM_SKY130_FD_SC_HD__NOR2B_4%VGND N_VGND_M1002_s N_VGND_M1004_s N_VGND_M1009_s
+ N_VGND_M1010_d N_VGND_M1016_d N_VGND_M1003_d N_VGND_c_561_n N_VGND_c_562_n
+ N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n
+ N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n VGND
+ N_VGND_c_577_n N_VGND_c_578_n PM_SKY130_FD_SC_HD__NOR2B_4%VGND
cc_1 VNB N_A_c_86_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_87_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_3 VNB N_A_c_88_n 0.0158002f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=0.995
cc_4 VNB N_A_c_89_n 0.0159899f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.995
cc_5 VNB N_A_c_90_n 0.0105081f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_6 VNB N_A_c_91_n 0.0705911f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_7 VNB N_A_419_21#_c_165_n 0.0159866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_419_21#_c_166_n 0.0154145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_419_21#_c_167_n 0.0157727f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_419_21#_c_168_n 0.0197222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_419_21#_c_169_n 0.0442418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_419_21#_c_170_n 0.00335056f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_13 VNB N_A_419_21#_c_171_n 0.00362507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_419_21#_c_172_n 0.00134522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_419_21#_c_173_n 0.00117446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_419_21#_c_174_n 0.0592139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B_N_c_280_n 0.0246248f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_18 VNB B_N 0.0153622f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=0.995
cc_19 VNB N_B_N_c_282_n 0.0391805f $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.985
cc_20 VNB N_VPWR_c_385_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_451_n 0.00218078f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_22 VNB N_Y_c_452_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=0.56
cc_23 VNB N_Y_c_453_n 0.00410518f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_24 VNB N_Y_c_454_n 8.75799e-19 $X=-0.19 $Y=-0.24 $X2=0.91 $Y2=1.16
cc_25 VNB N_Y_c_455_n 0.00484696f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_26 VNB N_Y_c_456_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_457_n 0.00202522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_561_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.985
cc_29 VNB N_VGND_c_562_n 0.0349306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_563_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.325
cc_31 VNB N_VGND_c_564_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_32 VNB N_VGND_c_565_n 0.00358901f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_33 VNB N_VGND_c_566_n 0.0136791f $X=-0.19 $Y=-0.24 $X2=1.33 $Y2=1.16
cc_34 VNB N_VGND_c_567_n 0.0155909f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.16
cc_35 VNB N_VGND_c_568_n 0.0335702f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_36 VNB N_VGND_c_569_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_570_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_38 VNB N_VGND_c_571_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.175
cc_39 VNB N_VGND_c_572_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_573_n 0.0166678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_574_n 0.00323631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_575_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_576_n 0.00557475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_577_n 0.0183638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_578_n 0.269564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_A_M1001_g 0.0250431f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_47 VPB N_A_M1012_g 0.0179946f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_48 VPB N_A_M1014_g 0.0179946f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_49 VPB N_A_M1017_g 0.0184925f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_50 VPB N_A_c_91_n 0.0108798f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_51 VPB N_A_419_21#_M1000_g 0.0185987f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_52 VPB N_A_419_21#_M1006_g 0.0176224f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_53 VPB N_A_419_21#_M1007_g 0.0181069f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_54 VPB N_A_419_21#_M1015_g 0.023038f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_55 VPB N_A_419_21#_c_169_n 0.021667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_419_21#_c_180_n 0.00628437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_419_21#_c_181_n 0.0013846f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_419_21#_c_182_n 0.00513483f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_419_21#_c_174_n 0.010199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_B_N_M1011_g 0.0293544f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.985
cc_61 VPB B_N 0.00365122f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=0.995
cc_62 VPB N_B_N_c_282_n 0.0106215f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_63 VPB N_A_27_297#_c_307_n 0.0133394f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_64 VPB N_A_27_297#_c_308_n 0.0309889f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_65 VPB N_A_27_297#_c_309_n 0.00315624f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_66 VPB N_A_27_297#_c_310_n 0.00269564f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_67 VPB N_A_27_297#_c_311_n 0.00422862f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_297#_c_312_n 0.00217609f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_69 VPB N_A_27_297#_c_313_n 0.00751666f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.16
cc_70 VPB N_A_27_297#_c_314_n 0.00131915f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_71 VPB N_VPWR_c_386_n 3.95446e-19 $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.985
cc_72 VPB N_VPWR_c_387_n 0.00221708f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=0.56
cc_73 VPB N_VPWR_c_388_n 0.0141086f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.325
cc_74 VPB N_VPWR_c_389_n 0.0516419f $X=-0.19 $Y=1.305 $X2=1.33 $Y2=1.985
cc_75 VPB N_VPWR_c_390_n 0.0155059f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.985
cc_76 VPB N_VPWR_c_391_n 0.0124915f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_77 VPB N_VPWR_c_392_n 0.0689736f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_78 VPB N_VPWR_c_393_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_394_n 0.00353635f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_80 VPB N_VPWR_c_385_n 0.0531792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_Y_c_454_n 0.00117101f $X=-0.19 $Y=1.305 $X2=0.91 $Y2=1.16
cc_82 VPB N_Y_c_459_n 0.00172897f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.175
cc_83 VPB N_Y_c_460_n 2.78665e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_Y_c_461_n 0.00309212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 N_A_c_89_n N_A_419_21#_c_165_n 0.0194866f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_M1017_g N_A_419_21#_M1000_g 0.0194866f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_c_90_n N_A_419_21#_c_174_n 9.19453e-19 $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_c_91_n N_A_419_21#_c_174_n 0.0194866f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_c_90_n N_A_27_297#_c_307_n 4.10066e-19 $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_A_27_297#_c_309_n 0.0138768f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_91 N_A_M1012_g N_A_27_297#_c_309_n 0.0136248f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_92 N_A_c_90_n N_A_27_297#_c_309_n 0.046205f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_c_91_n N_A_27_297#_c_309_n 0.00213789f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_M1014_g N_A_27_297#_c_310_n 0.0136248f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_M1017_g N_A_27_297#_c_310_n 0.0118246f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_96 N_A_c_90_n N_A_27_297#_c_310_n 0.0404893f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_c_91_n N_A_27_297#_c_310_n 0.00213789f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_M1017_g N_A_27_297#_c_311_n 0.00167295f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_99 N_A_c_90_n N_A_27_297#_c_311_n 3.67829e-19 $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_M1014_g N_A_27_297#_c_326_n 4.50937e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_101 N_A_M1017_g N_A_27_297#_c_326_n 0.00997294f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_102 N_A_c_90_n N_A_27_297#_c_314_n 0.0132812f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_c_91_n N_A_27_297#_c_314_n 0.00221654f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_M1001_g N_VPWR_c_386_n 0.0129691f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_105 N_A_M1012_g N_VPWR_c_386_n 0.0110282f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_106 N_A_M1014_g N_VPWR_c_386_n 6.32588e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_107 N_A_M1012_g N_VPWR_c_387_n 6.27883e-19 $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_108 N_A_M1014_g N_VPWR_c_387_n 0.0106598f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_109 N_A_M1017_g N_VPWR_c_387_n 0.00279634f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_VPWR_c_390_n 0.0046653f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_M1012_g N_VPWR_c_391_n 0.0046653f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_112 N_A_M1014_g N_VPWR_c_391_n 0.0046653f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_113 N_A_M1017_g N_VPWR_c_392_n 0.00539841f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_114 N_A_M1001_g N_VPWR_c_385_n 0.00886468f $X=0.49 $Y=1.985 $X2=0 $Y2=0
cc_115 N_A_M1012_g N_VPWR_c_385_n 0.00789179f $X=0.91 $Y=1.985 $X2=0 $Y2=0
cc_116 N_A_M1014_g N_VPWR_c_385_n 0.00789179f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_117 N_A_M1017_g N_VPWR_c_385_n 0.00949176f $X=1.75 $Y=1.985 $X2=0 $Y2=0
cc_118 N_A_c_86_n N_Y_c_462_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_c_87_n N_Y_c_462_n 0.00630972f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_88_n N_Y_c_462_n 5.22228e-19 $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A_c_87_n N_Y_c_451_n 0.00870364f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_88_n N_Y_c_451_n 0.00870364f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_90_n N_Y_c_451_n 0.036111f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_91_n N_Y_c_451_n 0.00222133f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_c_86_n N_Y_c_452_n 0.00262807f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_87_n N_Y_c_452_n 0.00113286f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_90_n N_Y_c_452_n 0.0265405f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_91_n N_Y_c_452_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_c_87_n N_Y_c_473_n 5.22228e-19 $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_88_n N_Y_c_473_n 0.00630972f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_89_n N_Y_c_473_n 0.00630972f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_89_n N_Y_c_453_n 0.00896662f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_90_n N_Y_c_453_n 0.00651491f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_89_n N_Y_c_478_n 5.22228e-19 $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_90_n N_Y_c_454_n 0.00659349f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_91_n N_Y_c_454_n 0.00132221f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_88_n N_Y_c_456_n 0.00113286f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_89_n N_Y_c_456_n 0.00113286f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_90_n N_Y_c_456_n 0.0265405f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_c_91_n N_Y_c_456_n 0.00230339f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A_c_86_n N_VGND_c_562_n 0.0036723f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_87_n N_VGND_c_563_n 0.00146448f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_88_n N_VGND_c_563_n 0.00146448f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_89_n N_VGND_c_564_n 0.00146448f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_86_n N_VGND_c_569_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_87_n N_VGND_c_569_n 0.00423334f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_88_n N_VGND_c_571_n 0.00423334f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_89_n N_VGND_c_571_n 0.00423334f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_86_n N_VGND_c_578_n 0.0104744f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_c_87_n N_VGND_c_578_n 0.0057163f $X=0.91 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_88_n N_VGND_c_578_n 0.0057163f $X=1.33 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_89_n N_VGND_c_578_n 0.0057435f $X=1.75 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_419_21#_c_170_n N_B_N_c_280_n 0.00457189f $X=4.19 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_419_21#_c_171_n N_B_N_c_280_n 0.00617045f $X=4.15 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_419_21#_c_172_n N_B_N_c_280_n 0.00323581f $X=4.19 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_419_21#_c_180_n N_B_N_M1011_g 0.00820023f $X=4.19 $Y=2.34 $X2=0 $Y2=0
cc_157 N_A_419_21#_c_181_n N_B_N_M1011_g 0.0032678f $X=4.19 $Y=1.66 $X2=0 $Y2=0
cc_158 N_A_419_21#_c_173_n B_N 0.0174258f $X=4.15 $Y=1.175 $X2=0 $Y2=0
cc_159 N_A_419_21#_c_182_n B_N 0.00350706f $X=4.19 $Y=1.575 $X2=0 $Y2=0
cc_160 N_A_419_21#_c_169_n N_B_N_c_282_n 0.0209283f $X=3.98 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_419_21#_c_173_n N_B_N_c_282_n 0.00164603f $X=4.15 $Y=1.175 $X2=0
+ $Y2=0
cc_162 N_A_419_21#_c_182_n N_B_N_c_282_n 0.00696913f $X=4.19 $Y=1.575 $X2=0
+ $Y2=0
cc_163 N_A_419_21#_M1000_g N_A_27_297#_c_311_n 0.00335853f $X=2.17 $Y=1.985
+ $X2=0 $Y2=0
cc_164 N_A_419_21#_M1000_g N_A_27_297#_c_326_n 0.00843121f $X=2.17 $Y=1.985
+ $X2=0 $Y2=0
cc_165 N_A_419_21#_M1006_g N_A_27_297#_c_326_n 5.45807e-19 $X=2.59 $Y=1.985
+ $X2=0 $Y2=0
cc_166 N_A_419_21#_M1000_g N_A_27_297#_c_333_n 0.0101149f $X=2.17 $Y=1.985 $X2=0
+ $Y2=0
cc_167 N_A_419_21#_M1006_g N_A_27_297#_c_333_n 0.00792493f $X=2.59 $Y=1.985
+ $X2=0 $Y2=0
cc_168 N_A_419_21#_M1000_g N_A_27_297#_c_335_n 4.89808e-19 $X=2.17 $Y=1.985
+ $X2=0 $Y2=0
cc_169 N_A_419_21#_M1006_g N_A_27_297#_c_335_n 0.00534818f $X=2.59 $Y=1.985
+ $X2=0 $Y2=0
cc_170 N_A_419_21#_M1007_g N_A_27_297#_c_335_n 0.00534818f $X=3.01 $Y=1.985
+ $X2=0 $Y2=0
cc_171 N_A_419_21#_M1015_g N_A_27_297#_c_335_n 4.89808e-19 $X=3.43 $Y=1.985
+ $X2=0 $Y2=0
cc_172 N_A_419_21#_M1007_g N_A_27_297#_c_339_n 0.00795376f $X=3.01 $Y=1.985
+ $X2=0 $Y2=0
cc_173 N_A_419_21#_M1015_g N_A_27_297#_c_339_n 0.0101149f $X=3.43 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_419_21#_M1015_g N_A_27_297#_c_312_n 7.12665e-19 $X=3.43 $Y=1.985
+ $X2=0 $Y2=0
cc_175 N_A_419_21#_c_180_n N_A_27_297#_c_312_n 0.0150382f $X=4.19 $Y=2.34 $X2=0
+ $Y2=0
cc_176 N_A_419_21#_M1007_g N_A_27_297#_c_313_n 5.45229e-19 $X=3.01 $Y=1.985
+ $X2=0 $Y2=0
cc_177 N_A_419_21#_M1015_g N_A_27_297#_c_313_n 0.00921886f $X=3.43 $Y=1.985
+ $X2=0 $Y2=0
cc_178 N_A_419_21#_c_213_p N_A_27_297#_c_313_n 0.0178299f $X=4.025 $Y=1.175
+ $X2=0 $Y2=0
cc_179 N_A_419_21#_c_169_n N_A_27_297#_c_313_n 0.00774573f $X=3.98 $Y=1.16 $X2=0
+ $Y2=0
cc_180 N_A_419_21#_c_181_n N_A_27_297#_c_313_n 0.0605155f $X=4.19 $Y=1.66 $X2=0
+ $Y2=0
cc_181 N_A_419_21#_M1006_g N_A_27_297#_c_348_n 7.04098e-19 $X=2.59 $Y=1.985
+ $X2=0 $Y2=0
cc_182 N_A_419_21#_M1007_g N_A_27_297#_c_348_n 7.04098e-19 $X=3.01 $Y=1.985
+ $X2=0 $Y2=0
cc_183 N_A_419_21#_M1000_g N_VPWR_c_392_n 0.00357835f $X=2.17 $Y=1.985 $X2=0
+ $Y2=0
cc_184 N_A_419_21#_M1006_g N_VPWR_c_392_n 0.00357835f $X=2.59 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_419_21#_M1007_g N_VPWR_c_392_n 0.00357835f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_186 N_A_419_21#_M1015_g N_VPWR_c_392_n 0.00357835f $X=3.43 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_419_21#_c_180_n N_VPWR_c_392_n 0.0210244f $X=4.19 $Y=2.34 $X2=0 $Y2=0
cc_188 N_A_419_21#_M1011_s N_VPWR_c_385_n 0.00217517f $X=4.055 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_419_21#_M1000_g N_VPWR_c_385_n 0.00525234f $X=2.17 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_A_419_21#_M1006_g N_VPWR_c_385_n 0.00522513f $X=2.59 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_A_419_21#_M1007_g N_VPWR_c_385_n 0.00522513f $X=3.01 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_419_21#_M1015_g N_VPWR_c_385_n 0.0065512f $X=3.43 $Y=1.985 $X2=0
+ $Y2=0
cc_193 N_A_419_21#_c_180_n N_VPWR_c_385_n 0.0124163f $X=4.19 $Y=2.34 $X2=0 $Y2=0
cc_194 N_A_419_21#_c_165_n N_Y_c_473_n 5.22228e-19 $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_419_21#_c_165_n N_Y_c_453_n 0.0117699f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_419_21#_c_165_n N_Y_c_478_n 0.00630972f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_419_21#_c_166_n N_Y_c_478_n 0.00630972f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_419_21#_c_167_n N_Y_c_478_n 5.22228e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_419_21#_c_165_n N_Y_c_454_n 0.00241567f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_419_21#_M1000_g N_Y_c_454_n 0.00322994f $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_201 N_A_419_21#_c_166_n N_Y_c_454_n 0.00293518f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_419_21#_M1006_g N_Y_c_454_n 0.0039358f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_203 N_A_419_21#_c_167_n N_Y_c_454_n 5.12484e-19 $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_419_21#_M1007_g N_Y_c_454_n 6.86349e-19 $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_205 N_A_419_21#_c_213_p N_Y_c_454_n 0.0158053f $X=4.025 $Y=1.175 $X2=0 $Y2=0
cc_206 N_A_419_21#_c_174_n N_Y_c_454_n 0.029274f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_419_21#_c_166_n N_Y_c_455_n 0.00468086f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_419_21#_c_167_n N_Y_c_455_n 0.0098365f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_419_21#_c_168_n N_Y_c_455_n 0.00262807f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_419_21#_c_213_p N_Y_c_455_n 0.0449595f $X=4.025 $Y=1.175 $X2=0 $Y2=0
cc_211 N_A_419_21#_c_174_n N_Y_c_455_n 0.00470394f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_419_21#_c_166_n N_Y_c_503_n 5.22228e-19 $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_419_21#_c_167_n N_Y_c_503_n 0.00630972f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_419_21#_c_168_n N_Y_c_503_n 0.00539651f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_419_21#_M1015_g N_Y_c_459_n 0.0012406f $X=3.43 $Y=1.985 $X2=0 $Y2=0
cc_216 N_A_419_21#_c_213_p N_Y_c_459_n 0.0138639f $X=4.025 $Y=1.175 $X2=0 $Y2=0
cc_217 N_A_419_21#_c_174_n N_Y_c_459_n 0.00222344f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_419_21#_c_165_n N_Y_c_457_n 0.00221107f $X=2.17 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_419_21#_c_166_n N_Y_c_457_n 0.00409494f $X=2.59 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_419_21#_M1000_g N_Y_c_460_n 5.53367e-19 $X=2.17 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_419_21#_M1006_g N_Y_c_460_n 0.00642186f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_222 N_A_419_21#_M1006_g N_Y_c_461_n 0.00611412f $X=2.59 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_419_21#_M1007_g N_Y_c_461_n 0.013606f $X=3.01 $Y=1.985 $X2=0 $Y2=0
cc_224 N_A_419_21#_c_213_p N_Y_c_461_n 0.0251164f $X=4.025 $Y=1.175 $X2=0 $Y2=0
cc_225 N_A_419_21#_c_174_n N_Y_c_461_n 0.00236161f $X=3.505 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_419_21#_c_165_n N_VGND_c_564_n 0.00146448f $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_419_21#_c_166_n N_VGND_c_565_n 0.00146448f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_419_21#_c_167_n N_VGND_c_565_n 0.00146448f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_229 N_A_419_21#_c_168_n N_VGND_c_566_n 0.00367742f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_419_21#_c_213_p N_VGND_c_566_n 0.0234825f $X=4.025 $Y=1.175 $X2=0
+ $Y2=0
cc_231 N_A_419_21#_c_169_n N_VGND_c_566_n 0.00739466f $X=3.98 $Y=1.16 $X2=0
+ $Y2=0
cc_232 N_A_419_21#_c_170_n N_VGND_c_566_n 0.0512575f $X=4.19 $Y=0.39 $X2=0 $Y2=0
cc_233 N_A_419_21#_c_171_n N_VGND_c_568_n 0.00117072f $X=4.15 $Y=1.075 $X2=0
+ $Y2=0
cc_234 N_A_419_21#_c_165_n N_VGND_c_573_n 0.00423334f $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_419_21#_c_166_n N_VGND_c_573_n 0.00423261f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_419_21#_c_167_n N_VGND_c_575_n 0.00423334f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_419_21#_c_168_n N_VGND_c_575_n 0.00541359f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_419_21#_c_170_n N_VGND_c_577_n 0.020984f $X=4.19 $Y=0.39 $X2=0 $Y2=0
cc_239 N_A_419_21#_M1003_s N_VGND_c_578_n 0.00225715f $X=4.045 $Y=0.235 $X2=0
+ $Y2=0
cc_240 N_A_419_21#_c_165_n N_VGND_c_578_n 0.0057435f $X=2.17 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_419_21#_c_166_n N_VGND_c_578_n 0.00571497f $X=2.59 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_419_21#_c_167_n N_VGND_c_578_n 0.0057163f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_419_21#_c_168_n N_VGND_c_578_n 0.0108276f $X=3.43 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_419_21#_c_170_n N_VGND_c_578_n 0.0124119f $X=4.19 $Y=0.39 $X2=0 $Y2=0
cc_245 N_B_N_M1011_g N_VPWR_c_389_n 0.00463894f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_246 B_N N_VPWR_c_389_n 0.0325355f $X=4.75 $Y=1.105 $X2=0 $Y2=0
cc_247 N_B_N_c_282_n N_VPWR_c_389_n 0.00580252f $X=4.61 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B_N_M1011_g N_VPWR_c_392_n 0.00541359f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_249 N_B_N_M1011_g N_VPWR_c_385_n 0.0119208f $X=4.4 $Y=1.985 $X2=0 $Y2=0
cc_250 N_B_N_c_280_n N_VGND_c_566_n 0.0023653f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_N_c_280_n N_VGND_c_568_n 0.00500932f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_252 B_N N_VGND_c_568_n 0.0239559f $X=4.75 $Y=1.105 $X2=0 $Y2=0
cc_253 N_B_N_c_282_n N_VGND_c_568_n 0.0063933f $X=4.61 $Y=1.16 $X2=0 $Y2=0
cc_254 N_B_N_c_280_n N_VGND_c_577_n 0.00541359f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_255 N_B_N_c_280_n N_VGND_c_578_n 0.0119208f $X=4.4 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_27_297#_c_309_n N_VPWR_M1001_d 0.00166915f $X=1.035 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_257 N_A_27_297#_c_310_n N_VPWR_M1014_d 0.00166915f $X=1.795 $Y=1.56 $X2=0
+ $Y2=0
cc_258 N_A_27_297#_c_309_n N_VPWR_c_386_n 0.0172742f $X=1.035 $Y=1.56 $X2=0
+ $Y2=0
cc_259 N_A_27_297#_c_310_n N_VPWR_c_387_n 0.0150746f $X=1.795 $Y=1.56 $X2=0
+ $Y2=0
cc_260 N_A_27_297#_c_308_n N_VPWR_c_390_n 0.0194075f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_355_p N_VPWR_c_391_n 0.0113958f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_262 N_A_27_297#_c_326_n N_VPWR_c_392_n 0.0190403f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_c_333_n N_VPWR_c_392_n 0.0286211f $X=2.635 $Y=2.38 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_c_339_n N_VPWR_c_392_n 0.0286211f $X=3.475 $Y=2.38 $X2=0
+ $Y2=0
cc_265 N_A_27_297#_c_312_n N_VPWR_c_392_n 0.0247353f $X=3.665 $Y=2.295 $X2=0
+ $Y2=0
cc_266 N_A_27_297#_c_348_n N_VPWR_c_392_n 0.0187749f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_267 N_A_27_297#_M1001_s N_VPWR_c_385_n 0.00399293f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_M1012_s N_VPWR_c_385_n 0.00562358f $X=0.985 $Y=1.485 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_M1017_s N_VPWR_c_385_n 0.00215201f $X=1.825 $Y=1.485 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_M1006_d N_VPWR_c_385_n 0.00215201f $X=2.665 $Y=1.485 $X2=0
+ $Y2=0
cc_271 N_A_27_297#_M1015_d N_VPWR_c_385_n 0.00225715f $X=3.505 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_27_297#_c_308_n N_VPWR_c_385_n 0.0107063f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_273 N_A_27_297#_c_355_p N_VPWR_c_385_n 0.00646998f $X=1.12 $Y=2.3 $X2=0 $Y2=0
cc_274 N_A_27_297#_c_326_n N_VPWR_c_385_n 0.0122896f $X=1.96 $Y=2.295 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_333_n N_VPWR_c_385_n 0.0178969f $X=2.635 $Y=2.38 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_339_n N_VPWR_c_385_n 0.0178969f $X=3.475 $Y=2.38 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_c_312_n N_VPWR_c_385_n 0.0144248f $X=3.665 $Y=2.295 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_c_348_n N_VPWR_c_385_n 0.0122096f $X=2.8 $Y=2.38 $X2=0 $Y2=0
cc_279 N_A_27_297#_c_333_n N_Y_M1000_s 0.00312348f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_280 N_A_27_297#_c_339_n N_Y_M1007_s 0.00312348f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_281 N_A_27_297#_c_311_n N_Y_c_453_n 0.0117136f $X=1.96 $Y=1.665 $X2=0 $Y2=0
cc_282 N_A_27_297#_c_333_n N_Y_c_520_n 0.0118865f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_283 N_A_27_297#_c_339_n N_Y_c_521_n 0.0118865f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_311_n N_Y_c_460_n 0.010246f $X=1.96 $Y=1.665 $X2=0 $Y2=0
cc_285 N_A_27_297#_c_333_n N_Y_c_460_n 0.00315368f $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_286 N_A_27_297#_M1006_d N_Y_c_461_n 0.00176936f $X=2.665 $Y=1.485 $X2=0 $Y2=0
cc_287 N_A_27_297#_c_333_n N_Y_c_461_n 2.43246e-19 $X=2.635 $Y=2.38 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_335_n N_Y_c_461_n 0.0159581f $X=2.8 $Y=2.02 $X2=0 $Y2=0
cc_289 N_A_27_297#_c_339_n N_Y_c_461_n 0.00321626f $X=3.475 $Y=2.38 $X2=0 $Y2=0
cc_290 N_A_27_297#_c_307_n N_VGND_c_562_n 0.0113923f $X=0.225 $Y=1.665 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_385_n N_Y_M1000_s 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_385_n N_Y_M1007_s 0.00216833f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_293 N_Y_c_451_n N_VGND_M1004_s 0.00162089f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_294 N_Y_c_453_n N_VGND_M1009_s 0.00162089f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_295 N_Y_c_455_n N_VGND_M1010_d 0.00162089f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_296 N_Y_c_452_n N_VGND_c_562_n 0.00835667f $X=0.865 $Y=0.815 $X2=0 $Y2=0
cc_297 N_Y_c_451_n N_VGND_c_563_n 0.0122559f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_298 N_Y_c_453_n N_VGND_c_564_n 0.0122559f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_299 N_Y_c_455_n N_VGND_c_565_n 0.0122559f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_300 N_Y_c_455_n N_VGND_c_566_n 0.00836079f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_301 N_Y_c_462_n N_VGND_c_569_n 0.0188551f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_302 N_Y_c_451_n N_VGND_c_569_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_303 N_Y_c_451_n N_VGND_c_571_n 0.00198695f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_304 N_Y_c_473_n N_VGND_c_571_n 0.0188551f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_305 N_Y_c_453_n N_VGND_c_571_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_306 N_Y_c_453_n N_VGND_c_573_n 0.00198695f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_307 N_Y_c_478_n N_VGND_c_573_n 0.0188977f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_308 N_Y_c_455_n N_VGND_c_573_n 9.11858e-19 $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_309 N_Y_c_457_n N_VGND_c_573_n 0.00118043f $X=2.42 $Y=0.815 $X2=0 $Y2=0
cc_310 N_Y_c_455_n N_VGND_c_575_n 0.00198695f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_311 N_Y_c_503_n N_VGND_c_575_n 0.0188551f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_312 N_Y_M1002_d N_VGND_c_578_n 0.00215201f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_313 N_Y_M1008_d N_VGND_c_578_n 0.00215201f $X=1.405 $Y=0.235 $X2=0 $Y2=0
cc_314 N_Y_M1005_s N_VGND_c_578_n 0.00215201f $X=2.245 $Y=0.235 $X2=0 $Y2=0
cc_315 N_Y_M1013_s N_VGND_c_578_n 0.00215201f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_c_462_n N_VGND_c_578_n 0.0122069f $X=0.7 $Y=0.39 $X2=0 $Y2=0
cc_317 N_Y_c_451_n N_VGND_c_578_n 0.00835832f $X=1.375 $Y=0.815 $X2=0 $Y2=0
cc_318 N_Y_c_473_n N_VGND_c_578_n 0.0122069f $X=1.54 $Y=0.39 $X2=0 $Y2=0
cc_319 N_Y_c_453_n N_VGND_c_578_n 0.00835832f $X=2.215 $Y=0.815 $X2=0 $Y2=0
cc_320 N_Y_c_478_n N_VGND_c_578_n 0.0122182f $X=2.38 $Y=0.39 $X2=0 $Y2=0
cc_321 N_Y_c_455_n N_VGND_c_578_n 0.00663839f $X=3.055 $Y=0.815 $X2=0 $Y2=0
cc_322 N_Y_c_503_n N_VGND_c_578_n 0.0122069f $X=3.22 $Y=0.39 $X2=0 $Y2=0
cc_323 N_Y_c_457_n N_VGND_c_578_n 0.001841f $X=2.42 $Y=0.815 $X2=0 $Y2=0
